
module DenseBlackBox5f433e8bf5(
  input clock,
  input [9:0] readAddr,
  output [8191:0] out
);

reg [8191:0] rom_uints [1023:0];
initial
begin
rom_uints[0] = 8192'h10000100cc1d0003f000000010030c00000c000000005003404c0000100c0c00100174f0070301001303000713440f303c00000f0347300c00004000dc0000100103030404030001000000040300541074000d330403000c04500000003c100100f4310003043300500071000000000400110c000f00000c00030c30c000c00000c04000030f00030c00400000000103001c00030004c0070c50000040c10003100040000400000104000c00000c000c4003000000000300001000c00c00000303c00000c40c35d03450003c000f53430c04470c00cc3000043c00001d00100031030000000000000403001c40500c00004c0f000000004000000301340000c403001004c0000f0340f41450000f001004cd5030040400100000030f5d03033400d1000003001d0f00000c0000405d103000340c1c000000010010300c310000074444000500100000040c00c000400f001101041dc0000003cc0451055001c004050c0c330703cc00300700011c4404c0000d10030c44310700410100000d000f300d00505000043c0c00004030010d0f003400041400000f4013000400000c000f4000f00400050400300004070c3c004c01cc340c10000d0001d0030cfc04004c00040000030000c300304c0000000000300c00301133cc34c30c0000004c000c1ccc0040040500f1cc1000000d0011003c51c0000000001044003c0000000044d30c0411730000001000010f00000401400005310c000000000004004c04040f00341403003f000c0400144000000c5044000f03cf0c30040303000000000000400010001c0c300c3000c0000000c00f03000000034000c104000500000000c40010f30004400c030700000011000c0001cc000000000030f00035000400400013000300030000300400440004031c103ccf003010c000f4c300470003000c00000f0c04000011434300030033113f001c04000001401c0000000cc0070011311703000000300000001400000c04040401400400030031000c044ccfc300c30000000c000000403040000100cf3c0011003700400000c0003404003031c30d00000000000f040000140403330000070c00cc3000003000003100070400c3005c04c00d040cccc300c303030cc30104001d5130071030c10d01034c40c7100c0351340c000c33000f0000000300000000f4d00015000c410c0304000000000000c0040c00000304010004c100c000001047110f0c000151000003c0000304000000000c00410400040003300c430400500050c10c000003c0ff44000000c700000044500030000c0c0003c40003c00057440c0c0030000000000004005c040c1f140400400000000141c304c0000000f0304001c3000dc00c103133050004400000001cc0c00000001f00000c00040d000c00c400000c000000c00c040000;
rom_uints[1] = 8192'h30000000001100c3c0000000000004000100000000c700404000000343405000000000001000000010001010c0cc3c0000d000c403003301000000c0000000c0c03000441000100000003000000100c00000c0000001007000c00000c103404033d0d0004000000000c000c0c000f001f000004040400100c300c00000000100400c001000000000001000000000030041001000000000c100000040c00000c000d0400003014000c100000143c003004453000000000c00c00010f03000000c1100510000c000c0000003400040f13440003300400000c101c00c10c00000f10300000000100000d03047000100004000400000c00040000130000100000007105000d100000300c04000000000000001c001000040004030c00000c0107000010000000010c30074c0000300f0300000c003413310000000030000300030c000000033d01400000001000000c040c10000404001444001010001000301cc0000003000103000000010004310c3c0000000000003000c4004cc03000000c030000000c000010040000000f00001cf00000000400000400003003300000300000300000001300000000040114040c30340300000000000000370c0c01000d001f000c0000000400000c00000000110c0c00001c000407000300001000040c04010c330440000c00041c00033001000c000000000c000c000c0000040300000000044c0cc000370403000333070001000c003c000003030c03000d000c0d030000010c0c000c0300000000003001c0000001000c00000c000c0c0000000010000004400000010100100c000001000c003d00000000000f0f1c1410030440001000000c0300000300000000000003100000041005000c000c0000000400040000311c0040000000000c0003c00000000004cc300c1004000000000400400c33001c000300000310005040000c001c000013c40c0c00000030f00d0d00000000100004340000010000000000000300000000400000300001000000001c0003001000000000400000000dc30cc0c00c1000000340cc0000300000001d05000000000cc330000cc00404000000300700000000310107000010000300c010070000011c7000000000000c00010000000c000000340cc00c00040000c00030000cc400000c00100c10000000300000074004000003400100400c00000c000c0310000001010c00400c0c0d0c00040030000044040000000010030c0c000000000c0400c00140000000000000003c0c000404000c0001104c300000710110000f00000c0010d000000000040300000c000040000c00000c00030c00000000000444000004100300000004403c0c000c0c0c0c04000000000310071c01000400000000003c000c0000101f30040400c01000000410000f000400011f10000004000c040;
rom_uints[2] = 8192'hd11000001400c40500000003000003100c0303001300010000310300c303c0107c0c0040c5c300c0000f00030101700c0041100c000c0c4401071000030005000140000c00c000d00000110331c03000040510004c04000043400000000010000c404c05300c0c030040c403044000100000003000c000000000c4000340c4c01dd0410010030001000f000000c0004000c0c00000000000070000030005307040000000000c05001000001001030c0001140110000c3410c00c0c00100c0000c00d01303000000c01cd00005c004400000030cc00100c00c14400000117000c0000000000c0300000140300c00010000c000707c000000000d0c0c00010000001cd0004000000000c0041010100c0000c0130c4000f000c030004dc30740074040c00000c000010c001c000400001300001c00300c30303d0000100101000000f01d04c070f07001340400c011c01000030000c03300004010440000000010001010310430003c30c0d0304000110000303300403c00500140c30000c100000141300004d31000010000000100000710c040003000003000031000f0c00000c005400c04f0100100000f300000304030400c050c00cc0d0c0301300454c433004c00044000100740c3c000503400040cc4113000003c3030040000001000c000c0014000001c30c10c3040c0310100d040100c0004c0000004501001000c004000043400cc000000034c000cc30f30c05cc71c00700000000004c000000c33100034313c000031000401c007400000cc031110004004303030300000100c004000330ccc003c00000030000000c00040001c0000d01030c34001400000c0c04100300014300000000003c00000400000000c37003c3100040c040000004000c00010404000c000f003030011110030000cc1c00c0400003000010100301100010030007300c00c000c0743d0c0c400c3300f000330c700c00000001300c000301000c00000003174000000000000000003c000101c0030044c34f0000c4000040000cc00700011100300c45cc00010000001010000000000f00400030cfc40400000000000000000000c0000000000003003d00400400c000cc0f3000030340f400000000311400030400000300130000400001444003100740040c05054c40c7430000400004400c000000000c01000004000c0010000710300000000cc31304000000000c0047300100007c00000700c10cc0000430070143004c131000c040100dd00000000040000c0007000c000001000100407c00030037053000000c0400050030000cd0c0cc400c370000100001c0030f00010400010c00f4c0100c0033c0c00c003cd0000170df1c430c000c000030003000001340040c07010cc41100000400000010440c00c30000100004f003000000103000040c7c53000000;
rom_uints[3] = 8192'h104000c000004040000010010000301040031000300130000330100000c0041001d0303000300300003000701000c00400003010c00000f100003030300000000040000000c000013000040030000000003040c10330f0dc040000000000c00010c0c4101001c00000000400000000010001304c0c30100000c000000000000050004000000000000100101000010030100000000001003010100c000000000000000001033000000000000000003c003300300000040000301000000c00c00300103030000030003070000c000000110010031040d050000c100030403010c0100000c003310000003001f0040000001010c01010000c0000400000000100000010100110100030030000c00000003004703300303300000310c100000013100001000003000000330030100c331000303070000c3030300000c03c00d0000013000c003430000040007030400001300010000000000000d00000103300400010401400d000d300104044d0003c000000044010f0004001334000c0000000304000ccc01000001710c0000050040010000030330000000000010330000000c001f0100000101030000000030030000300705007001010000011c03010c0c03000d4c7043000c1c000000000c0000300d01500000003400000d010000000100c3100331040033003fc03000000300040300030400070003c0c0000c003004014111000d0300000000040000010000033001030003000400c00003140400000404030310030c00c0000000000700000000000700001000000300000000000000000004000000000004010c03031c00030300000001000700001104300100304401030000030300003011c300000000010c00000430034f0030001d0000000000c000004c0300000f000f31000000500c00051c3c03c0050000d00c000c000000401303000001c003011c000734000075000cc11000100003c3003c00c10000000c000000000000010003000300040003000001300000000130000c0f00000303000001000f0000000003014c30c00001000403c10c000f0000000104000000103000000001070004030000400001030300040300440003040401004004030000000f0000030400040000000400000c0000000001000303000403001c0704050000100004030100010000004310000030000300001d330000010c100000000010010000000f000000000300053c030004000000440000000c0cf00003000000074003000000003000010c030000000d3000c40f001c0c03000310030441c0004303003c00441c0103000c0005030003c00004041043000d3003000100030000000100000c0330030303000c0010c300440000030300000100100300010d04c1c000000000c30000000033030004000c030c43000000000d000001004000000001;
rom_uints[4] = 8192'hc00000000000003300500c04040c0000c00000430001000000c0c00c0040c000000044410000000000000400400000c0000000404000cc400000000000000000040001c00000000400004c34100011000000c0104c51000000004040004010000400000030000000003c000000000000140001c001040000001000130c00000400c040000c0000100000000c30010000c00000000000300c0004430350000c0c00040000c0340030c0103004300000d0040c0000000040100000010010000c4004000c00000c00003000001000005440004dc0000000000004340c00430000004c00001450000300040000100110c01cc003001c00000000000000000000000000001c0010005c00131000000030010005d0000c0cf1030c004000000400000004c000030070000401ccc0003c0000000030c00000cc0000000000f004f44000c0003000030d000000000cc410000004d040000040c001c410407d000c00000540007c0c000030c0001000000034000004000c0000d4c03004000030000000000c40000c107000001000000000001440c0000000000030000c4740000000300004100000030000c00c000c0000c0030000cc00010030000c300010400040040c30000c001000405007003000400cc000004000000000c00000700030c0c0fc00000003010010fccc0d10c0000000c40c4000cd000000000030000000c00104c00000001000000100040000001c0c4014003000cc3004000030000115f000300004c000c0ccc0000000104c44440c0c40104000000c100000f030000440004c400c00000000000000cc0300c00000000000000000000c0c01040000040000c4040c000000000000100c4000c00c051000000c0000000404404c004000f0c0c0000044000000000000c000000403005c000033c00010300000000c000c000c40000000300c003000410c0000c0000000000000400c000000100000404000c00005300000000000000000040000000130300400c000001040040000000010000004000f4c04103000000000107000041000000c00d0041000000000000c0cc0c000040c00001c000010000030001c00c000c000000cc0000004000c00c04000410040000004c0300000000010c3000003000031304004d0c00c0000000c000f0c000c4040c3404000000040c0001000c0003c0c044004300c101c30400000000000100c073000000c0044000000300000000c0030000001000000c000c0000000c4303303c0000c0c0c00000000000040303000f04000000003040cc0c4003010c000404301000000c000c40000000000d001000000004000000000c00000cc00c0000c010c0000030430444c00000004000000000000c000000000403000000010c0304000c4000f0000c10004c400000000000000000010c00c0c03000000000;
rom_uints[5] = 8192'h1000003c3d400c0114400005001c0000004004003cc10030073f40001100000000000c00370000010300c0c00000cc0004100c0000400400400000000001010573c0f404040004000005cc41004c040040010d0000040000470410000d04c700031c00410c0100300c340c0000010c1001000f0043440330c1c57000000000c130104000dc011cc00c00400000c71c000004c000000c004c00010c000440000000014c00c0300000cc1c000c1100007000003000c00c00030003000100043c000004400c00000c0000000010001100011c000000000c00c41100c003cf000141000001c0c000000c00001d0c4000000000c10100c400000400010000010103010001030140403034011000000000000cc4c003c403000043140001140f101000000c00c440f741c003c000040040000003334d000300003040c000010403000c0fff0f0000c00073500c000001001c3100c1000000010304d0004c37c100c0c5400c00000000010d070000100c0007000c37350000340300035c43100400c4011c04000500000c004f00c0400074cf0000000000003700071000000000000000010004000000400001003007030d0c330040c0034435c0300d0100001d000c0c5d100000040044c10c4000070000034000c010300c401d00030d003c04334c4001000c00400c0304010000100c0051c3000d0700d000001f300304003044cd00000001c07c030000100c000304003d070003400f000040c40d00d004004130000cc000000000c500000010414030444040700001c11000c0f0c00000000040300004c000003100c00104c1113000000d0104000c000c0100070c0c0040300300000c0000c10001030104c00000340001007000000d3000100133004040000005001001400c000c0000400000000004400004c0000031c0000000447340c0c040c00000000c0000040050000304f04340c3404c03000030c00017004104001c030001000000c00cc0001000001000c4cc3700770301000c034000cc04c001001000004001000400000000000c0100000004304d330300000000700c5c400410000c300010c30c001d00034000000c00300400053700003f00c4c103000010c440000001c00311c030413c000c00c14c000cc0440077c00004000fc003001c5c0151404000f4c300c440000c010040034500000c00000034340c0000000300004004c10c001000c0104c000013c0000000040c40010004400d030000f300f1000000000000000340340100000010010400070000000300400cc0070400d0c001040c0330400c10cc00000100033000000010004c00003400cc00c00000000c10000004c40040000103400001ccdd010c0000000040000404c005000c0007004130c0400001000c000003c00034c3400070c00c000c00c403c430000c00000040;
rom_uints[6] = 8192'h30000000000c000430400100d04000050c0030000004404000005d0000c00400c000000c000c001c0010000c04004c0400c00130d0400c3000001040c10001c00c000000000010c3300c003010400003c000000fd1f000000cc000400300cc000cc03000000000000050010c0c004403011034500300f450004c001300c0000100c0c4c040000100d04000001040100000d04400004000001000c000c03c00000c004000000300000330c1000000100000300340000c0c3dc00000c000cd00000000000000c0003c001040f1c04003341d0040100030c000040c040c004400c00000c00000400000003040014400003000100c0c00000000030000000c00044d0430000d00000c1f100c0000400000000d00401000404000000430000140100037000c00040d030700000d000c000c00f00d000100003001300000400000140c101dc0010cc40d003003034c0000000030100000140013000c00003007000440000ccc4c0150100300d001000044040c003410007d03300c00c03000d000300c4c000010c0301c01c0010400000010f0001440047fcc000d000700044130000003c100001c000040000c00300010c110330c0400d000003000c030000330401cc00c000000f01000000000500000c400010010c0400d00000000c7400000470000301000c0c04000030000010003001000cc0cc0f010103400c003f1000000031c00000000103110000000300ff3c0c0103cc30400004044f000001011000000c000000000300000400c1c01000000000043000000000000000cc00c00000c000c0d00001c0c00003130c0000010300000100000300000100c00404013c0000441f00005503031100450300c030000300c0000300000300c501410f00000300030c030000010000c00c00040301c703003c0400004000000c01001000000000c0c0000040000c00000043c140c07f000000000000d050400000c040000f00000000c00400030000000103000100c000400300010101473c005030000000000140000000100000c0303c000030010344000000000004cf00c13310004300410100110000c00001c00044400c0104000c30000d000010000001000003000c00c0100d00440000c0004000cc000000700000c1c1000144010345110004401000410000400100000c0d10100c00000c0004c00040001404040000000c30c00104c1030c000030030000c4000000100000c00344c044fcd40003000dcc000015d401030040000d0004d044c000400301c10000001000000007c01044000001cccc003c0000cc000030c031c0c03400c30100c1000001c100000000003100000000010003c401000001000f050c013000000000040010c1114c00470dc0000100c0000300040000c0030000007400000040c0007003c1c000d00f00000000;
rom_uints[7] = 8192'h4000000005c0000c000d300000f41c040000cc0c30000000d03430740c04000030c303001c00001c000c0c00003000001c000cdc00400010c01c004400000004000000140c000000000c00300050000c300440000044c040d030000030c0c4000000004000c040004c04304003000c0030ccc000c004c0000001c070040000c0c00c001000000c003000c40000001000d400000000000010103000000c040c000000000000001000030010c400000000001400003c0003d000000040400000000d00007c00c0013c40000000004f00c0c0000000f500000000f00004401000000100000004000c3070400040000000c00c0c00000000000400000c040c0034500c0000010000400d00000070330010000000400000c700050c0c0c0040400c00003000000c000c0c140000000000c3d010c040345003000104303043d4000000003c3000f04000030c000c70001c1c00040010040005c00000011000401000000000000f3c000400410c0040403030000043000001000c01c0000400003400c00000c00040000040000000c000143000000000c000c00010103c40f0040014005cd0300dc0004000000103000c70303000103401c40000c40000000c0030300040000000000c0c00f00000c0c000000c00000000301400000300030140c400010100c01000c0c400100000040c0040000400030000000c3000000000003040d01c00c4100030500044400410040c00cc00d000cc10400000001040c4000000004000303010000c4000040000c100c040500c0040003c00c00c3000c000f0044004104043001c0000740cc00000000040000c000000000000d000030004400000000000000cc01000000001000000000c00c40c004040304c000000300004000030301c0000c00404c400400010000c340430c000cc003000310000c500300303c0044c70000c00d4000003f00130040040000c30001c0c4c000c300000000004000001000000c00000300040000400407400101c30004000040340000040000c004040c30c0000c00c000c0000001000d0c43030000000300045001c0000001000000000340c0430c0100c00000000f0041000000000c0000c0004000c00735000000000004004034430d00000001c0c00c430300c000030c0000c10d003004040c000c03044c0000000001000000100000004000000000147000030000c000000003c000000000c7000103400040404010c000c30c0011c0400cc0004005000c000dc0000000010004c703c0000040000300004003000000c0010300000004400c0c040000c1040040c0400000000005000300300c0000c0030001000dc000004040400d4040c30001c70004c000c0000004c004000c43cc000000004405000000000000c0000000404000007cc000400007000001030300030c010000000;
rom_uints[8] = 8192'h44000030010300000000010003004403000001053000c000000000000071000003001000c0000d0400000300030330040c1c01140304040101000030000c00010040700d00004100010000000d04100010000704000000c003000000051001000f00100340c0000404000000000f00500000c0044c10000101010700c1300103c30cc000000000050000010004010000000000000170140000000033000303100300000000033140000000440101000f4c0000000300000f000001001000c10c1c100000000140070001c0c00014010c000000014fc0000f030140034000030000000300030000054000000c0100310011010f10000000000000400000040000570c00110014015300004c00000400c30000040030030cd0000d7033c003100034c00103000400400001000043c030004d00c3010400013000000000001001004d4300000030043313011100000003300033400f40d100133300400400300303ccc0030003010301100043004000040007013001043301400000300000c0003301300110c0400001400103000c0314000004300000000003000c0d430000000c0140000c0003000001044000000104c000000500050000f000000003000d034113001d30000710000000004000000113000000030130c010c0430030000100110000400d000301c000010f00010704400003000303000005000040000003fc0000001301000170000d0c00c1c40d030f00c00000000004000cc0d0074300c3054710000300003000c33303010140110fc010040100004173000300000000000400c3300001000034000300014000000501000103c300000050400001314070000000000140003cc00000000400000004110300000c0c001103100100c003000000303c00000000040c0c3f710301000104404140cc010001000000030001040040300000000004000340c000c000c000000c43000310d41000d000000003030d0101000000030300001000000101000000040001000f04c000040000000000000000050300c0004300030303001000c000403310000000c1c0400f500000000001000c04010701000004030003010c0df31403340400030000000c0000040c30000c01000300000000000000013000000000030400000004070003d003004100130c400000c3000003c0031441003c030010000400000103cc000c0043000000004001030000030d000403d0000030000000003305510303000c000000300700004101f00300000000043c000303030c00000034000103000050c301000003000303003000050000300134c03000c000400004000104004000100c110440000031000001c304c300030d0013000003001003000040000041000c0040000dc000300000040045c71000000303c0100103000340000d00017000c30c0300000;
rom_uints[9] = 8192'h70000c0070004c01004100030c0041f03003000007400005430004004300010100c00000401100300000c0c130034031000c101000003300000314000000010033014000000100000000c00003cd0031c15300040110004140c1c100fd710003c300040000c00000000110c400000000d0130140000030004003010c0400c0100040c000c0005340c0010100004040030000000c003000000000010413000003c00000000000000000004110000011000040000400000000400000404000030c0d030000000030c1000000100f4000030000c303c3000c0fc11d010c400000000000cc00003000000303070144743003c343c00040030000c300000000000100000000010030000ccc00000700010007004f4003300000104030c4030003400100000103300001101001c011000013400000011341c00000c00000000000033100c00004114000000007c01000000030001300003c0300300cc301010001007010000fc00304100c7100030300c1c03044c00104110403310001000141000301c00c0d400000434330000000000043000130000000d00c00003400000300000d410000c00000440003c000cdd000c00000403c00013000c0001401330003c3f0000404003000300c03000d000000000140c00003c07300000000033053100000054c330c1003f00c4300000030c1010000013301000000c04000130cc01000003000c034c0034300c30000c10304d00f00000000000000000370001000030d403000c000c0000000040400000000000d3f00000330000000030000c00d00d400c000000007000000004000040300c000303000030c001c3100000c0000300300400000000030400000001cc00041004003c0100003000000030000303351010013000000000000c0d010030000c001dd00c00000d3301003003c1000000030000310010fd0311103cc3130300100440030000300c0c00000404000c300100000010000100100010000001000c001000000033100000c0040000044010030c00000000000f0c040037c470003c030000101c04000004000000c00c0333400000000300311030d30000000010300010c300000170030000000040300f33cc10004000300030030130c430000c043033000c0c00000100000c0033c00003000037030c000014007000411c01030400000000c000301c00401000000000003d30f4003d0100c1000000303c007d001d500010000000300130000000c0001007000c0004400000000000000000000000010000000c00004c00000041000000004010cf000c4000000035030004cc01303000000f4000001c0000000000303030031040101d03000000003c003c0d040033c0003300000000110c010000000000fc301c0014340000000034d00c100c3300000c00500c04000044100000000c4000;
rom_uints[10] = 8192'h300010000030400c0034101c34100040c0c00004004c040000d03004000c0000000c3cd00cc000000c0000100c00303cd000c0f00010040004000010000010003000001000440000040000c00c00000100500040133001301070001000cc00143070001cc040000c0100c04000003000004000c04000047c00c030300000100000d0001100c0004030140000000000000c301000000000f0f03000001c4000000000004000000c3040300000000000340030100000100040000000000c100010303410c000100c00007000700430137000f03c000001c01400140000d4c0000c000c00c010cccc000000003c40d0000030000470000000000000000030300000000c0000300cff0050300c0040d000400c00001c1cf01c0000503074041c304000500000000c00000001104000cc1050003404007000000000005c30400400003c0c301c3c540400c0000c104400003c00f00400c0c07400c10040f0103c300000003000000400000010c405000000100000c000004010000010c00000000c14000004c00c0000000010000c0c000000c00000000c00041030ccc0140044000030d04000303000c03000c0c030004000000000011004400410500014004000003c4000005000010030ccc0100c00000030c0c0000030143c003c0000c01000030404000c400030d000f0000040f0000050f00cc010c0c00000000000300c1000c0c00010cc04d070003c300000740004c0300400f03000fcc430000400c00040000c0000c03d0070001030f00c40300040300000000404404000d0003000105000003004d01000c000400000000030001010f000000c00403c3130dc0030000010100000f400c0000000c010000c000030f0004004c0001c0040c100000030c010000000000400c03050c000000000c0400c003000000050000430043000000c0c00301700000000043c0c10c0000000cc00300000400010f00010000000440cd1c0cc000000cc00101c0000001000cc001000c110403000004000f0000cc00c0000003c0400000000c000000004103000101c4cd000c000101030c000c0300000000c003c0c00507c000400003000003c00c400001c00403c00000000c03401dc0c00000000500000000400000c00c0000000c0000330c00ccc0004c00c0000000000000050c00000001040c03010400c00000000c1001000300400300000003000447000c01030c00c00004400000000000040400010c00c00003004001010700010000000001030c0000d0010403004001014004c4000440400704ccc00301cc00000000030004000cc30000040fc00c010300000301c00c0300030043000005100430c0f0c041010000004031000003010300040000d000400303004001000000c0cc01000100030000cc030f000c000000c00300c0cc00c00d000300000;
rom_uints[11] = 8192'h3430000000cc070000000000000000403c0000051c03050000003000000c00000003014033000000400000000000035000000000c0000010c000040000000000000000330f340003000000000000001010000003000003003110004c00c01000000c30030003000310001003000100400001400000030001000003000001003030000d040003000030000000000000000004000000001001030000000334001c0003701000000c0400000000000003c00000030000000000100000000c0000c003100000000001c00c1c00050000000300010c300044000003000000100000000000010000003000000000f300030000000100c3010100c0300000000000000f04000001000cc0011000001000000000005c400c000300000300000000030c0000000c00000000000000030000000303011000000000000000000001c0300000000000000003c3000300000c040000004300300f0000c0005000f000000403310000c0000000000073100010000003d0000003300004400c100c03000c00000c0001000000003001000000000f04100d0000000000000000110c4430c0000100000450000003000000000010000000000000c00f000010000300004000c300000430014050010400000000001c03000000030000010000cc010000000000000000040003005003000000010000040010c000000300000100001000034c0000000000040001440010000f00000c00000000000100010301000000010c000000cc0c000000400c00030001030000000000030c0000001000001000000311003010000001030400400000034000c4400000010000000003000003100400110033000030030331000000000000100c0010004000004000004404030000000000000300300000000000300000000000043000300040300030010000000100030000000c000000c3000000ddc1c00c00000010000300000100000d00000000000000010330030300003001300000010100000000040c03010000000000300c4000000000000003311c4000000100000000000c001000010003010000000000010000010044000003c000c0000010000c000000010000004000000c0053030003000000000300000430300100300100000000000000000000330000100010000113c0130100000000c00c0000040c00014010100004030004010100130c0500035c0000c0c000000000001000000000010030010f0c0003040001001000000100030000000000100300d0c0000000100004000300103004003003000d005000730100000004030d73000300030c01300100000c0000000000000c0010000c00000010000000000f0300000000000003000000000000000000100003000000000030010300000000000001c4000000001c003100030000003000000f4000000500000000;
rom_uints[12] = 8192'h10000000cfd000000c000030104000c0c00c0000c4000d000000040cc0cc0c40cf340010010c00c00c0c000101000c0c00100040000c040345c00c100c0000000400c00d400c00000c00c303c300000c0040000000100c00c3000440100001000044004340000c000c000000040000000c0000400c000300001cc00c100000000000040000c00000000000003300c00d000000300000000304400c003c0003370d01cd0000cc000000004000003c000c00000c0000c0c0000004001cc000400000443c4c0000740000410000000050001000c0040000330000004c300c0c00340400000001c1c000c3000050010c0c430003c0000000004c0000040000000033000400003400000c1000004c000c1c0000401c040c000040040f00040c0000400070030000140c050040003000000000000000000c000c000000c000f00c4030c3030000004000d01000304c0c00000d00000c00001003400c0440000c0c400010003400f40000000410000003d00c03000010100c0100000100000000c0c34c0000cf04000c010400c00300040000c45c000ccc4000f0000c40000000000000000c0000c000c00440300300044000cc00004400d003000000000c1c0000c74cc00000000010000f04004000c030004000000000c0001cc700c010c000000cc0000000040c1c0c04c0000c0cc00c00c40fc400400400030c00400000104cd004000000c0304c0000010310000000004c73040040000501c0001001010000c310000000100001003c00003010cc00d4004013cc00001ccc00c0c3100003000c00400041000000400400c4000c00cc00000100410004003000000000000401cf00500000001c0c00c40000030000000000000c0001001c10030104000040000000000c0001cc000030000004010000000000f000c00f04000000c30000103440000100000c1000004c000430340300c003c00c00030301000d00000004000003030000100003000007000000300030000000134041030010c400000c014c041100300000000000000000000c0c0000000100000cc0030000000010004100007000f00004c304400045000000400000000004001c40000c000400040004000000000100000000000400c00400d10404cc010000000300034c000000700c000c0000d00000070ccc00004c4c000000000000330c000c5001300000c740000001140000000000000c00c0700c00440fcc0040101d00004c000c043c0c0070000c4f000c40c0000000700c0000004000c003300c0000c00c4000000c000c400000000c0030c0001130451000003c001000000000000030000c00c0000000000100011000000047001f0300000040001000004000400401000000300030000704400011500040c400400000000c00f00000000000000000c000c40c0c00000000100000;
rom_uints[13] = 8192'h51c00000cc0300000300c00100404dc041003f4000f00040f0000010000000000000540000000000c30003f0000101000040010340000f000000000300010000400000000300000000c000f000010001c1030c03c11110f4ccc0000c000c430fc010c70001001000c0d001c0c4004751313dc04050c04700c00040ccc14010fdd41300000000400033c00003040300c0000000000c50004010000000c000010100100000d0000c004c0000434000030000c7000000111300c00001cc00000c104000100500f013c4300000000c40014000dd00c30cc4c44041400470440000c040000000c0100300040031400c1130003c000030c000000000c000000000d040100004404c01300340000cf000007004700100f333c00000c0004030000030c044450000000fc34d400c10c300d00000c004104000c30000c04000400000401404034100343c0000004013041040510114c04c00c1f001000004d00430000400c0004044c10cc100030000c00030c70000cccfc10103004000c00003c000c000c01000c30c41c4011000000140000000000400c300070040c010f0c4000000003c00c04d04000c0400000c0040110000c0c01000741000c00000004000c03330c101c0000000d00010003040000040c0000010c00000404000110003c0000040030010c03040f4cf113000c3c000000f0041c0c031000c000100403f0000000c00c00334c00040000000c00040c0c0f0d00003c40003d000010300f4cdd300cc0c3100004001000000c430000043d00000000000000143c00110000000c0030c03000000037000c0c0c000004000000000000400404000000c41000000140030f1c010300100000cc011c000400004c003137000004004000000001003c10000c04103100000d000030004040c01c0c3404100000100cd000300c0c00c30000c0dc00000c1074003010100441030c00c0000000040c07030003c70100004c0c0c000000000c000c11040000004c00000c00300140000c0300000014000cc00000000000c00000000401000000000cc0000000100000000c0001c0071000100c000000000304d03c1000004004000100503000000000c0050000c00100d03c00000000000040010c00434400003010000000303c0c10000d10000703f0000010000000401c051000030f0013c40cc0300000000c04000400dd00100004d00c000c3030300410000041000003000c000030c0000300034113000004100cc0004000c0d40cc0000000000000c050104010004000001cc400034005030000000c10000d100c00300030000000141c00000001d03114000030040030000c00000c4c004c0c0400300cc00000000c00000000000c400004100400003000040c000c00300cf00c30010c000000304300000c053000cc0000010010d00000300000000;
rom_uints[14] = 8192'h4000414d0040c50400004100c01403000004050300000cdc000040010d0040000007c0100000007300c00343040c0c004cccc3000000c000c004430070000000010300000000100001004300014704000c00c04070c54c00f000000003c40d00d300400030400c0300c041030100000400000c30400103010000400500000d000c0000030c01000000c100c01450001300c000430300000100c400c0304010000000000c000c0000000500300313000033000000040c0100000c400f0040000c0cc00c00c010001f0001c0004011000c0d3300c0c00cc30dc0001c440001c04000000171000000000030000c040000010001000400c000000cc00001000143c00c00033000014003300c0c03000000074c0410000c400043010403430700400c030070030303000344300403030cc01000001c400700cc000dc040c40040c00fc03d400000000f01001000c00300cdc0400c310c33c10400c000000313004000000f31c300000000100000401d0400004340000003001000003403000040f400c4c0001000c4070000000c0c4040000003c400400300000000730004c0005041d0000400040cc0c0c40300000c0030010000000040c004000100000c000f004100040300c4400400000000c00c00c3300000000100f100c4000c00000000010004010c0000030400c740000000004040000300030c00c000000400cc00400dd00c3c0f0f0010000100503d00c401300c0050341140c0070c300ccd0c01dc0000000000c00c0703004000400c00c44c4c0d401400000dc0c1070100003c004c401c030c00cc000c430001003040004c10040c030c00030307030300004000040ccc4000c0c00c0000041430014001000001c0c4000d0003fd0003c0f00103000004000103000005030f00fc0000c04f00300c10f40c040c3c0000c000330010000c0040cf40c40f010c00c440c403000c05c00d00000c1000477040030000130440c10000c0010007400003000000034300d0c001004cc400000000404c00cc00c05f043007000000010c30000000001003c103110c00004000007d0cc0000d0c0000c10f000c000300040100004171010c00000010cc0c00000c40000030015740030c000101004c000000040450400000030004c00500750c1010c0000350430330000004000d0000000000000000c0030c0013001c000000000010f1c000c04cc000c000003c00001c000000400440c04f0c34100510400000ccc04c0cc0000c0000000c0000003040003c3c40030f0c03001f0000010c0f1000c400004300000d4303000000000140000c003400030000000004440000000000040cc0300d00000000400400030000c001000000c4004000430000000014cc30000c0040000c00000000c4015c4000004cc10cc000047cf000010c400000d0000c0300;
rom_uints[15] = 8192'h1c0d000000000c000100c50d030c0c043100c00040040000000d0000030043141010000500c30000c000010001001404000c03070000030c000400000c010c00300000040c00040700000314c4001014100c0000040c0010341c00c1c0070c4c0c00040c00100104003c00000014040c1710401cf03110000004040444f00000005030000001c410070c000150000400050c01000004140445040000000000c030d30400003000400400000043c0000330003dfc0030000000000414403410301c170000c0000004c00300000c0c0404040313000050073c100050f5400c0c0c000000000000dc0c001004340d000100440c0014100c0400011c30c0000c040004000dc00400070000000c00300c003c310c54003d010c0000030044010401300410100000f0000030013c3c30000300000010040c000d044c0cc000041400341400001700010c3030040c0f0000c300410400030c007000100f0004000400cc0403004000003430010403cd3000000d00043000fc711000030104400400cd3000f0170c0000343000044400310004c001000c00d0000000cfd400f000100c300401000c101414c007540c0ccc0f3c00cc3c03340104144000050400000004000000073c000404000000000c10000400100401000c00344014c0100c1c3400f10c040c410c00003c31030407310000f0c00d04030f100300c000000400001401130c7c7c00000104400000011c40001000d700000c0c04000405400f000c0000010100540400c014000c0300300404100c03070004000000001000dc0c00004d0000040c3c04100c0cf03045000444400000c300f0040cf00c10001c1004f30c14040000400400040c040031000c040000330c0c3c04030030000000414043c0c40c4700000014c04d0d0c0c1007140057000400000000d0000c0000d04f00c10d000c0414d4000c0c00543c0010014403040004000c00c300000030000004000304c4000c0000000c00000c303c00c000040cc00d0400040c010014d03c00101000043400003c1000c0130000300000c00c0c350000000001000400140051100c003000100d00310400300000040c0c00000001400c0c3d5400cc0cc4040000003700c41c033c0d00f40000003c010400030c300c010c00413c0c100c0000040d35c30700100c001040010007040000003c0030003c4000040c000000000c04040c000c0f040c000400003004000c010c0000f0000c1004000000070d00c13300100100c0000000000000000100c004000c30cc50300c30030304c00500000c010000c13400140c040410000c00004300c33003140000000000000000303c300c3d0d0c040d1403000030001fc00400001000000004010104405030d400c003040c103004010014000c30cc0043000000f0000031040403c40504c10030cc30;
rom_uints[16] = 8192'h4000c0000000c3314000340450035010c350004050c04cc400f0400010000000000c04400050001000000040f000433000000f5040c4454010000017500010c001001430c0c400c030010000400040f00030c0c04444000301404000100cf001334040c000004010c440c000033010301030c34043c0403000100000143007007051340007004c004400c0c0304040401010000000000100f000c000c144c00040f0c001000ccc50000001404010c0c0f0040000000010f0000000c001f0000010300000000c4000c00050c3c410cd000000d0c040d000001f0c0000c0c00040c0404000001450c054000030033030c01040500050500004d000005000000400f0c0cc410c3c5041310000050350c0000030004010000000f0311ccc3000c13000ff0000534c01f000c400f07000f3c400400000c004c0c0c004c054cc10700040c010504000c05030400040f000300030101f0000500001f3004014c03030510300304c50000050c1f0100c004000f4510700c01034c0400000000c40c437400001c01003001c40f0c000f0000c3040c000c014300c30405c01c30000005004c0f1300400d0cc00000000004c51f044004000c400f10000c0c3034100100040400c7000000000000040400d3040c000c00000001c000310000c10100140c000c00043d00c0050300050000c0040f034000054c00030c0c00400c00c003030cf00c0c00c50f0c01340c000304c001040cf4000005000f40000004c404443c010f3000000c0100000003010004000c004f010004031c140c0400000400000c0c0f0f04000d0c0004000c100c0f00304c004d00000301700000000405041c00330c00054c0410c03000000400030c13000505050430010d030c0c04000001050c0f00cc000400130c04000c000c0000c403c017f50c3004040001c101040c00000c0404000c4c040dff440003040110030c1f000444007005030d030000000c000c000c0000000f054137000400000001000c03c0000fc00c03010c0504400c040500000c1f030c0000050400c0f00000050f0f0c040c0100400c0c0034040c05050710010c00054c01050d0f0c003041011f040444000c000c1c0c0f00040c00014c0105000c000503500445000000000004000f0441000400000303040c04004c1c0f000004040c01000c0000104400000f00030c0f000c1f00040000c0310010010c0050300003000c050c03000d0f000cc00c0c040c04000f0004000c0c4d0f00501c000007040104004c04040004050c00330000000c04000000c3000000430c00000334df30010c00000500040500430004cc000004000c0300000005000004010c030c40010c0f0300000000c400040000000100fc00300000c0700c004c0d0103c00cc000005330000000c5013c000444040c040f0500004530040c00;
rom_uints[17] = 8192'h70000300000734300000001c07000103c30503030407470000000100070130000300000c0cc3000031000100000000013701000400c00011010004000f0013010f01100300370130040003000000070c01104030000303011c00000301000d4000000303013f03034f011033000000000000003000330001000f0315000d000003110c0000030300010400004015030000050000000000003000070101030d00001d0400300100000c03000c0c0400040300030000030303050000003700010300040300030000030c0000000000000303010f0100400003030c03100000330100050300040003000c0300350333000c400104030100000000010003000c000c0410030113010411030400300f00000400c10000030303011000000400300c10031701000301700f0050033c3d040c430000000400030000010000040344030011000004003073000c00103007030004030133330003010711000d30000030010c0c00000c00000c0f1100030d0c0f010000300f0f01030d017003000313000004010000010000013c113003030303000400000000004d000100300000000000013300000033000001000d1400031c04031100010c41330000000130033300130d03000c07000003011c0100000c000401000311030f00030113070000030c000c00033700300300000001100010030300030000101c000f0c000301310003333100735300030100000c030c0c4700030130000011070001010014000f030f000004000303400001000131110d1000000033010303050030010c0000110003000000050c140005010003000c03030000133701000000030000000c000c04000300000000130303330500101000000010301330000130030c000000000100010c00000f0430000f010c030f0c030700144c001101cf314d03030301000f00000003030000000011034d0503c0010303c00400000010040003310300030001000c0c000100030040013f0f00000000030c03070d010f030303300005000000073000000105310dc004030501000000033403000c0d000000000c0403003000010c30000033040104001000040d030000030114304033000300001000000c00000c0030300033004c00000300031100000503004503003f010d1300110401003c3000130110000315000004030004010f0001c00c01314d1003000c0103030300050000033c000c00000c0001000d00004300400133300c0001000000013c0300000030030103000100300d010001030c010330000003010d04013014014c11070001030f013d0001000000000d000003000000000c3c00010000100000000404100010030d03c030040003f3000300000003000000000330440000030100301031070c00010007100300100c0001001003010000000c0000000c00000505000003;
rom_uints[18] = 8192'h44401070f015001010d103d100031d100303000000331000303000000100c000c0001c003c0000000000001c00c54c0f00000105030c4000031140000040000304c0c0030530001100044101c010c440c700305c40343033001c100101c40000d00c10300003004043000013003f0f00c004d00c03c0c3d003c5040c00704304401c00000300143040000341000101034430000031403040035000131c1c4f1004000000c3100003330c301050c07400000f0c0000c0c0000300010004001c401100050001c0100c01c041103014d0011c3000000400134410dc004000050010f00300c1004c3000114015303000100330301430000050400100404000001345c0030000340c01041013cc0040000003441c0003077fc0300c0034013c10100004c0000070001000440004103101530c0100c100455300040c40cc00c431c0c0403043400000c00310c3031440c5c014400003100d1000100001c00000000300c03030d300037000050040c0011c0000c00c304033000f011c1c00c3500010030151707000000000700000407435cf000013000400100130104004414c003000c003c5040010c300c300440f3000014000340305d50440c00407000c01034140c0cf0034000003000000007300000534d01003300c05d3030000001000003103110340101f00d3c070100000300000410c44100514000010340000305010000000000c0f151f340000c001c0c4000410c10c703400110004c0c1005f03d300c0404cc0010c00400000100cd1303c000100013011500030404c10030c105100030000103100003003050303001113030041040001c330c000c5400001c033435130c040c004000004d00570014301003100d00c334c430000004f0133040000c031140100100040030f00501c05000401001d30500000004000c301c4f0050173334004001300470441400310040034005d000040110070304034030303d030c1050000000040cf03030000000303171c05c0030c1400004330030c30300d0f0f000100c500c030007c030c001000000040004300313010101004100f0037000300300cd443301c0400101c000000c100040f005313430330014310010010001005003000c1003000d1003034f3003000c0000c43130c0040300011350040003500000000013c430004100fc3c4110f00030300107c30410403000000000050010044100450100003010000c000000017000000100005f00c370014330301331c4555000000000143c0030033740c00414130004c030c0010d170000043000330000cc0c1001000003000004c50c0c300c43c0310000040003007000301001010001403301700114011dd010033001d0000033000001343443411c00010400011000c30001333440030c0701c000030500000330300340c000c0344000c0000;
rom_uints[19] = 8192'h30030000014401c1c00000004001c3000300300c10070000003c4000000004000000000100cf300004011c013c000400f1c31c04ccf00300400004007000000370000000001000000000040c00301c03c00d00410f0010054c0c301303070300000d30000400000c000f0000000444010400350c401000030c040701000010703504000c1003404000400c010c04030304001c00000004400304c0000401010c30003400c0000070340330045d00000000000000000000050c0004051000003303d11f000c0030140c30000c3c003f01000040300f0004300c01c110301cc000001000051c00000103040004000404c03707031c104c0000000000003f3400300700c0d00000700f101000c00100000000c000110f03f4c000330410370704c0003d030000330304300c070304100301413000003100c3030100040004300c0005011040100c030003010000c543c7040130300c000300f4c40c0c030300000c04f00313030c310701113c31f003010030c0ff074005000000c004377000040c330c33cc070c0033cf04001c5000000c00300033000000404c00004f04c00c004005d40004400030000403000c1c05c0c3100c071c00071035140500000033110f0400cf1000c1000000c000c000400040f30cc00000c035c0000530000000400003000d0000100f00030000400004000f1000ff010f0d300c041004030d040d0030f00c000c0040003c041100004f000100c0300000003400c40c004d300f03f4013004000c0004000c3c03011403170000000004034300100100040300000100033f33000c10000403000500000100400331040433130410c30143000404cc01304f0030040040103010d00030001400000c1d0f5305410f400c030000000300040100c0030103050c404131103c0400000033103003000100040003000f0140043f000300c0000c4713010000400000d043c44c013c0f0041fc0044300135c000070070000f00304300014c0000040c00c43cc3050030f13330400f0001c001004300003c00050011000c0c3000000c0000050c1000c0300031011c0c000030001033313cc000310000100004000001100000000140000000040c05300c33cd0400430400000040303000000000400c0300d0000c0000030000070c00c0c70c053000340000c10100400130001c0400010040c00c4000040001100407004001000c41001001d100140c00c303400c00034f00010c0c34000c00010f3001403c00000404000c000004030401030c134d0c003001000000000043030104013000c0000cf300100c004000034c00000000c700000f001300134c00000c103330004c0c500704470400c0000000c0000c00c0040000040c03010300c0000c001f10000070030040c4400303000c0000000f4c003c31c000000000030cc00c1000;
rom_uints[20] = 8192'h1000000000003c003400030000001cc0cc0010003304130000000f000c3300010104000cc0c100c04041000f3000050c00000030000f0301f00700c013004c0004050013033000100300040474300c010030c30c3f1111003741010f00303000c00030004c0c300d100cc1000300f1000004433c0c1000fc0030013001000c4400c030000103003c0003c0000000000c0000000000000100c40110434004c00ccf000000000440c0000c0c00004000010400d000000400300030007000000004313000000000f0c54c000c0c030033cc00300130001400d731000005c030000030000000f00f0000000000470c03c504003000c000010430c0000001000000003400100105d1300300000001341d003f30100030004f000001457401070000004110000001000007001010000300f010000030f0dc0000c0500000c0cc040030c10030c0001f0c0000000c1000000500000003cfcc0173100d0333d0c3070005010440c0301f03130c00000cc000000500751f0000041c1c010fc0c003c003cf4037c00000001f43c0c10003c3000030010030300400000041c040430010003003f040c0004100c044000000100134040000c343f007040c0730004000c000f0c07000101000000c00313000010014004504000000f0303000f5010c0001137403001f40003041c4033104740300c4c3c10000100710700003040101030304c001400cc0030000c0000303004001001003300300cc0003441000c130c3c3c0c070d00000004001400010100043c100040c0040000045400c0003c10000003100000c0f00f00400c0003304000400cc00000004007403010700044000f100014000040c40c1c0300041010d05000c010c0c00c30c0c0cd04000300004054010000441f40f000304c0431c744001030000040001c100000005003d000311003f0010400000000030000f4c0c04010d00441000c001100403000000130040104000100400000c0000033000000c003004010c0100100c0401000000003c107c430c310000000333030000110053000400000100c0000030000000c003004300040c4f000c003410003430000c300000000030c403100300cc001041100004c000013100000400040000400004004cc0c00001030c04400000c0000c00f07310040004044400100550000000030000d4000000000c000f13000005c300000c4d0000040c004000c00001000000c007004000c000c00303403005404000000030000003001100040005c00f0030004300310000000003100000000f0001400041000c0001000f0c0100000000c00000000d00000000500f00040000cdc00000000c00000c110000f4400000c00000c070c0000000030000c00000000000303103000c000c010030c00004c0040c30cc00f0000003004000300000000030c0430f5000;
rom_uints[21] = 8192'hc000000300000400300c0103000413000400000000070000000300400c00000000c14c010000000000000040000030f1440000013100010c04000001010000400004051000c00c0c0001000330030100001103000040000000010100040100041400000040030f014301010000c03400000430030000040003000c0005104000300400000c000c00000001300000000000000000000010cc0c3c0000050c500040040000000c041004c3040010300c00000d0400000c00f0004000000000000000010c0000000c013c0000c1000c53000003000c4043010c001001051000070104000001000300000004cc0000003410070730000000000000100000040000100031003c3000000070000001c40004000c000f05000100000004000c03300300010000000f4000c10c1000015d00010404400000100100010000040410100000300000400101030100000000000c07000004c00c0300100040000f0101000000000105000040040001433000000005040000000403c004c0dc03010004010500000c000c70000c000c0000000c000d000005000100001c00000004c00f00000cc100d1000300000004c00100000300000f0000001011000100043043001700000303000400004004000000000400014001040404014f070000010140000c030050100007000300000300030004000001fc0c0c0000070500000c0004000c330103040000000c03000c0000040003004043000104300d000000073300040d0c03c00000000010000000131000000c00001000000301070401c50c0000010000440c0c0100000c000000043004000400030001003000000000130001000401000d00c00d007100070000000031040c00330000170151030000000000000003000c0410c40300000004000004040000000d1dc04400034300000304000001011401030c00001300000d1341000d0041001c010340000003303000003030000c440d0000000000011404010000000000000101010001000c00000c00000c3400000000000cc1010034000300000000000003000504700c003004000000040001c3040000000701000033000001000c0304040100000000c000010000c1000000010350c0000000040000000037040034000c40001105000400010000011c40000c000c100c0404030000010404071c0000105004400001c0c1010300000000000000004001001040000000000000000400140c1000000001300001000f0104040004140d07030004000000000000300001040100c00000c0100c40001c01003004010c000041030c00001000000f00001000100004c1000000000000000c00030000000005400400000c0000000000f000003000100003c000100000000301040140000040070c040034040050001400330c0003000000000c00000403040000000;
rom_uints[22] = 8192'h10000030000010100300000100000000003c00003030000030000030003400c0001010003000c10010100004000030004c30000000001000000000001000000000014400300000000000003100000000000000000000000103041c003000000000001c000070000000040030c10c10000040030004300000000000001000000c001c000000003000000000000000000104000100000010030c000010003010010001000000f00000000000040c0030000c000000000c0c000000000000000000000000100000000030000c0003145004c0f0000000000c3000000034c0000000000000003000000000000000300000000000500010000000000000000000000000100f0cf4c0001000001400000000050400c30100040010401001003000000003040000003000003700001010300041003031400010000000000c01400000300000000000040000000401000000000000000000001404340000003000300c00000030c00400000000c14400000000001000000101000030000c003030000000000c00000000000c00000010000400000000004000400003f0000100000001005000000000100000001004003001003000c01c003004000000000000001033000c00000c0000100003000030000000000010000cc30410000100000000300d00000cc000000c0300c0cc0000000000100000003010000030300000300000003000031000040000000000000000000000000000cc1000000c0000010000033010000000340400001010030013000010040c0000001430000044040000004000000030000000000030000101000000010000300010050300000000000000003400300000300400013004c0400000000cc00c005030000010000000000004000000000400000000000000300c0000103000c000001443001000000000000400100010004000000000300314003f004000f0000000001030300700c01000c004003300000000000000000000300000000000000004004100040000003d00100c00300000f00000c0000030300000000c000cc003030003010000004000000500000000000000000010000000000000000c00300000400000000400000010000000c00000000000000001003400000010003000100040000000010c00040c0000001010003000000c0000000c0000040074000040300000007000004c0000000000000005040000000c010c30c00000010010000000500000000100000000000030300010001000000c000000340000100330c03000000440000300300c500000004000000000001000000000043c0000000030000004000c0000000000000033000000c040000dc4c0000000000c110003000030c00000004300340000000000000000f040000000000000001c30000c000404000000000030000000000c0c0000;
rom_uints[23] = 8192'h40c00c0040000000000100004000c000000000404000400400400c000000c0040000c01000000000007004000400000f7030000043003004c00000045100000000004000000000000c000000030014c4000400c0000100000000c0000000c440c03000300c0000000000c4000000c00010c0000000000004000c000300000040c70c00000000400c00000000400010000000004000003c40c000000000004000000000000000134000000040040000c000c000000001000001040000c3000400000004000000000400c040003000040340c00000000000c00d3000c00000000c000400400040000000c000c703fcc00000000c000f00c0000000000000000040c3c40000c0100000c00000000000000403c000000000cc0400000000040c000c00000000000c0003c0000000300000f400000000004400000400000c1c0000000040004c0040c000300000000444000013000000c4001000004040c430040c000000000000000c000000000030003000000030003003000c3000c00c0000f1000000050404f10000c3340004330004c40000000000000000000040005000c0000000000000000400c0004000004c00000c0000004004c00000003000000400000c000040000000400000000c4000000004c00c004400104c000c0c000000004000c00040000040044000100000000000040010c040000000040000004000c00c00000c0c00d40030004cc004000100c04c000c000000c40cd000300c0000c50000c030001000f0c0000000000000f0000000400000f0100c3030c100000000403000c000000000c00010700000400001007000000000c400c0000000c0000cc100000000c030000000000005000c00004c01000100f04000000c4000cc0c0000c000100000000000000100004c03100004c0404004000030004d3400c000000c03c000000001cc400040000c004c3c00403044000040000404000000c000000d040014000000c0000c0c0000c0c0150c0004c4000000000c0000000f004c00000c00300004cc0000000c000c00c000030004043000000c00000000c01000f0000c0000001c00c00000000000000c0170000000144c00000000000000c00c04040015000000c0000c0c00004c00000000000474f00040c0000c0030003c0000c400c004000000000c00004c004000004010c0000004000cd40440300000007000003000003004000000c0000000004c00000107000000f130130000c00000300000003000000000004000f004000000000d00000000c000041000300c070000300c000000c0030004100040000c00000c00c400004400000000050000100000004010000000030d0030d04c00000000000c000000000000c400004003000100000000000010000000001010000c0000400400004000003c1000f0000000010000;
rom_uints[24] = 8192'hcdcc0000130050100400000334004c5000c5000001104000c1c300000c03541047400c0c0000445354000044000000004c0000c4400100030404c400c0c403c00c0c00c0000013cf0000400c30c00c0cc140c404f00010001403500c0f00c4500c000000400500fc0c1054000143010703c000130401000001000c00000140000000000403c000040000400c0000401000000000c0404030041c03c50003010c000f000000040000004007300c0400000000004000400004000000c00c4400004003c10040000c00000141300040404300430003cc40030100000000400000000300000000300d000040010c000400300044000000000c5000000300c04441c73c00cc00000c350053000c3004400004000c041104101c004dc00c000030000c000000000c000c04040000c4050031c03000c00c010000cc0074000c3c0000c0000000033c0000c0000130004c0000cc440000000000c0100000c000003044c0000000000d001400000110c000070000310100c0c740000004000300400000005043000000040001703400510003000c0003000c01431000c0f004c0144c00400000010c04ccc400403c040100000c0c0f040004000c3100010c140c0c03c40d000150000430000c0000050340000013001300400f103400c040004050000000005f07040c040035000400c700c1000c1000400c01040c0030c3004030043c00430040440c0c010c41005c000070050d10004003000440003304410c400403330f4003000000300fc00400110040c7000400000303f00040c00c00400104030100350c000004300000000000c400500cc0000040070c000c0c03c03c000c0454c0d001000000001000000c10c10c0040000103000cf7100c004000c400c0d400000c010300c030c030c0000003c00cf4000504000000c00140c30040000cc00d000010030c4004030040d44c3001000fcc003301040440dc04000c0414010c004000030300c00000040c0c0003030400000c101400010dc400c100000003000004040410000100003030004004000cc3070000c00c4c0003cccd000503c4000101000ccc040c00000d00033d00440000c00000000000c000c00c444c40c00000300000000c0400c00000000404d007541304000000000404000000040d10040007000401044c3c0c0d0150300430c0000400c0040ccc00010d4000000000000000f000c3110000c0000cc0040c00400443000000c3400c30003400ff00051400000430c0000c300400000c40034000c0000c30030030010c000000000000000c0000400400050c00500c03000c400c30f00c4500000040000000cc0000004c71054c0103c0004c0000040000400c00040330033cc000000c00300150000000c40043041000c0000340311000cc000000000c00c004c0000000000c0;
rom_uints[25] = 8192'h400300100c3d33c0000000c000000001040000d34c14400000f40000743000000000011000f000344010001f100047c031304100104c33dc000103001000100c300c043000303001000000c40001001000035004000300470c0cc300010d00d000541c00000c0010040c11003415070000003000fc00444c00003000000100040000401400003104000000400000000c010000000005100d0000c4c00010101000100c0c00c01c0400300400010004c000000400013c100d0034000704000c0001000c00000c013001d4003400035c10004300000044003cd00c10c014d0003000000047c030000001000340dd340c00440400100000000c0c0c0cfc0000007c500c0ccc7c10140d0c0000030410c443fd000003cc300000471401304340141004400000c0301044cc01fc0300c00c000100047010cc100003040f040701103400300c070400000030000030004000004cc000000c00010d001401000400f0cc10140500310400330430f00d0003000400100c30c030043100000000000400c4747000cc3cc0f000003000030c0003c0c00004c054040c00c0c014000010000004740000030000000000000301d070000000007cc00c0000007401001040310d0c0447cd400111303011133cc00c010104000000303030040311c00003c4031ccc000fc0300010c00c000047140040031300300c00040c0400300c003010004070044d0031000005400c0430001c1c0000303430c00c00c4300cdd1010040003043000404010000000071004003c3d000c7000000100100000c03c00000c001004d013c000040000000500010c00000000000000000c00001c40000140300c04000000000000004000000f00000000c440ccfc1004cc10041c3c0c0c0014000300001000400c04c01c0c34d0050001c05000000c000045000000003d0000070c300c0000003c00cc100c00141c0003000007150c0043000400040f3c0000043010001c0c0007103300100400000c000400100000100cdc00d004f040030031441000c0344004010004c3401c0010040004000430c000c000c00c30d4304c70000007c04410000f40400dc000000003c4700000000c0000000c00013c3440001c041000c001004c0000043c000d30040c000344dc00140000000005000c000000304000000cc40000000000000030000003000000401000013c01000001c304004000001047000c3000000c74500c00403c000c000c1300d71300000007c41001500c01000000d00c04007d07100c00001004000044305c003000cc03540004000c00030c0011703043000003100010100013f0044000000c0c00000000343000030000001c003030001711000400000c000c30030cc00004000c10f1000000700cc040044130000c030003c1004000040000030000030000cc00040433300c0;
rom_uints[26] = 8192'h10c000051400400730000003405ccc10c0500c00400104003000f0440000070003300f11711000000430001030000c0f1030040430d050130043100c1000100000300010304000100000000000000000410000031510c03cc433301000007c1033f00310000330c054111000c0f5033c003c0c0c011004704c1003d0f004130000131000000000f000100003003014110d00400000041031000000000c0100001c1400c0000330c000c0000140040c34cc3411c000c0c0000c3004034100300100500013000c34301cc03010013313005dd1f00014d10010001000001c00003007000000713000000000005131140000100303003100000100000030c000300050711303743c30071444cd0000100c00f4103173040110003c0003000c040000073c00000c141030c00400c0104140d00000003cc0041000011003300000300031c000300411131014300405000c3f100c0010d004400030000c440010000330000cf3030513c010c041134005100c31dc34d131c3c10000100c00c0c0013010001050304d0013000000000000030c00300003c00001c0000004d0d0400000010c10401000300c000f000101c030030110000041cc304103000003105114004400f005c4105003c00c4010d03000000f30000000c01c30c0103040005c011f01c444c0c0130040c001330000c1c4001301300003050f001040303000d10000304000d410311c10c01000c01031c0d400504d01fc30000cf10c000c0001001c0000030030300000110300000c003144000530500c0f10000c00c011c1400311031100011003104000100300c03450000010500331400100100c7c000c40000300100c041130000c00304107340000003c000df401c1101000000000000001030001000354001031000000f01030441c004c3010044c04104003c0000400000040fc000010f000000c003003330030c0301053c3010013d400301000c013104cf01000303100010300043030000c0000c0330f00030000c031d1f000f000001403000040001c001304001030100033003001111710400f00000000c00001043cc0c00030000c000000d401033001010000000414001001d000300000004c0004300c000000001c10100100c0c0000c1003140000501710000010013c1f0010d030311cf000000130000f1c00100c011000100000175001370300f000000100c0504004143001000030710001104013c00001101400131c3fc300f1000400cc00101c574300100033010300c003010000301140000410040c000301d0330104001001010100c44400000030003d00500000000f0007100c33011100000c004c100030000d31033003105010000000100010000300000c003c0c10103333c330403101000000c0500c0101c50d7c310033000010c0001c11010000000050c004300;
rom_uints[27] = 8192'h10330000100005100001000000000103cf000000010c0000f000000000031000010d00000004000000300010030030030000000000000c43010004000000100000000040000043000000010000000011000000400000c00000000004c30001000000030000000c00010400000000300001000000000330000100017000030040100000000000c00300000000000000000100003100000000c30000000300000000000010000003cd0000000303300000010300000303004000c0004400000010000c0004000000000001c000000000000003000000000001000000010000010000400001000ff100000000000501000000000304c000000000000300000000c0000101000000c000000700010000c000000303034001430303030003000001000003000c01000000070000000001040004000c00000103500000000300000000000000030101000000010003c10000c00007003000000000400000000001010000000041004413c00100c100000c000003014044000300000000000300c3013300000303000300000100000000004000030001000000030001000003110001000000400000030001030000000000004000010000010001000000400000000000000101c10000010100000000000001000301010000040300000400000000000000040c010000000100000040010300000000030300000103000001300000000f000c050000c30101310c3000000000c10300010104000000000000000000000000030001030000000003c0430000010000005001031000c00001000000c004000000000300000000000040004001030000000005000001c0004000004c00410000000c0000003001000001000000400100000000000003000100000303040100000300010003030003c003c0c00104000cc10001410000030000401000cf0000010105000303d00cc003000c000100000000000000000000000000000cc100000001000000300000c000000000cc010010030003003d00004100000000000004c0040000400400070001300003030400000000000000000001c000000000030000010000000300013100010c00000000000000000000030001000dc30001000000000000000100000000000001470004c000013000031000000000000303030000000000000100000101010000000003000331000000000100000305000c03030000000000000340000001000000040003010403100000000003400000000c00000100000000000003000003000030030000011000000010000100000000030000000003000000700c010000000003100000010c00000000010000000c03000c0011f00000c4000010000000000000000003000103000000c003004000000000010100030003010001000300000000010000c0000004000000030;
rom_uints[28] = 8192'h14000000100010001010300000003300700000001000000000000040c0003000003001000cc00000000000000005301400000d300400f0001010000c40001000000100c010c000400000000c00004070000303c000000003003404001c003c403000001c30000c0c0000303000110410003c0c000000043000100000c100111c300030100c101000001000304003304001000c0000000030000000041c0300000c001000300f0c001000c0005c000340000000100010100010000400000030301030011000000031040010400013c030031c000c004030005000000000110001000000000c1001000410013000f430000010003c00100041110400011000010031000c0400300300001451c00d1003000130000c004f00000030101003c1300c0000000010013c0003003430000000041030133000400000000000c70040303000111010d1000000c40040043304301c001c00004df00c3d300110000100300000cc003001040010c0000100000004000000301314001010000f30000000010c0000010400000003c0000000003031305010100000000000400cdc010004103010300000001037000000c000004400000000070040303000c0000c000004c00004003000000c04000d4000003000300010000000104044040000003c000f040000000010004010c04300300000003000c000100c00301133400c00000c030300000c00400030000100103000004c003010c00000000070003035340f103c30140434c00c005000001000100300000000040c10000000000c0000300c000c0d000c30000030c000301000003300300014041c000000003000013c000c30003040101010103000000050000fc1041c300c1000400001000004001300041000103000000d1000003000001010100001c00d3c4000040400000003c4000044c000000000001001003000700035304004003c30330000d4c00c04001134000010003c00000000100104044030c000000000101c0c3c0400001004000000100100001c0000c30000010410000010d00c000300101034000000c000000000003034000010003014000007c410001000000000000040c00003000000cccc1034300004030c0000003f0400000000c01c000000000000003001100000000030001014407404300000000400300534101004700000030410300000033100000000307000101000000000300434000003003000140000040000300000333130504000000014310100000000f00c101000400001313c5c0000100000000000003000f00004040000010030003450300001031000341000000100d000440001000000000000001000510030010c001000010004003000000000101000110c14000c1c31100c000c1c00004000000000040010000000113000001004000000101001301000100;
rom_uints[29] = 8192'h333000000330000300000000430000000000000311300300004000000300000100000100003300000041000000000001001000001000001040000000010000000301000401000000010003000000010030030101131000000004000000c3530100000000010100000000330000000000010000000130011000030300000100c03301033101000000000000000000000030510300000030000001000300000100414000030103010100000100c00000000013030300000300100100000003000033000003000000030340000300000000010000000131000003010000c0400100000000000003010003030000000300000000400001033000000000003000000100000011000001317000000033000003003403000040000110000000300000000001000001133000034100000000000c000303400100030300030300000100010000300000300003300000300003004301030001001001040001000003030003000001010000300031010000000000030000030300030003000100000000000000000010f0400003000300000000000300000000000000010003030003000000130100010003000000000303000030c000031001000100000000000000000103010300000003000000000300100000000000011000000001003000000000410340c003013000300001003013011c00000303100301c0010101000000310000013101001000c1304003000040c001000001014330d0000100000003500103c04000010000010003c000030113000000003000330000030001000303000000c000000150c0030000000300030301010000000300c0007000010000000000000300000003001001003100000343000001004003004100000000030001000000030000000033030001010000001000000000c003110000000300000000010704c0000000000000000001000041000105034000c00010001000000030030000000000000300000100c0000300000040130000030004400000000031000070010003040000000000000300000301f3030000000003001303000000000001000300030003000033010043000303000300000000010143010000030000013000004300100000000031000303c30003000010000000000300c03003000300000043300100030000010003130101013100010001000040010100001001000100000000030100034030100100031000004300003101300300304003001001c100000130000004010013000003000010030000c30040000000030100400000f0404000100000030003c00001450300000000000000000003030030000000031000000000401000000001034100300301300001400000013000030300000c00000311010303c10000010000011000000300000000003000010000030010010000010310000300;
rom_uints[30] = 8192'hd0c003000400000043c04003d0000c000d00000c0340c003014300010f0fc0010003f000001004c0344504c3c0000300500f00010340cc43c1000000c004050030000c0301c000000d0000040000340cc00700003000c00011430307c0001000c0403004c5000f00d030400000003003cc10c03000f0100000c30005330fc10004110f00000000000000004000000dc000f100040001300301c0030033000103c0340400005003410001000000cc1000410040000003014f00c40010c30c00003100030030000001051d0c010440c70410cf4030c1040000f0c04004000300000313000000c10400c1c33001010c0700c0ccccc3c0cd100400047000f00c00c3c100400347c000015000c010401f000d4744d00c00f570c473dc03340001470c0043c0000031c0000001c043c0d00c1004c04040ccc177000004034333041c3c0f040001c04401010d7f0007010003c001dcc03003300333d040c10005c004030001400cc30040c100cc000010c1c043c10001004044c100cc10044dcdc003c00440f7c0030000c04130c1034400041f04300003c001c0c0c04c001000c00f4001070000030703c00030030001357d000100003000031dc010400c00400003000034c00000040044000011040000001174dc040004000103000f0003010005470000004704c3c173040003c040cc04005000000c1007c0c00001000000c410430303c04100013031c03040c10011c4000100dc04cc000000c001003100c3131d0044100400f043000000000f330101043030d000c0c3cc300010000040004c440400c0004c00c000000d0344f0000000cdc0000035c000000000c00040000ccd04400004fcc000000030c04340000c00cd00303d30c0f4030030071c70cc0007033003000010004004400000130500c30311c0c074c0c03340300f00c140c00047c4000000330300c0c3c044001013410040c0c000330003f1010304c000004310c3003003004300004300050040050000d043c0433000400000c0c00043cdc10f0003c1c00007c401c000c0040000c000c0107003c3004000000400000074000100c0c0371070750000304000f000001111004030730541044c030041c1701301c0000000010000003d10c1c040070003000000c0070000000001c0d0000300000d0700c31cf0000400450000cdd144c4070000100400011043c00000000c0500004000030000010cc100000004001004ccccc005030000470000007000430040c013c134004700c0030c0144c00001dcd10c040500300403c000c070f000037004030330400004010007f00d03cd0c00c340c3000000cc000000000071f100040f01370000001100004100c00004010440030c00c0300400c0034000c000d101040140d0050300cc00c04000c1cc443000030074c000050043c00000000004;
rom_uints[31] = 8192'h100d0000404140403c0400000c400403c40440f1000041000403000043c0000300c000004340000000740040000000cf4f0104c00000c434004000001003000000000cc00010000000000000c00000c40000000cf000d000000000cc000f010000ccc04040c00c04100044c000000fc0000000440011f000000c0f4007c040403c4cc404000c400000c0000000000000400000000000004000400c00404004c0c103000000000040000000000000001000000140000c330000000000c300030004c00040c0c040c0000000000003f400cc004000000070c40000000c1004004030400000004003000000c00c4000c040000c00c04c00000000000000000c00c10000004000c300000040c000000703110300044000000003000000000000c4c000d1c00030c00000c01000c00100044043000000100001004000d0001014c0c300004c4040dc100000c000c040000400003000010000c00d00007004000440000004c0c000c0010c0304700105004c00c0c004000f0040c00000c001c10c000d010cc00000010000000004c0000300cc0000000300005000000400c0000000000014c041404300c4000030010040c000000001c074000c4c40010cc04004f3000000c000000003f40c3041400000044000c0c0000c034400c0c0430000c30040c4010144d0004c00004cc00004f0000000030f01c00000c1c1404010000000010040c001c0c140400040030400c100004cc04c40400001000f40740100000040000000000c10000f000004c055404cf001154003000400000c0000000000000000c3140000300c0000c00c0000c00040410f0c00c00034000c144300c00000114000000130cc0c000c00c000f140c0003cc041c000c340000400c040054040c4004000003000c00c100c440040030000c000c003c30010f30030c0003140cd03400040000041004cd0c0d0104c00c0070430c000000100000500410000000000000000000100c10000c000130000c04300400005000c00001040000c000300400000c007c0000140404c04014000000003c000cc0040030001000040c0c000000000c34040010cc0000040c4000f0040430000c0004000004000010404c1f0c007d400000c44004100000c004000c00003000001000d00000c0000c00040000330c00000c100000000d0300000d0c5010001050000dc0c000400c0000000000040000040c1c00000c1000010c0000310001500005400030300040040c0c04000c040004c0000700040c0c0004000c0c03040000000ccc0000010c000c33c400340404000c400c0c0030000444c0fc04040c000c0d0000c0c0000f00000c0000040000530c00c0070000401c0000c0000c00001400043001000c000700305000000c04000c000c07c0100d473401033000000c00000000c10c040000cc3000100;
rom_uints[32] = 8192'h40c00000c3474100c34000000003f04001000111010044000140000000c1004000c000430140000300c00000000000000300000c03004000000300005500010040c00300000c0000000000c000000301c0000000c30301030040000300c0000100c00340000000004100000000c000c0c000c000c00dc00000030100000000010000000000f000c00000000001000300301000000000010300000000cc01c4000000c5003000001000003f00c0c3000304cc400300c000030000000000004000c0414000c340000440400050000340000c01030000010000000d00004dc14000000000040007c30000000070014c00000033c00c00c300000000c0cc00030004030341003004c30004c00100c040000100400003400001400000c30c40f301c00030c0000300410330000000c0030001c0c0000001c04000000000000101000cccc0c303c04101000300c100000003000500000c0040010d000000000000410300400000cc00f01070c003400000c041000040030300c400cc010000000000400c430300001400cc000000000000430c00000000c0004c000003cc000000030000503c00000000c30000000000c1c40007c04104d54c01004000030100010300c0c0010003000000000c0000f001000040000000000004c300c3400000c00003004000c00000c1410003400001c14044000004400044c300000001c003c3010403000103010403c001c300000001030001030000cc0004c040004343c0414000c0c00000c44c0300c40000c0cc4003030011000003c0c3ccf03303004000004503004500010071010014000c014100000040c30000000300000100000000d04000000000c300000000030003000300c00000c00000030c10c00000c0300000004000c1403303000000000fc00000010c4130000c4333000300c340000300c03740c000c30400cc010d0f01000f00c30000034000c400000300004000030003c34003c0c000000003c100000000000000000143000000c0c0000000c4700003c30c00030000000000000cc30001010000004041000043000000c4c00100c300c00000c300c0c300c0c000c10000c1c000c3c0404100c001000004440103c00000c44400d00100d00003c00000c00070004301004003000100000000400040c0c0c0010100000003700001c1c000c000000100c0054030000000c4cf00030000000001010100000000300300004000004000000003010000004340c00c00c003003000040000000000000000c40300c0c0c040c311013005000040000000c100000000014f01030000000000c00003c0000003c001440003c0c10000000000cc00c04111c0000304410000010400c14000010000c0000c005d00000003c30043c3000000000000000000c4010040000c0004000000000003050300000003004100;
rom_uints[33] = 8192'h4000000000000000040400000c00c00000000001c00c30000c0000000000050000c00000c0400000000000c400400cc070000704000044c00001300c00000000000c0c000000004000000000000400000000000000000c0f004001c000c004400000000014c0040000000000000000000000c0c0c00000c00cc070c000c1700000c4f00000c000c00000000040001c000000000000000f00000100000000c004c00004004cf00000000c0000c004000000000000000000c000000001c000c0ccc4440004044000000000040000700c01000300000440c000000000004000100434000000000004000d0000010c00c00c0000000010c00000000c00004000001400400004004000444c047000ccc00000c1003000c0330040000004d04ff00000c0400000c0c0000000000400c400000000cc4000c0040000000000400400000000000400004d00c00040c0400c0400c00000004000004c40c44400000000000004030000c0000c0000340d00000c0ccc00cc000c00c33c40010700300000004000000000ccc000000c000000c0040000000001c0000044040000c0300000000c00c0000414000f00000000004000c003300c00040041004c04c0c040c04c0c0000001c404000c40100c00000c0000c4000000c0000c000cc0400000000dc4034404c000000000c40c0001000c000000010c0c0000000c0000c00040003300c000004c0000000c000000000c40740007040400000d00000c010c000000c00000c000c00c01400000000400000000000004004000005000010c000c00000043400c00000011000000c0040c000011003000c0c0000c000d000c010cc0000003c000c00440004dc000404000c044000000003440040040030000404000c300c40000000010000000000000000004000000400c0c003000400c0074000004001010000c000000000000015004c0007c000000c3000d000c0000000000000000000cc000400c0000c1000c000000000c000c00000034f0000c00000000c0040c0300000000030000000000c00007000000000000400c000000000000000034c00000000c00000dc000000004000cc0003000007c34040100000040c404c70000400003300c00000000c00000000000400c00000400c00c000000cc00000c00070040000000040cc0cc00001c4c00001030000040400000c400c003004c0000010c10130414001d00004004cc0000070000c400430407400c00000040004000000c000000500000000c00c40000c000004c000000c000000000000500300003cc000000000000004104c3000000000c00000000000c00c40000c00c00400000000000000c000c000c00540c000404010000004c000000000000000c4014004c040040010000c001040000c0300000c0c0000c0c000000000040000cc40c0d00000400;
rom_uints[34] = 8192'h34000003c000000741000434030000000130000303c000000c03400030040110001004300d30000c0c0000300d003000c1000030040044003c300700040300000c0704010000300000000c1f00330010003000044300440001100301003c0010003135c007000000c040c000000400041c1010c004101c01037c100000000003040c1d0003000000000000d030301030003000000c00003cc40d00030403041000f04000000c000403100400304103cc0c0400000003100000c10c1fc000c03030c00430000030040c0c0030003704000003000000c7040030d404000040030000000c00033030003c40001400c30040000030000100040000030003000000100100040f10100000040010cf00000303c001030000043100010c374003c0000c0c00300c0000000033c00c00c0cd00d03c41003410040c0c000c00071700031c0404f400010c0000000001000030004010000014301100301c3030103c3034030100000f00000444000c010501c0000033010cc040400500350004c1340c00700000c0301f301c0c04300c03000f10d3000070300004000f0c3301400000010f07c01034000410300700300100030c0c300003cccc1c040133044100000c51c000400100000300100f003000cc00010c7cc40000031f140010001104f0040c310d000040c0130c03000104300300000300000131300000400c03d05000040000c00450013004c0300004000c0000004c0d0100034000c3000c0000341035c00c1c0007030000044000014c00300c14000c10000f00305313c404300d00000cc041c0000c004000000c00740000130c3001303700003300000c0000301c040070c10300070c000c40000400011400130040000050000000cc00700c0030353c30000c0c0000000000040d0004000c003c00d340300000c3000004010c00000000035400030300000fc030d04433010c1c000030001000000c000d3c0010004000c033000130000c070401000000300c00010030c003033c11000000000370303100000c0c0000000c11340100000000000c00c7140030001000000000030003000c00c0000c000c13310700000300003303010100000000c00005000cf0cc00100c40000c00ff04000c000c0001c001000100c00014444000000003410000100000000100000031c0010f300c0f00c400000000c01100000c00c03000000c30030100044c0000000d07100001300000000cc40c070440040440100000033f0c050000d070c0003001000403000c000c1400000004000400041100300010030000f300001cf004c3340000c3403403000000000c010003000300030000000000003400073007c405044001000000700000d40431010444100300103003010f4c000c0c30330c0004000400c03f03100c03010c004000040003000030334c1c400;
rom_uints[35] = 8192'h100030004010040000c0034340034000300000c0c1405000030000003c5c00000000c4300000003001130000340000c040c00141c07000c3cc000004304304004100700030000400000c410070000c344130010001c0000000c330f00144000001c444400100c000000331c00c003000c00000000000d01400001000330010c00d0000000c400000000000000001111030c000000000c00000000000c00340c031d1004003000304003700400100000000d070000000304050c003c000000000c0c03c00000311010000000000107000130040000010340403004370000103030300000003004000000001d00c00d000d01c1c001400300040000000000000001110431000000003d000003031400000301000004000c004d70010c0504000000cc00000000000000000410010003c43010cc000301c0000000d00000300c30000c00000c00c00001140001c000300c00030000003030030004000c0000c0010000000034100004030c00000000000c0100000500000000010043001000030c010000007004074000010004c300030300000c000c0000003d07030c11110000010f0f00030000740c04000000000405050000d00103000030040305000c03cd001000010300f04300040000c00000000c30000000040c0000c3000401331001cc00040001400503050000000001000344030000c1007303000003000500000500000040000c30501d0330c10000c40040000000031000003300cd3c0043040c030000c00f0c04030000000c4c000400010100000000000c400300100c00100004000c0000000d003004400000000703100000001c030000004c0c00300c030c03c000004dc00001040003300d0000c4003000000001000000140041000c0040041003000100000300007000400000001c0070010000010000040d001d00c100140c0703000004040c010f000c043000070c400c000c0010c100300000000000c0000033000003404313000000030000000400010000004004040131000001103c000000000000000001001c1005030c3100000f030330040400033330010c00000004011000000c10000300000d0430000c00011003000003000000410c0c03701000031d40040150000000000100000041053500530c41f30001100dcfc1000d013c0000000d004003040033010c00001700001011000130440c0000100301000004100dc0000c00000c000c040300040011c00003cc0003fc043cc4000143d00c00001000cc0000010010000404000400104100000c030000cc4c03010000000343004c4000010010041c3500000300003c0c00000500000000000c01410304007010000403310030c000030005010000444000400c000000000100300000010000400000000000d000007c0001000d000000400000000000004000000100;
rom_uints[36] = 8192'hc3c00000c0cc0000400000000000001f0010000007f070000c30c1000050314000f0401000400000001040000010001c73d0405344c0c0c014400001cc0000000000cc3040000000000007cc0300040000000cd0c0140c004044470000700041003d040050c1034000c031c0000000400000d04003c100000010c040c03050004301c4401000030011c0004000000001f00100000000c0c000404000c0c0c0000c050c00000000c3000000c034004003040041c0000cc0f00010007373c0440000400000c4004300c000030040001c000000cc13001103400c070cc440000033040003405c000cc000430070004004004000003450c00010000130c0000000310000c00004000f4c4040430000d00030040140300001c4404013031303c000000047010013c001040000c001400c443100c00000c00c000000003300330000000c0001cc0c0000c301c0f001c00430cc3dc401007100503540530100004030d710010001471000c03310c0000001003001c0010000300dc0000170f00003040d0040005413c100c04400000000004134d000c050010c00010300c00f300cdc00074cd0010c0440c00040c0c14400f00330c0003d01f0000141c000400004303c034040010000001400cc000000000000030000044000c04010000000000101c0000000430004107441c003c00c0000000004001070cd301003414000c04100304040c0144301c0004033c00c005c10000110c040c0c004c00000400000004000040040000c4300d000440000c000d0443107c140000000c3004cd030440000110000010003034000c000c001000000c0001100300000f103f00100004300c007000cc000104c001000c000c041c000401c00c40710000c0001301000c04041c0400040000100030cc4c0000ccc0c041c300ccfcc4100511400dc0040c5400300000c0000f3c0400005303137004c0c00c00000100c00400c030c44c0c0430000004000330000c0040000000c000440cc000c44410033c0004100100c40003c40030000004004050000df407130700000000140d000000000c400000074c044c00300000003cc00c40040010100000140000040400c0700303c004001c00c00c0c0fc0300400004c100050cc0c000430000401040000001000c3001c0100dc000040013000d00c0005013c00000430d41100d004d444030004033100000c1cccf440000c13f000000003d00c04000cc0000c1d0000003034c7041c0400040030030001d00300000000040c0c040c00001c010cc014d0003001100cc1030134000400000400000401000000000d0000c0000050cc000000000c0c100000040d130000c1404cc40fc10cc0031310c1040004040c00330c00400dc0104030341c040f10050033c000010c0004000013000003400400304c000710300c0c05400c000;
rom_uints[37] = 8192'h3c14001004d430305003044010001000001000001400d30c0030100004103030000070700150000c0030100010100c00c000001c04f000403000300440000c000000103010f040000000003c000010040000c4d00000000013c1500100100410004c003010005030301c01101d4c1c0010000000003001300040003c0000f0001c003000040000c300000000000040030000c00000000c003300c00000410030003c00000000040000000404001000cf0140050000001030000000004000c0004cf0300000004000c0750030c0000410004c00c000cc00100f0c004000700100005000001010400500440070000000004c0000105010000c10000013000000003300c1401c303030313c000c0010100000f10030100c00cc301004cc4000c4500c301000d3c00c0000301100300004010010000700400010000030500300000010000003003c03103004000c3000000cc050040000101030f1103c000010000400000000000100000430d0001004c03000000c000004003100100000000010010770000000101000000430000c00014010000010000031004000000130000000303040000c0000000000000000c00010000000f0c0f0000010001011301c000c4c00403000c04000100000000410400000100000005034d0005000003c0703f400001000000410300010040000700000100000010000c0000000010000001010f0000c300031004000000400040c101031dc00001000301004000000141c000c14071400300c100000000100300030000000000000105030500000500c0005f000000000000ccc000c0000010030100000c04400340c1c00000c0010100c141cc00c00004c4010c0f00010100d0000000000101c0300f03030300c000c00103000000000000000c101000c00f0f0000001100050040f005000d010001130cc1004100c00000000d0300430c40000043000300033403100001000c013000300000004c01000000010000c0000000400c00004000d0000703404040053c4003000430000000000300030001031000000001031303c0030003000000c1000000050d0000710f30010401c100000000000010030c00001400030003401c0014c00410c000050303000000044000000001000101000000c100c0000003c0000300c0c30fc40301014033ccd0c00101000000000000000c03d3030c01400000000d40000d0000c0010001c30001c30c00000001400f0000c50c04000fc004c0000c0000c3004c000000c00d0000030005000401000f000103000000c103c3c14000010440040100c003003c40000005000000d00100c004000004000000c0000000c50000030c04004001030000d00000000000010107000001040000c0000000000c000000000c4003003004031100000100000001000003000f01000130cc0100000;
rom_uints[38] = 8192'hc000003041000f1100000001000401c000c000040c00003040003070040c0c30c00000304400000000004010000104400301050413033c00010000c1470f0001c0c044300000300000004300000134000c00c175c3f500040014400430d004001f104c300f000d0000040c0000000330000c01031c300cc0c470f0101100330105041000100000004000000000400010001000000000c000dc0001130301c03000000c000004000000000010300015000334000044100300400000050000f00f0c00000d041444000000010400010d3504c0c000f140300010431410140100c104000004c000030000000103c00100cc01700100c40000040000030400000100c0000c0d013000c033c400034403031113000c100010040c00c30070f0040000c1100001700001140c0000050030c0300003040000400010000003f0000000fc0c0c0f03401304c3c3000040310c010c0c04000011c41c0c3011000404400300cc0003054403c013000c4c13c1101304030005003100400000010004000440014541433003040001000000c0000c5300000304cc00c300030000440c000000c0000400000f0c00100100c3100f0c001000310c07d03100000130c00011040f0cf14003034040d0003003030000000c0cc50000010003c00000004405040045c011300c0430001c0400003c0000000030000117010d0033c1310c000000000001c03501100d10c040d00d1100c00101d0100700030c1430471070001000051fc3040011000000c4000000001000000100300d003004004004500003100003000010000070700000c4050000000004000077f0000000100100cd0c0300000343300c0000000510000034001000030000f300010f0004000033c51003d3030001040f017400003c00101000030030c0000104f4033000c14100000401c0303414430500f50000000010011c0c003104000013310c000330050000040131000d300001cc110000400030000030000010301341101003f000cc440034040030430400005100310004300000c44f0c00003f30c000c4404300000045c10011110d303000100000d7001001000010000c000001004300510001000c0000100d300000c03000003000040301100100000001100005040300010f000070031403c00400000c030c30340010303000f1310000c0310f00400d000001c0000000100300040c4440033c400003d04f0c101c000c1035000000010010000c03003c10040703103c003331000000000000001040000033c003300cc0d0044c0000c01c00000017000f040101cc1400003100544000000001000054000403001000001c0103030043c01350d400044c010c40000074303d0c1100000c00cc00000c000c004001034001000010000503c00003103c0300400000341000300c0100c17100500300;
rom_uints[39] = 8192'h3000000030010c000100000400043c103010000400100c00000404000400000000000000000000004c00040c003c0c0c0004010000340000c03c3c100000000000070d0301000305000c400100010c00d010000f000c00000000c003000c0344033000040005001c300c0000000154400c300007c3000000c0300107004000050100000000000000040c00000440040003000000004001cc04000c01040f03000c000000004c000c04000004000001000c1c040000010500000c300c0d0030001000000400050030000001100000050004000c00000c01100410000054000300c70400000c300c300000cd000c0c0000000301000400100000000740000000050c0400011c040410031000300400303c110030001c0c0c00040040111c0c000011030004330000000001000c0c0c00000000000000000000cc00300c3c0040000c00040c000004dc05000001000c00000034000005000040001c00000c0c0004000000340030c0300c04040000000c0004c00c000c10300c0700000c0000000004010041000004100c0000000011303000004400000000070cf00c0c000000000d400400000000000c000c000700050c00101c000c01c0c0000000350000400000000c1103040004040c00000000003c0000000c00000400000c000c000fc01301103c0013443300041100f0000c0c0400000c0c000000000c040003130000000000010011000000000000040434140033000c0400100000000c0014000cd00c5c3c001d073001000000003400001c000004000030040043003c0c000030000c00100c300c0c000000010f014000000001c00000030000000400000400000000000700043c00010c040400c0000d043300000410000c000c000700000033000000100001c00c0c1004c0000c0100041c00300c0c00000300040000141c000c00003100003c04135330000c0710000c0c0c0034330000010cc00130000004000c01100003000004000c0000000cc00f3001001c0000000c0f0000001d00000f0400000cf1001c0c00000c300005000000104c013000000001100c00c403000003000f010c0004040004040001003000000c00100c001003000c00000d030004000000040c030003000f000400000c00000004100000030005030000000c00400c00000000000ccc041000000540100f000c03130010000c0c0000000c003330300304000c0f0004000000000000c4100000000000000c0c011c0000c00c3c0c000000000000000000000300000004000700000000000000053410000003040c0c0040040c470c10000c0100070c0000001000000000000c000c15000441000700144403301c10340000040000300000000000000004030000000c0000c7c00000000c0001000cc4040c000c000004000c000100300c4c0c0000003000040c00;
rom_uints[40] = 8192'h1001040000400000000000100403440074040004000c000c0010c1c400000000300000c00c400010000000c0100cc0c04c00000010400030000c00000000040000003340000000003000003500004000000044c030104100f0100c0000301c0000300c0c00000000400000000000c00004000000000000101030410030100000cc03000c340000c0000000c000000000004000000000040c000400000c003430000000000df00400000400003000303013004000000000c030000000000c000c0003004005000c0000130c43000040000000000c0400f00004f030cc40001000c00000000000f0000000c05d000c030040003700000000300040000000000000400010c01d50f40400c00000c1000040000700040c400040000000004001500000070000040040000000700000000c000000000044044000400010c0000400040d00c0000000000000d000000400cc0003003000430400000300c1004040000000c000000000030c400cc00c0000000fc0000c000c4f00303040f0000000003003300000c100000040000000c40043c00000000c0000000004f0000000000000000c000000000030c0330c40d00400000c040000340010003000004000000c040000000000000030c004000000000300c0003003000140c700000040000c0000004c0000410005433000400000000040401300403000c00040000000300004000000400100400000000410010004c10040c10000c00010000000000004000400000000000400c00c000000000000100000010100000c0004c0c00c0c10000c000000000c0400400c00000c000044000c000c103c000000000014004014000c0c00c0000000340c01000c303c000040cc04000c0000340100000c00000dc00c0c000000000030040010c0c000000050c00014000c0c0c00000030000050101000500400007000000310000013c0440c000c1c00c1f0400300400010000000000040000000000000c0c40c00c10000003c00405005000000100c0003c044000c00c40000000000030000f000030c00000000000ccc0c0100000c30000000000000000c0c0cc40000003000000c00003000c000000000000000000000001cc44000404000000004400000000030000c0001000001500070000cc30000040004310010014004000c0c000000700033000400400c0001000000d10c40000000040000104000c040f500000000000c00003000700000000004000000c000040000000030000000000000000000001000400c040011000000000000040000101cc00030400000004c00113000003000c40000000000c0400c000400040000004430000000404100300c4000000ccc0030f0000404000000000000000003000cc4000001300c0000000000c0000040101304f000010c000000300000000c0000c3000000;
rom_uints[41] = 8192'h110c100c00c04000d07003007000100410d407000003c0000143003010003c00000c30c00c70000000000307000000c300dc003c01400304c000000010000301010001400c4c013400001130030d004000000304000100c0d434c0300c0054000034c400000300000000504000cc00004c40030c404000c000000034040000001d00314000000c4000001c0c0305310004100000000cf000c030c0003000033000010000c3c30301400000030d3c0c3040031c000014cc0313000c01104004130070400000000000300300371030503003000400001cc010003030700c0000030f00000c0410cc00000000100130d401100c003c07000004c40000000c00040d70300c043104000040c04073c0c0000fd03310f41400000000000000400414c00043c00001c044d004000100000000001100cc0c45001011000d03c1044f704cc10cf0ccc03010000c30010c000d001110400044143417c00c04cc004110030000c000000010100404400103c0d03000c0030000105000c00140000044000004c01003cc0000000140c0000c0001433010000000000000700000cc0dc100000100110040fc00000001c300100030c0c0000000c430404000000d0001331301f0c000000d000c04000000c00c00004000000400004f004fc0000c001000040010440000041c40074010330100000004074000004004000c00001000400100001c00001410c044004000000000747fc0300c00300000044000440033030000000000c701000140000004400004004c000000000000001c710011c000340003071d07004003d040400414000000010000000117000000100000303c0003300d3000003000000c403000000004d100c04001c003043000c1300000070004d000100c0004100000030000000400300d3300004c003c000400131003d0c0404d00000010401c401000dc000004350cf34000c7000340c001000c401400400004d00cdd000c104000001c0300000cc00010000000701410c000300040d0ccc0001000133000400050103d000cf0000000400070040100c03c3010040400700434300000c000c000c41037c0000404000c300c0c000c0400300404c0013104000003440441000000d4001001100000000c03d00004d31000c0100000c004f00000000004100010001c0004c0104411300004000000d100001c40045143c0400ccc300000040000c0000000000d003400000004031470f00050c0400d00c00000cc00d00000000c0dc0000000d300040cc014043f33000000100030000c017000f0300400c00000040c00031100000100cc00000400400000101000cd00000000140400000434141000103010030070000cc0113003041c000444004d3040003034400c400300100c04000003c05c4c343033c000c0000004d03d0c03000410001001000;
rom_uints[42] = 8192'h7304170c00000030050030304004400000301000c010100c3000000cf0051400000000cc1004115c000031010000000cf4000c10303c0030034000300400300c0000000000f0044000003003000c0c010c441000040300103f0c0000000cc11000000000001000305013c4003000001000405500f03c05101c0000f010007c305000d00c30000c50141400004000c00013330c10dc3c0f340c04003c40f00011c0000030000010443c0000041010000034004000000030c03150c05f0000003034100017400300000c3c0034001d30110000014370007c44000310000000000000103000300c03df300c0303c00c34100000403c10000000000040000cc01404540040003010c030003000100031100c00cc00100703304010040000c00000c10010103000ccf0005040001430100003400000000c043f30700030000004000ccf0000103003c040003030c100c30015c100c40c01c4430c30000400cc000030f0003000003000000030000070100c03c1530c700400c030000100000c04000070040c0c000000000004f04c00f030000c00044000c330100400000c3030c03c0400000000001000500030000f001c03300010f0003cc0c300000410000c00300400431013c00c100400330000300000504000000f0100100040030000c00000c0410c1014704004000c710000003314000034000000030000310c0000c0400c010010000300470040c0301000c0040005400c0001400410300400004000011040303000400104000000000354400000040f000001000010010c00dc100c0000c00013007030000c0000000c00040000007000043000040030300c043400054344001c5040500c00004010c0004400003030c030001000000000300c0c400000001040001030401000000c1000300c400444300d0700040c0c0000103d000000370c0c00003017001430110c0000001000c000300000301001000040300000000004000000c00003c0300001001010c0040000c010c00c1c1030c5c000300cf00cc4000004140001003cd400003331000004003c0037000c13040c0000000030c0300340004100040d00000c1c0001001000100c030000300c700130cc003c104304ccc040c00c00d03005001c5c0001c0010400101030c00c000050000000c00000c000300000300000000d1c000c0403131034003003300c00000030c00000700000c0000c3d000000000c001000044034000c3004701c30000030010cccc007c00000000000000410404c000c11c01c00003030400c070000300044c10d000c1000000000011c0401100030c01c0000100000000000c030143000031c103011030030301c0030c0000000001004000000503000000031d0300000000000000000c0044010000054000c3004003000001d143000011c3000000;
rom_uints[43] = 8192'hcd3000303c0001000000c0030c000000700300c300f0000311c0003001c0000000f0500330000000c00004000400400444000001f040c4010003c1100003004000c014401000001000c00cc10013c000000c00000300c00300d004003001c00000100100000c030344c0c000000104000cf03cc0d100000100c0030050000030f000000c00c0000000000c00c0010000310100000000110c000401c5000000030033000003c103000000000003c00440c0ff00000000000000000001c00000001cc0001c0010030000000c000000000000f000000034000301030140030000000300030000030000000030004f50431030c01000000003004000c300000040c0d0c40c000000003400c01130300000c0500301033c004001030010003000010003000000700000010c030001000030030403c0c0000000003000c03c400300f3c0000530050300c40000331000000040c14300fd101001000c150040001000004000001c1001c00005004701004014000100000400303000c00005000030040c0c0c000410c0001101000000001000000000c000000000000037040100c000004044001000000c000000000000040030300cc03000c000001003c307500034000f00310000040000404300c100000003c0000104c0c0030000000000004c0101003c000000300c00c40000000f03400f30000000c0030000000010000c0c7f000000014000300c1430c100000c04000013400000000c03c04c43110f00000000c00010c01103000001030001000000050c300000000300004040c04400c330c000410330430000000004cfd000000000301c00013000000100400000000410c0c000434ff040003000c104003004c03300000100000c00000c000010000001c00100000000cc70100040433fcc000010f003000000000000031010d0044030c5000000304000c000c0104111000340040400100000300c010015410030110030c0c0c10000000000000004000000300000100000000000000000c0003c0403000000cc03404000000030403c4001003004001000000000030050000000410000030000001c00d0f00300010000400030013010400000000014030000000000010300c030400010c314000003000000000cfc000340c000000c0050430001000001000330030040004c01c000c0000000004404010400c00000d0003000300000000040c000000014330000110001500c30014101000000031400004000033000000000000000c0030001c000010000c330010c0300000004000000010000001c0000431d03001110003000043000c0001000100400100000000000001c4c000000001130c03000000c440000c00400000c000000c000cd030400c00030000700500000000c00000130c00040000c00c0000c00000cf040030c000000040000;
rom_uints[44] = 8192'hc000000000c1300040c000004340c000c0003003cc014051000140035c00c30304303d304010000103033c0073010410f03d00030c31d1c37c03000001100c40010007c5000c30c000000000c3003cd0030dcd0034c000041031300100001000300070010400f1f4034041c071000170070500501000c4000017d040f0003c005500340040300030130c00343000c00001100d30000030133104301041005c74001c0000c000733f04c130001000001d01c7000300000501000000c4301000101c04003c33c040104c0004500040cf040007300f00c3470000700011c05c004000000000304400000030411000c40100c0340330c001c003010d400f01000004d010fc00d00103001c00331733000000000d740f000c300000c00730c1000000007000000300c1033030d13103c000303000300330d30000300000d00010c0c007301070003dc010c003000dc0040004c40310000f010070343c41001001010c04130c0c1f7070d40470013d0000050c0004c1c040011001400400010004001c0c0d400004d0c000010c000000c1d4d0000c040003007000c003370c0c0110001004400c10030400c03400c0001f0330101000c34c44100001001700031103000c30c40ccd0400000c1451400000c0000c00400cc000f0040073c0015000100c00c014330300034d500004031cd7c000c003100d4f10071000100000d00000340040100001cd41130004cf0300c30dc0041001001400d0070004c3c047050c0103003034040c4000400040003400c10130f05410040000400004001001000f0c014cc00c0041f30144c0040400c0400cd00043400033dc0000c4030007c0cc3540100030141704000f0400011041c04007dc00cc00d00343003d43c03c00000003000004c403f30c051d004073003113c10014d40040040000030100d0317000f10471170003c000005f3431134f050104f10013001c0013000000f000000334000013003000c1040400004000000c3040130051010000c3010c0c43400000003000400f470010c0000c0001014004004000013500000000414c0400c430f00034071004774130ccc700400001c0400c17400000053001010000000c1014c0c133130000f340c0c00000130c100030000000030cc4701000011040341c310c030ccc00c010040f41374070007003000000710040304000c11300030000000c400301c00700100000f41000f503000f010cc00cf00000c14000f000000000740001030417000000100040000000c10c04d300000000005c0d3004c00005000000410007400100001d000c44004000000400c1003130000d001001000030c013c04030307d1031000070000c0f000c004000000d00000700000300303c47401c4f400c3001000000140013c0014504d400300c03c031040000c43000c000010000;
rom_uints[45] = 8192'h400c00000000000004000404f000c0000040040000300000000d00000040000000c00000c000000c00c000003400000c0000000c00004cc000000000000000c040c0000c004000000000c040f0c4000000000c04f000cc0030400404000cc04000c04004000004000000c0000000000400000c10c04c004040c000c40044400000000000044c00000000000040000400044c00000000000004403000c400c00000000cc0000000c00000001000c0000000000c000004c00400c400040c0000c00c45000c00000c0000c000000c00c0004000c0c400c4c0000c000000000c00c0c000000000ccc000000c00040000040440000c0000000000000c00c00000000040004010c400000000040400c00000000c000000000c000000c00040400040c400040000c0c0000000004c000000000c000c4000000040c004cc000000c00004c00000c00c4040004000cc4c440000c004000c0000000c400000c04c00004c000440c04c100000000000c044004c404000000000c0c010001040000c0c00004c000000c0000000000040000000004004c000000000000400d0c0c0004000c0001000100c040004c000004000401f30000000404000040440000000000000000000c0004040000400000c0c000000000004c000c0000001c00000400000c0000000001007000000400c00000c00c040000000c0040040000040000cc0c00c00040000c00400000000000cc0000040000c00400000c00000c000c0400000c00000c0400000001000000004000004000000400010000000c0000000000000000000004c0000c00040000000000c00000c00310c0400040c0c000004040000c00c0040c00000000c0000c0040c0040c000140000c00000000c00000000c0000000000000040000000c000000c40000400400000c00c000c04040000000004c0c000040c000000000000c104c400c40c00000c00004000000000c00004004000004c00000000004004000004c00c0000c40c000c040000000c0c40000000c40c0000c0000c00000000001000000000000c00c00000c000044c004c4040400000c44c0c0c00c40000000c0c04000000000000cc40040400c0000000c44400c04c00000c4c000000400000000c00000cc000000004000000c000cc0000c0300004c00000000c4040c0c0c000404c00c00000000004000004040000004c000004000c00004004000000c0004004000007000000000000000000000c00c00000000c30000000000000000c00040000000040104c04c40c0000000000000000c00000000c000040034c000040c000000000000000000c040c04c0000000cc0c00000000f00000000c000000000000400400000000000000c0000c0004003000000c040c54c0000ccc0c000c004000c000000c0c0c0000c00c00000000000000c0000000000;
rom_uints[46] = 8192'hc00000040011500fcc0c004f000f30000000d0000013000104430004011330501334000f10000000c4000c00c00c0f04400030111010303c30c007033000000000030c00000330001000070fc000c10330310cc0c100034c401c004000113140c3c3300300c3300407014000004040130c004000000010c000000001cc37400c000dd4310000000003000100000033000010000000c70001000401013304c43c3c1430000030c4f004c00000c030504104f4400000c0fc000c340010003400040c100000c00c305000030111001070005000dc0000100000c400c114000000f0414300c0070400010043c104030c00000303000000000000050000070000000140c0400c30c3c00c40100040004401031c10140004143c000030c03d540103f0c0110000c3011000000031000000005053010010c4000000050000f030004003000304c4f00030045001034400c0033003000304000c401000c0031040000cf000010f3133400333c040030030000040010511004c00c04003030500000c3040000c130100c300004400000000000c30c00030000000000c001403400000300cc043104000000033000004400007d0140001300410004000400340000cf1c400000c000000000500001100000000000000000400100440000cf01000043f01c0001014c001000000030cc41d40014c0000030000000300730001000c40000f40d3000c30053030c300c0000c1110030003c03000004c000040353000003c5040c010000401c00c000000c00cf140000000c00000717033000300300000010010011000004003100400c00c0001300100050f0040040000100cc0300fc00440000300c0444010000300c0000c00000043007003c0070700c00c0c0004c070400c400cc4140000d001003030300001c00d10c0330000c00300040d0000c04c30c51004000413d0000d03c000300300013004500034003c000000001000c00000c05010030cc0000031001000000001000001400c010c04f00004100300000404103003d01d400c004403030f41100000300040c303000034010500014000c3000ccc000013c0000d3001000130000000000443404f0c003030000044003304c434f0c00305013035440300453004030440000000030c00000040004c0c04400c0541000c040007cc000100030000c01c000000400013d0004c7cf0f0000003c00000040000d3000030c73030000000c1404130c30000c01070054000cc0040c3c000041d4000000001001004100001000040003c004f00000300c400030300000000003001001c000000c010030340c0000c004c0010003000000d00030003340c000100f000000043003100004f0004000c00000000c0c15cf040d0f0c074040400c40c3043000031c0010000000010000c0c00c00003c4400100030000c0000;
rom_uints[47] = 8192'h10000000000c001000d00000000030d000000000c000000000301000000c000c001000047000000000001000000010000000000c0000300000000000000040000000c000001000513000000040100030000000c0cc0000100000003c000030000050c034441050001000300c30400001c00000c0d0303000001000000030001000000030000000c010000040000000000000000000001000000000004011f00000c01c300003701000000000303000500010300000000000000400101000000c0001401000004030c07000300c000000000050c00000003000c010300504301000000000000000040100000c30c010041c00d00c000000000000103030000000404440004400103070541440000000000000000000f000000010101c000c100000000000003000300000300c1010f0300000040cd000300000000000df001407001010400001000000010000401004000300000030070440c0004400c0d000040034000000000000003000113030040000000000000144c0003500300100c0000c00c00003c0c0000c00000040004004030000000000c430100010000104000044c30000401000000010c000040030000c003030300400000000000110000004401000004000000000033000000000001c0000001000400000000000003004d00001f010001000f0f000305c0000000000000000000000013c3030000000c01000000000003cc4004070400000044010000100003000f000c30000000001c0000003000040d00000300000000000300001000000000000101010c03000000400000030000040cc000030100010310000403100000030000000514000400000010010003000c0001003000c0000044000d00030000000d0003000040000000000000000000000003010140004100010000033d0100000400000c000000d00000000100cc000500300c0004000000300405000c00000001040c000300000c0400304007000000000100000000000000c0000470440300000100000c0030030010010000c00cc00301000000001000000000000f3100004100000301330000010000000301c1c30013010003000301c00000333000040000030000000040000000030040000003000004c3004000000c00000000004000400004000001000400f00c00000400001c3100010000000400000100000000c01003c400040000000001c040000100000000040f0003000001000000000041000000000100010001010000010300010004c000000003010300033000404040000000010c0c1000000500004000004000010c0400000103000004000000010c10000000040300000300000000c00040040400c0000f00c001000000000000000100000000c0100000430303004c0000030000000301c0000001300f03000d0000000c0d010c054c0000100;
rom_uints[48] = 8192'h10104000c4000010c31003330000050010000000003c03c100c00000400004000c040c0030c000003100c00000400044c0000ccc401000703010f00400001000000300000c0000100000c10c0000000000001000000000003450c00000cc30300c0c300000400000000010001140cc0000400cc0034000004cc001d07410000c00c30d00000000700300000000000000030000c0000d000000c14000004000400000000c0430f0c01000303c0cc0101100103010000000043000000000000010030000c030030c00100000c0000300000c00000000303400400000000d00400030000d000c01000010100dc034000000c01003c400000000005040c0000000001cf00000300040004000003004c1000d31100cc00000c000c40010450030003000003000444400c400000c005140000004000cf00014000000001000103004000d00f0000004c000000004000000000040000000040f000000100c000010100000440000c4c0000000000400000010100000d000f000140010000030000000000010c0010000003001c00000040444000000000c000000001000040000000000d0004000000030300300c00010000d0000000000004030c00000000c10c0004000000504c000f3000c00c00000c0000cc0300040c00030c001410000c00c011f0000c1dc00004400000c100300500050700c00d00c401330300000007c104c00300003c000000003000030c00c00300010003c4000004000004004301003000000c04c40030000000000d00050010030d300104004304300301000000000c04000000030404000000010000011101000001010000000000000401040000300100000000000c0100000000000001000cc50c030000000001400c0000cf0000000c0cc0510004c0000000000007000c00000740001000cc0000c00000000101004300030000000000c4cc05100000051040000c044401400c000000400000c00c00c0030f00000300010000000000000000400300000c0003000000c05c0d0c0004000c0001000401004c000100c000000000010140000c040c00c00c0503000041000f00000003c00000400c0c0400000000000004000000004000000c430004cc0c0003100130030101000c01030f0000c0010c0004000004000403000000000500010440000000000000000c40c0c40000000c00c1000c00040000000401000000000000000000000000014040010004000c000030000000000015000000000500440000000000010000c330403c01001700140000000003c050c004040004010004300d07c00000000c000100cc30000c0f010000040500000000000c0003c00c010300c3070004001d00000c003000330300004000070000010300050c03000400000c00003000010c0001010000c00001000004c0004001004300001000;
rom_uints[49] = 8192'hc1400300004f000000040030f000000404000030014510000000300040000004004300c100010000000100c10000011fc3004005050c30f0c1000000030000400305000404040000100004c0010000340c000000334c0000300001000c0c04c400c0000c440f000000003c0003007cc00004034000040001000c000030300000c3000c04000c0000000340000501000c000000000000000c40001c30000100430400000000c0000007010000d0000505000030030000300000000001d40c0000001000000000000d000400000001400110000c0300050300c50300c0070c01000000000000434000000100dd0044cc0f300101c00500000000000cc000000004010d030011010040c01c000c000c00000f44400000430000000001d0c5404d4000050000040c010100000700000040000041c04c0444c000000c1cc000040100000c00400c370000400c03050000000c03400300440c040c4400010c0000130c01043300000000034c000cc030000f0100c040000000000c100400000000c3000c00030c000040000040001000000401cc000000000007040c0003000100c00001103405000dc0430003000000300c0143000404000001c0040003000c010d01c30000000400c10000004000000004001000000030004003000f000c0003041c0000001cc0000000040c00000000c0400c0cdc04440300c40000000000cc001f000000c14c014c04c140040003c5c0004000004403001000c400c100000000010c0100c0100000100000c0000f01400004300c000c0c3c4c00030c000c00010143040500010001000000003303000300400cc00f40440d000304000000000f001100004001010c000000700cc40cc10003000000000c0c00400300000401000f0000000100000040030c00101010c100010310000000c100000100043000040040cc0c440c0000070741403cc0440000000c00100c0000c5000045000014000c000000000400c000030300000003000700410001030101400300003005000c000c00004000cc0700000c000c0c4040000000c40d0000c00000000400000c0003004000005c0301cc0c000000000c3c070000000403c30030004000000c0c00304003000004000c00033300040040004c010000000000000cdc000c000410014c0c4000000000400000051f7000000000003004000101003d0043c00000000000cdc0400c01100000004c000c050003c007c3c000000000000fc400c004040000c0c400030300300000000051000c0c44000c005300040000040004004c00000003c0000330000000000000000c1000030040c0000400f4010c00000000c01f000cc000033004000000000000c00c00000400000000000004d00404030000004400000000001000040c70000003000c001c0000000c0000400000040c0000000c;
rom_uints[50] = 8192'hc4001000f044000c10c000000c000040000400c000d0010300303000000d010c0000100000000000000d1d3070004440003c300000000030000c0000041c303305000030000c0cc1c0000f000030001c3110c30040000c040030004c0c500034000000000c0000000000c0003000000c04000000000c0cddf4000000f3010040000000000c0030400001c00304000000000300100000040000000000100c3000cc0110000cf00010430040000c0074c0000cd0c000000c0c30000c04304030000000c430c0000400340f4c00004c04300c003c4ccc0d1000530000c00f00000033000000040000000c10000744000cc10cc00030000000c000000004400300c00100000005000ccc403c3000000c40000030400431000001c5c0000000100000000004c00700000000c40f404d700000003000030003000040400030000000000040300c010c5c0100000030100303374c0c7400000031300000000001440070304c0330040c00100000300c0000000044011f001040110000030004c000c000c00c33000430000c0000c00c0000c0040000c00017400f00f000000330701000000000000000000041000000c00330103400c0c0000000000440000cc00c00400001000c00300000d0003043000000000001cf0004dc0034303c04004000104000c003c000c0cc004c00000c00000100030000010000000000300c500000404400c4c00000c0000f00400143100000000001c0000c0d0100000c3300000c0004003000000000cc000030003003340000000c0c003c11000000003400000c0c0c40503030c000400000000300000010c0007c3000401010004c300d043c000301c30000000100c03000110003003f01004c0000003000cc00040000c000100001300030c0000000c0000000000300c0000c0000c00d00000cc00400c40c0000030030330314003411d00010000130000004cc000000000004cc00cc11033000000000004c0000400000300c00000400c0000d00c04003340100100300000000004c030040000cc0000000030000000100000030003000f00370f0c0030014c000004003003c000100000000100000704000d0000000f0000010000d000000000000004c000430400000030001000331100103403004d00100044c3030044010000000cc0000001004000000000000000007d004000000000000000c000c30f07000400d030030003140000003000030000d0030100c0000c010400400000c030400030003400000005c30330030c0c0000100100c00000011000000001c00000030003000300000000001030000f040004000000000004000040000000170400c0770003c01004400030000000000000000000000c400c0000300330c00c00000040000001410400310000004000100c00000c00c00003c304000100;
rom_uints[51] = 8192'h300c00001300010000000000000c0000000003000000000001030c10000003000f00030c000000003c0004030434001c100004000010d30003300030000000003000000000000400000000300003003000000c00003c34003404cc00101f00000c0000000000000400c00313030003000300030000c00003000030f000000400140c0040000010010c000000040004001500070000000001000000310c01000c003000000003000030000000c100000000300000000000500400007000000000500000000004000010000000000c0c00400000047400000443000100030010000300040030000000000005000000c040030000000000f0000001000000000030010000c0c1000c0c3000040000004004053000c00c100003000c100000c0100010cc00001100000f00040c400510000000000440000c00040000000c44101033001000010c4400343301000000000540030c00000404001410c0000d00001000001000c0040330000f00401004000001000000000000000040000000003000040100c033010000041304040d000000000000000000400000000f0000000000047000003404040c0000000000000f0400001030411300000300c0300c000000101c000d100100c0000000000c00000100010000010113c0000c0000040000000c543c000000000400030007000004000c000500000000000001000301030f130400400004000c00040003004340003040100c0400000400c0000000000000000000000000000034000000000c000000004f030000c00000000000040c000300000c4130100004130000000c0000000c00311000004000000007000000000c1703010000f400004000000000040100000001130100c00400011001000000c10d3cc000000000000003000c0c30040000300c0000f00004000000000000000000000000000000000043003001c1000c0100100000000010000000040c00040003000000c000004000300c00000000000c0000030000000010c0000003000d010400000000000000000000300001000000000100050034000c000c000c00000400400c01034000000c00000000000000000000040000000100000304000000500d0000000000010c010010000010100001000140c0c00004100000004000003500c00010100000000104403c0c0000300000300c00040000040c1c0000000000040400000000000001000c001c4030000400000003000037c3000430c4000d00010c0434000c000000440000040001000c04040000000000000003010100c000003000000701001405000c0400000c0d0000f40000300000c000d0000000000100000c0c000003f0000000014000000000000000000000000400000010000c00000100000000001030000c001c03000c001700000000011001f300000000000000;
rom_uints[52] = 8192'h30c00004000000000403c00000c00c00010c3c070d0c000050c0004c00010c00c000040c0000000070c00fc00000c40000000000000400c000003c00000000000400510d000dcc0000004000004000000000000f010000c400030000400000000000c0000c000003030404c0000d00300c000c000c40400000400000c040003000000c0c00000000000700000000000100000000000000000000000004000300c0000407000100000000000300004040030000000000000000040c00000000050004000000000300000c43c00cc0000004c000014040c100c00300cd300400c044000000c00000000c030000503003000dc00000f00000001300000000000340000004404c00000c0101000c530104c070f04c0c040c05c004010004c004c3c030c000c01040400c00400c0c04070000004401c000000000010000c1000100000400000c0440000000cc0000000f0700c001400c000530350ccc000c0440000000001000440c0401000014c000c3c000030400c00c0001400cf3c000040c0c0400400c34000003144000070000000000000f0c0001c001000000000000000040100400000000c000000001010003040007c00704c340000000c000000400470040000050000300030004000003000403c00000000d00c00403001000000000004c47300c300400040300000f004000000000404c00cc00000000000cc3c4c4040300030f4cc1000000000001003c400440c00c0040040c0c070400c4030004c000030000301cc000000303d40000450000c000000c0000000310000c0004c0000000000c000000c00304c0004000c00c04000044cc000001000000c0004030c0000003010f000c030f03000001000000010c000c0c000000000004c000c000c5470c03100000030c01c100f000000300cccc0000c10000000001005750cc030000c300000000050c0000000003030000cdc000c000000003000000000004c04000304400001300000000000c0000000100000004033400000c00c00000004000004000000c04000000c00000030000000010c30040c004040404c0c040400004000000031007c000000000000c00000000504c00c340040504000000000000030003040000030004000000000c0f00000000000c100c03000000100440000c0410c4cc004003c00c03d0c0c10001000001100300c00f0004c110000000c00000000000010004000040c00c000100104000001c00000000c000000400c304000c00404c000c0000000000440000001000400000000000000000c000c000000000070c0cc005400410000d0c00c000000000310c0000000c0300c000004c0003000c0003010f04000000340c133c00000500000000000040004004c00cc000000004030010004c40000c143c000f0003000000030004000c04400f100000000;
rom_uints[53] = 8192'h4000000040000515c000000400040c0c33000007003300c0cd3000434403000331c00000c0000000050000c50000000311401f10330c070c0f0300370000c03001403004000c030000030041c0000101030001010c400040c000040031cd030103003001001003cc00cc030004c40400010000043c01000d44010c0100030001011510c3000000040000c03000000c00030103000100400c040000130c000d00000000000cf10000000000000303f00c0c040300000f44f30000100501000c330c00000000c44f0f010030f000014100000300f10005000c40c370c3000104d0100007c4cc000c0000040c40400000030000341c0c00030000050d10040000410103100c014c4d4100030d1103030000f30f01013030001010000430000d410000c000014d04430001c0c007033d0000010304340000000307000304c000510100c300000733000c404403400010000c40c007000d100ccd0300010c00cc0c00c33001100030400d0100310000000030440c010343053000000c000000030030000000110c0001000000034400300d0000001000003c004c030000010040000430c1000100407000040c0c030344040f00000413c00d03c3040003010300030d04000303c0101cc00000c300000c0ccc000000c000c00403050000c000300c0300031700c040ccc0400d1304030030000c000c00000033010c0c0003030400000c0740000c004503030041051ccf0c00c300000c007110f430c4000030300c0100030000334301000307000003cc1000114000000c030000c303000000101300000fcd43000c00034000c703c3000f4003000100000000100d00001c00000c70000000c34003540004440cd000014110031004030003003104c00000c0c0cc00000303030c000000004001f703030c004c0d00034c0001000004014c000430c00c03000001010c00410cc071c00041000cc4010c30000c0003cc40300000070104104000000c00000003030000030300c030310c44100d0000000100050c000c00050030c000040003013c000000010400ccc40000000d00c70d0f00000305030c0007040c5c0047000c030410c30004030313400003000c0d0000100c0f0103001013030c443300410303c00c40000300c4010000030000004c31c0c003401040cc0c00c10100000007340300c10400c30000c00c440c0d404000000000000c0003c0007f00100003000c11000c0000134000c330c000010c00030003c30031001d0004000000cc00704c0c0c000003c0300000010300300073000c040004000301c40d0d0000030004000c340004000c0040000000c0000010000c43c04c000010040c17030c00cc00070c43c300c00000410140043f00000003000001d003000000000003000004c013c0000000cf0000000000c50c0d00130fc0000000;
rom_uints[54] = 8192'h100000003300c10040010000000005000000100000000f0000004c000c0700000000004030040000000010000400033443c303c0000000741000000000000000014001c103c100c0000004cc000000050010c0cc040000000301000400c00100c400cc1f000100000403000000400300010000c0300104000004000030000000c4400000010700000001000000000100000000000000010cd30103100100033000c00300000373010100030001430401000000400000000100d4cc04c400000701c10401000300c14300030010c0440000140003000100001000c01100300001d000000304003000004000d700700000101c0c15000000311301000000000004001401001000000c010000000000000400110300030001030034000d0400041000040000c04300000000300003000704003f0d100500040001003000000030000c00110040c004040000003c01d043000000c001030003cc000010030004c07c000310001017030c0001c100100000000000000000410c000034000d0000c0000300c404400400400400400004010500000000300c00430040c030000100000000f4000000c0000c010d004c000101000000d04cc31314000001400040c430f04c00f04f0004003400004c00300000001c00f00c00010cf0000301000000007700103c000000300000000301030c000c7500000000000c0404000003300000000d00000000000c0000400101c01400c013c0034c0c00014c3c003401000304040000000001000040000000c0030100000113000000410001347000000400c0040004000300003000000400040000f40010000000110030030000010000000c10000c14003f000c107c00000103300500f300100140400c01031030001d0c00c40000000000c0003c000010000100000004c4330000030004000c00030000100310700040c10030000440010d0cc1030100c0140030000030040003100000000c04c000c100000000c03003004000000c00c00000300000100010033c033000300000100007140001000c000400040000000004404001000010c000004000114000003c00cc00000100000c00000000c0000004d0410cf000304003c100000104000300000000000d400c0301000000000000030440140000003000c150001003000c030000000f00041000c00000003000000004d403001c000300000c0100c01010010000c0003003300000c0003103c00401d00040040041400010000010007401340c01007000000000004004100004000c000040d00010100040100c00000001000000000100000000000000300000070041c00000000100010004004000000001c000c0010040000000c77000c000000c0300010014000110007103100000000100c0c000000cc0030003c00c00130300000c0000000000000c00001000;
rom_uints[55] = 8192'hc413000010d03c000c00000c1010d0340004c00404c0310c00cf001000400401303034c000040000c030000040000040f00c0010300c001404c00300040c00000c030500000030c00000000070001c000000c00040004000c13f000000031c00003130004000c00000301030003c00305100000c440110c404000000000000300cd0700100dc301c0300003c0000c41000040000003000301400000cc000407040100000c0044c0500000135111000f30034c0c100001400044c004433c00c0010140010000031d00c1500d0c00450300c40c01c400c0004041104104030400000c000300000310000c40043344c0000c403140f0000001030003000000000000340030500014431000034404010330470c0340030f0000c0c0000c304c04c0000731000000003fc003c130040005c30030000004c440313c0703f34300040010c3400000000c710040000fc000c0000300030001c31000011030150070c030500700310440c33f0311100f0100040000000340000c00c0000000d0c1400f3c0103c1c001c440000031c040c0cc03c701000700c000001000110300000001003307f3fd100f350001c3410c01410410000101000130c00d31000cc04305333040000307430101c00004000000c04101cf300300000001503007000000400100c0000003000430530000001000003c000444050d0000c34101cc3001003c000300c00301041dc0d340300541004d0000030c00c30d00300001f00141400335c0140000000704010cc000030000401030c4007d13400dd14f0c03011003000c473304004000300f400c043f00f030c000000131031000000007400400000300c071d10000010ccd0f70c000c00000c51c000d01c741c43044c430040041cd1d00f1c40c0000303001c30304001010007d030100c341000c1300001c000c003000c3c4030150000dc50000c7c0010400050c0fc400104303400430343400134003c733f0f0000000f04403c0000000010303000100070cc333000040c0040f3c403010000c00f03430034444004000001f034313c0c0c3cc0000010700d000d3304300003047c0c033450001000001003c00010440401c013000001c0101010404410733010341df0c0fc000000c000c00004003000330300010400100000005003100c00050c04003c300f000000001030403c0000103f000cc030c00c000f0010c003c004301c100c00000001410000f310105c0c000453003c00000133103ff0430010c00f00300000c00000c1500000d4310030013c00004c34d000405c00333000740040001c130000330400c01000001f0030f00003040000000000c114c130d1004f00cc40d000000d1c4430c0040000010030044000430030f10000000c100340f0004304c004000000c170c0003f00340000000c3014000070f0c0c000;
rom_uints[56] = 8192'h5140c0000000000f0000000040050000000000000003f000030c00000f0000000000c50000000000c0000000c3c000c33c00304c000300404000040c00001000000030000000000000000010c0040113700000c35110030c30d040c00000004000000003000001001c040000000003c1000001f1110c0040c00000301000701f300000300c4000000c00300c1004730f00400000000c0000300c30000000c0cc10c1c0c000000004040303000d0000400030000000010400000000cc004003c00000040000000000c010000c000400000000d300100c000100c0013014000000344000c00000000000400c30013000014000040c0700000004000c0c001000003100010535001400000005000001c0000050d03c0004000cc000010010000300c0c40000000000300000411301400100400000000500000030000031000010c030300400030140003fc00f0000100100c000000000004000d0000c000000001100c0004031000030040000003010000000003033cc34ccc0000c10c30010030033f3000000c100003000000000001000400000c000000000000000000000030300001400031040000100000001000000000000000c000000000000000030030000c000c00c0030003405000400001000100000000030301040010014003c0010330001c00c110003003030000c0003010000000000c00000000000030000000040000000000001000400000005000cc30f000c0c000000000005005010000040c03300300400100400000000c0005000000000004000000001c00034000000d000040c00000f300013000c13004000000013000000003005001000000001430000030011300003040000c3cf0000c000000001c0000c300000000000010000100000000c000004f0dc0000001070000000000100010c300000000c4c0000000014030004000c01040c3000c40400140400001004c000c0000000000000000000c004000000000300c000cc003100000004000000000cc000000c000000c0000000000000300f30400030001003c00000000000000040000030000400010040031000001000000404c00000000c010000000f30c000010000040304103000000400000000c0f07000040c0400003000003030040c00100000000000004400000340001001011030000000100000040030001000004000003103cc00003000000030000000000005c0000000000003000040003300000404001000000c43001003000550000000000f10300030000104c0101100c00010c00000300000c03000000500100400044300000000000000cc00040030c040000000014000010c3c4f00050f0000cc0010300030c00c00300400000000c0010005050000100003c000043004000003000104100cc03000cd001c30000000000100c00c0000103000000;
rom_uints[57] = 8192'h1c000000000000c040000000c014040fc00000340000000031000c0004300000000004040000000c1000040ccc01000c00000c000000000000000000001c0310000030000004003004440c000000010001300c0003100004100000000400070107c010101c0c035d0030000c031004410000c4044000c00c07400010c0000330000c04400000000000000401000000040000000000c00f000000010000000d000c000c000000100000c0044cc00c300c030000000c00143003000030000000c5430000000434040100c00000004000000000000740c0010700043d001000000100000103010c03c0000300101001000000300050000010000000040000040c0407000004c000040004040c0cc000051000000034c4400c0ccc00300000003310040000c0c010c0040300004003c440001d00003c0000000001003d003000040c10100d004c0000000004700c04000c00000403031004340000001400c00d0000000003000f030004000130045001000003040d040000000400000010000003f0333003001000000c000000100103d10005000440003400001f0c04000030000374040003000100000004030c0c10000c000000010400003000330cc00c000300f000170000000c0c00000000000001300040000000000001000004030470c05000010404cc003c30c3f11c0c00300dc00003007300040400c3050c04000000000c034000100400000310011c00050000cc000c14441c00c0ccd0010003000c0001000104000000004000000004040000d41000000030000000000c00000f4000c0030c000000000000010433000000100400c40003c0000000000000003c0400003c00c0000010000007000c004000000401000000100c0400cc15000404000000003c0303040003000c0100c070000300000000c7403000000307101000c4c33010001410c10140c70504c00d30030cc000000c0c000000030000103000000c04140000000c00040c000c1000040c100404c1003000c0000c3c00000014cd0000000c300000000000040010000003000000330000300000004004000100000c00000000c005310000000300000000f00440440034040303030300001000000000000d03d003000000000304000400c00033ccc100000c30c000000003001c1010000c0300000000300c0c3000d400000c0010000000040c0d0010300c030c000000100100000cc00000010001003430000000300304010c0000000c0d000734000f30000010000130000000041410000c001c440100ccf00304004c00000104001100100344000000000cc000101000c3000300010004140140000f3004010c0447c30000174d0400000c000c0000403000100400347000300000044000140004000f3400003000004cc00c01000030033000000300030004000c3c00000;
rom_uints[58] = 8192'h100000000000000c10010000000100400000000000000f300100001040003000000f1000401000001300000000103030000000000003000000000000010000000001003010000000000300000300004400000300000000000000000001000d4c0040400000030400000000000303000101000000000000000130c0004000030000000000000000013000c0000000000000430100000000000000330000000000030000000000400010301000300000033c0000003000010030003000003000000000c00030000000010000100000000000100300100010000000000000000000000040001300300000010000011000000000000000000000010000001005140000010000f003041000030003010000000043000000014000000015000003000000000000000010c000010104000050000000000000000001000010000c100040000100000300000101000100303c000000c00003000000000c000000003000000000000301000004000000040000000000010d0100440003003003000000330000050000000000000000000000000000030f0000000100033000f000000000000000010000001300500003000310c300010001000000003000100000140000003000000000c0000000010000000300003000000000030003003c00001000001000001000000003000011000000000000000400000000000000000000000003000001000000003c4c330030000000000000000000000000300003004000100000000000040000001100300c00003000000100300c00040000000000040013000000003000030000c0004000000000000000c00000010000c04000000000400c00000c00000300000100000030003c0004000400c040000000010300000401000000000000000400040c10c00000110000f00040000000000000000000000000c3130000000001c000000000010000000004000000000100000000000000000000000000030000c0001000000014400050000000000004000300000000000000c00000000004000300000000000000000000300000000000100000040001c1000000000000000010000000c00003010000301000040000000310000400004330000000004000000c00000000c00000000000000000c100000000c001000c000000000000003300d000301000001300040000c003000000010001000000100000000000000000300000000000c0c03000d1c00001000000000000341010010000c000000000000003000000000000000000000000401000100000300000300010000001c00001000000000001000315000010000000000001000000001000003001030000000000000004000000040000000000040140c000000033000000000000000000cc000000000001000000000010000400000400001400;
rom_uints[59] = 8192'hc00010000000c000c00000c310000c1c00000000000c40c000c000000000c00c000000700000000000040001000c4c00c0004000300000104000000440000000000040c0000000001000000c300401100430c000c00040c0400004001000c00000000034404030c00000000000000000000000101cf000000000400000007030c000000014004000000000f00000004000100040004c00000030400000000040000c000030d0000000000000007000c0000c700000004000100000400010003000000c000000004000d000300000d0000000040000000040000000c3c00000c0c0d00000c00000000c00007000000000000c50c000000c00000000403000000004000000043440104c0000000d0000100ccc00001040c01400c000c0004100c0004040000000000000c000000014c400c01c0000005d0000c00000000000100c000000000c4100000c4030000000000000000000004030f0c400304000c000c00040c0004030c03030004000000000cc00cc400000cc0000000000300c1000001000c010d0500010003050040000cf10000000000040c000000000000000000000c0c0000030004000300004400000000004107410c01000000000400340330000000000c0c000400c0000c0c0000000000000c00334c33004c0000000f040d0000100c0000000c00400001000000000100000d0c00000000050000000004300000c704014000040000040500000004000401000103000000000d01000000040c11c4c00000000c000140000000000000000404000c00000c00040000000c030c0000000100000c0004cc00000000000000000000c4050040000000000000c40004000100c400400000000000004103000440470000040c00000004030c000300040041000000001c03000c03000004430c41000c04000000040c004003400c0c0c0001c00041000c04c01000040c0300030c0000000000c404d000000543000000070000000c00000000000000040004410c44000c0004c70000001c01040300000c010000000c0004000000000000300000c300c000000000000003430300000400000f00040c000001000003040d0c0c0504000c0400005c0000000040c403040000000100000000040040000300040701000cc3000000000000010000000d400001040d003000cc00000000000000000004000000400c400300000000000c0000000000000400c0000c0400030c0000000000000c0c0c0c000003c001000c00150c030000000140000400000000040000000300070000000100000000c000000c00450000000000000000000400004c014000004c0c0004000000010100000000000000c4000c000000c4000000000003000000000c0c0300000c0000000100000f000300000fc300400d0400000c400c000c0c00000000000c01040000;
rom_uints[60] = 8192'h4000000000000404cd30040c07000310330000001300470c00000c04000007001030011c00370000040000130c03300013000f000d0100140c031003000040000430314441003000000005000400c4300410343101c00300000d3c0000c03d00000dc01000000010301003003030001005c004030471003000003f40f00cc30017340d0f000000013010000d0000470000000010007030003f041c0000000011100010c030c000000100070333040030000000040000c000041000c01100000c33004c001004700000410c00010500011000c401300c1400404c00010003000000000c0c000010030003003001d0cf4170000300000000000c010103cc34003c073c0c300fc1c40000003c0c3017c010c0030100003434000030030d00370c000001cc00101300050c000331000401001000340c01000c0000000030c1103000c000f311001003100030000c340030130003000100030d0c01003000000004c30000ff003c000007000000104034003c00000330003034001014140c00000043000001000030143043000000000301c0000001c000140000000714130100030000141d00000400040c110c0033070000330000300000000000c1040c00300014000510003100031100000700000034043100100000c0070103c00050040030cc0140001d0101070c0103000000000000040003030303040400000040303000000100110f0300104713300030373014c00000000d03003404040300003453f00c300100c000010010000c340c4d00f0c10c000000040c031100010304c0004001300030130001000000301301015001010300000400000304004c00000000074301c00300cc000031340c00000d000004f0030f000fc007010d310f300c00001c00c13010c0000100300c0c5730040c00010013000c004000000c0c4037010cc010100f34c000c00031000000c0000c3100330010100c00000000131000110110c504c0310000000c010c001000c10000100410030001000001300ccc000c1000c0000104000c001500d73140010c10000010000d1337100000000000c1300f0011030301d10010fd0000140d00300c0300000000400110000001001c04001c0c0305000340000003003033300000d00003000034000c0300c003011d03003030cc70c03000000300101100011d004004001c30000c00003000000000000000150013070d00070000030400000d1330300c4c300314330c001c0c00003c01d1000c0010041100040000000c30000030303730000053010000003c3030013000110c00040c0c4370c00430100c0304000c0000100d1c0000c0000d0c00110310030104714c03050030140d0c0004000015000000001004010100003100000c170544000c000404000000307c00030cd00ccf000300130f00040000001010004000;
rom_uints[61] = 8192'h443000100043010001010100000003010000010c0001000100000000000300000100000000000000000000000000010000033003030103030000010334100003000100000330000000000000410131030013003001001400000030000303130000010111000000000100000300013030000000000000000300031331103000003000050000030000000001100000000010000000000030010030010004000001100001000100010001030000010000000070000100030030003000400000000033c00303000000030000000010000c0500343030000301010301010047300000c003000100000000000500000033000007033f000300000300000003100000310000030300013003000100100000100000c300030101130003003133000030000000d000000300000010100030003c000000003000030000000000030104030000003300000307003001000c01000003010303f00000040000330100000c001301003303300001000110000303000130030000000330000000110110000000133000330300000000030300000000000500001100110005033f00010300010000303c0000000300000000000003030700000300c3100100030000001001040400000300000000010000000000010000000301000000003700000103000000000040070000000100000013003000030000530003310000000300000000030001010300040300000100030100300017000001030030030001030000001f11003103000003010003030000500103410003000700410031000300000100000000440330000000430c030300000000000001000013010000030303043000000001000000000301cd00117100000000100000000000031303130111000310001010010c010001410000003301000001110d30030000c11303000000000003000300000133000000030100001433040001000000000000000000000c03003c0000003100030013000300000000130000000013100101030000010001000003c100000010000000300000030c000000003000000000131001000000000100010000010300000100003d000300100001000003001001000303c10000000001cf00010003030441000300000003010000000003000001004100000003000033000103001003330101000000003030000003300000010000000000000033010300000000300130000001301300000101000141000004001410000004030300010000031301000100100c01000c000300000030000000001000000110100040303000050300000001030101030310000300000100100000130040300013000000100001030300010405131300000c003101030300000000130000000000030000000300101303000000007000000f000303000500130303000000000001040300130100000000;
rom_uints[62] = 8192'hc000030001000000000014000c00030000000000000000040c0000000c040000000100cc0000000000010400040c00040c31000c0000c00000001000000c000700010400000400000040c0040400000c40000400000000040f00c0700030074400400c0100000001000000000c4100000000040c00000000000000000c00744c001f0100000000010000040c004000000000000003c000000000000400000000000c04000004000c00004000000c00000c000040000001000000400000c0000000000000000c0c00040000040040c00c004000004000c00c00c0407100000300000000c00000000c40cf003c00000c000c0000c300004000400c000000c0f00000000c03c400500007c0030d0004001000300010cc000310000c1000c0040050c300c0000004c000d00000c00000400c01c00400010c000000000c4300000004300c004100000c040050000cc00c000000100000300f00003c000cc00004000000000c04000c0000014100000c400cc00c00044f00100030000f0004000000000000c0c410000c000000000000050000000044000c000000401101040000033dc50000c000000001ccc0000000000c00c0000301000000000c10040003000007001010c0010000010c000400000000c00100c400030000040001000c00c100000c0703000c000f0013040000000004000f0c000400010c0000000c00000400004070001c30030d00004d0c03c00f00c000400c040000000004040300dc0404030c000c30000c404000100c0000c000370000000000410041cc0c000031040000100c0005110000000103c411000000010000000c00000034000c0004400100000000d00c04c00000001cc0001c0004000c530c0c40000000000003000000cc0700010c00040c0003040004000000c0000000c0000f04000c000013007c000c0cc00000400100300c0cc0cc000403c00004000000041c10001c030c000c00010003000000010030c0000000000000000c0010400000004c00000f100004300000040000c00041000000154000c3070000f0c0000c00000c00030000030f00c40cc000010300340000000000000c043003000040000000000010000c00c000cc0000000403404000030c000000000c0c10300000cc0000000000c1c00c00000000000000040000000503000000000000c0004c0141000c000030000c000000003c1000000000c0000100001000040000c00000000050c045000000000000000000001000000000040000034cc0000000c00004030413000100cc000000000000000100d40000000f0c40003001040000c00014010004000000000000000c00044003c001400c0001100000000000000040000000000400003004000004010c0000c000000100000400000c00030100000000000d0000000044033100400000;
rom_uints[63] = 8192'h5001000141000343c00040014000c430f0c000010334000007c04000000c000003f00443010000c004c14040500301f340014d030c00000040c000010001100f0001c3300000010000000401003c0dc00310c0000410c000400400044000c1400003cf0c10000d0000400000000147014400304101004030000100030700000100047044c100014040400000c0c00100010001100011c3d100430000044000413000010300c3c010013300501100c003003c0100003110c000030034f340000d000000000003103110000c0301c13c403100003000d00331004040101300c35c040700c031c1c301433300400040c000000000701400000000003140c0004331c0c000000050444000004000001000030000030000c300004100003000f3030103010001004003c0001cc00340034003000003f140000003000007f00c450040f0001300001131030000034001000100000100410100031100104c4000c0c00100c000343353010000000f43000113c1003000c00ff00000014cf303000000010431034301c1c40c330003c11001043c0000003140004004003003300c000000cff70000cc0000c000034040510000c0014000c5cc00c103300c4cc04d04c33400000010c00101000130030000003000c00400c000037dc04700c0000101003000000c1044010301c040000044030ff10c00c300000300300cc0010000c0003cc0030003c0400100411301400141d100000443c000510c0300000050100c0000d0c0000300000c000040c4005000000003004000031500050c00000000010013000143030000303000c00303c0c0000001030000000cc030043050050000c00d0001000404f000000100000030c0000100010510400010030004000f03404cf333d000400000cc03c011010c100110030100f1000c0044000c4000411300000310c3407000000005003103d04000070c00430000000c00c3c103c10c000c30000003c0000000037d00c3000000000100007300d0cc4044000300003003c003d0300003333000c00004c3010050400300030003330c0040c0000c00030103c1400c00010303c007c100001040000000004303404d4c00030300000c0d014041f010c001300c400400010300c0000103010000034301140040c30001c043144073130300403003d300000100c3c40100000f0c0100040003cf03c00000000c000c00400304313000c3000000000000030001400010010003030f001000000343300000c00c000040000030000300c10101c0c301c3c3010c0c4041000003000003c000004101cc000000c00015400100c003f000030001c3c10000c000003040000040101000ccc10301014100430000400000c003000001000030130100000301000000c0cc000007003330cc4004000fc0040040000fc300c30000c00103130;
rom_uints[64] = 8192'h410000041111003000400000c0000000030400710c3040010400300101d0c05c0050c0113c0005413040104000430374d4101f00430000c40c0c003d000030003031d030410000100004130140010d4300cd01c3330000c1404000c000c340003000030000000040000300000f4300000000300000f000c34000077030500010403300100030000000000100000000540000000000710041c00100003f000c0003f00000400440d0000013c0501300044330000000c044c3000001c40040000003013100430c710303004303303034003000400000000c7f0c0004001f404000000001540300100005c0303504140003041cf030470000300130054004000c40000010000303007100051c0001c041040cc034100301011001000cf3f0400300411300000c0007c000001330c000100033300111c0000140030000410100000010040310000150000050c010c5007404f101500d0c4c471cc0104511003f03c04050d0004000300030c0000010701fc03070011007c443c0704053c0300d0000f40c00c50010004014c0c0000c00011300000c50000000000310300f000400004030305000003004130300301034300030050c30000c400033f10c005113103c00c3c040cf000030dc00c00c10140300d040003400041040030030c3040513000c04000033301343101c01000c03c3ccc000c110013000400000000703000054540130001103003000010d000340400c041400410010c0440003133001001040000c0000130000c000c01fcd050000000c0f40000070c003030000403001c0400c447fc0c041f003cdd00f00440c00100004130c4040c000035031c3043030c0374c001fc07000340040000001c1300c001035011040000330c3000330030c700000c04040403313d4101f03000100314c03400c0c400c401f307000000001000f31c000c0400000004c04030c1005000711504003300010300141000303000010510000d0011000030000100cc00c040d011c4000007c000000c30003c000330000040c4400ccc10f0313c0c003c70000003440300000000003301300341c011003400043c00140cc0000000df00000701000130000030c0100d3000000110501104040041100330003000030c000031100d01004300303c013004400000101c031100007030000400000004430000003f00c003c5c00c03cc4310050305104100100000013040c0000000c00001000304c7140c0c0010340c003700140c47cf331300f00005043040010030ccc004040c003000fc0c00d001304400c30c030010c400030404011103000001000c30003330c0d1004003000c000004400304001f1450c000d00303004000040c000003343330000300300101100100340444f00c000111c301000c041c10030d000044c0000030300f30300c00000c000000;
rom_uints[65] = 8192'h14300000000c5140c3000000400100c00000c0c0000030000100403010040000000c30c1501c0000401040c000c010307cc300c54303c000c00000404000c03030004000000000d14000c0000330013003004000fc0f4030f103007000c000043070c0004000c041000cd00001c00c303cc170017040400000030000c00000103010c0101040000100004000c00040c040300000000000c34700c03033100000c030c00040c00351c0301043100300140030400000ccc1400010400034f0d0cc0d11000000c0ccf0303c400040000c40414401040010403000440400d4730000c0000000300050000000000000c00000c030c1303003000c00d000004000000033c00040c140c5430c30437000010000700c000c04007000003300cc0c40004300440000c4000000400000c040013c30010000505530c00050004030000430443000d000001347004300043cc000c0f0c0010001441037100d04d3c140100dc0c0d4cdf0f0d000400043d10140000030043300300c0c00000000c0530000000004300300030300100cc000003000c0f7300000c000300400701c000c00c0c0004000300040010004003400005441d0c31c30c000c03470c0c0c07fc0001330f000c030400f00c00dc0034c0030400c04100003c0c070407000301400400004f00314030041c0c000f0300000c000003c5c30001400c001c001c030004334f440504c04c0d000130fc0704c004c3410c0000100c000307c301030c0c000c03030004051c00034047c00c040004000d0d0c0334100c1400c040001d0030000c11c00404100f00f000140403f30c0cf100000d10000c0510cc0040040c004000000c3d011c01040004000000000f01041033000004310010030fc1104034000400cf000c00cd00003c0c00041000030103000400041c1f0700c3000c000dffcc0000dc0101c100c7130003404000000000c4040000dc000cc0cc000fc00003000404000304c030010303440c00400400000c05003300033c0c44700c0c130f101d104003040c340c00000d03c0010c000c030f1000000c000000000401010100100f3c030043013d003100000003000c03000000100cc000100404c4040c0cc10f01000000000000040000000c0c000040000c4003030c000430033c00400400440c0d0c0f0000003c4001400000071c00074004000003000003d430000c400300030d01010400100c0d4000140c70000c3003014001440007c7c000034103000100f035400c0000c300003000404300000400000c000ff00c1510044c050c000c0300101c0100000c05000c03cd4400700001010c010003010110000000000310010000400c04050000000c000cd00c000000010300040037500d0c04030c0404000c0400000c000ff0030510011100101f3000000000140000000400c0000c030;
rom_uints[66] = 8192'h1c0000000c00c40010000000c00000407700c00fc0030000c0c000c3c40c00510fc03474c54000cc37400c400300730f004301000c400f004103000030000cc00d03cf0c103000c43000001c40c070000500d0014300d340000f00000043dc0d0f334c45cf000f000004400000140cc30000044703cfdf0cc004ccc00004c00c00000c00400000c000c0000100004000c0000000000000000040c004001100404140400c0003010d00f04c0140040fc00c0c040400c0000c0300003000000040c40100000000040c0cdd0040030701ff0030f40cc0c0000000030330f0d000000c040000c1000f000345c33d150c0040010f0400c00c000000001cc4cf040014340df144400ccc404f03000c00400c01cc4c000500040303c00304dc30004040300f1000c0310004c001cc00cc001c0000ccc0c0c1c010000d03f00cd3d30000ccc1700c03c01d1000034003500030c000c0040c4c0fd0c103004400c30000030c13775003dfcc010c01c00d41300140041404d000c40407c10c7000000c000004405c03f040c00d014d000110040173c000c40000000c00043051df04000000104540000dc0400000000000001405300400d1040c03c0c0c30003304130001001cf00401c000000050f40004c000040c34100403000040000030001000000000000410001003530004c400fc3031401cfc0c070014c04100004c310c00007d30100c43f0001300100050053ccf00f0f40dcc00000100400040040c4144cc0c13400040f000c010000ccc000034c3040c50000004470000000034040000003000433c0000100004000000070005c40c700040f00000003c00010040040d0043414ff040400030c0f00403040000000440303cc4c0307c00000001001000734000c414001441c40dc0403c00050c0c00303cc0f0c000f010c000700d05d41400c01000104c0df000701c4503140303f0fc0000013003000cc00003000c30314004300440c0000cc004c00c00c000010cc00cc4000c3f10003100400c0740400500c0000010c00410000000013010c010c0000037d0000000c43004041c0101000014304400c0001d000000300300f00000000000c404000000c1fc700400c000305000000000f0001334700c0074c40030000004d703403cc0350440100414040c04400c70400034300003000140cc0040341c34451c000440001000030cc000c340c0140c04c0000030000014f000304010c0cf130010304c007000500c040000c10000000004c00c7000004030003c03000000301074000000134c0404300070340c003731c0f030c0c4c0133000030004000000100000000400c000100000c0c701c0c000cf014cc400300d0440c400340000000344000c004001c00c3f0d0c013c010450000100300000301000c0031000c00000007040000004d400c0040;
rom_uints[67] = 8192'h100000003005000003c0300d3003700010030000cd030430743400301003430310170c0cc5400000c3000101004344d01c031000d130cf00031003400c500410c430010001c030000000710000cd00ccd004400f00dc010350101100c4d030001c040c050000000000c0000113400c003040cc13d04400000001c501033003c100d100030000140001c0000c00f00d0000000c00c100000400100c10004c00040300000000400000010030d0311c0304013c00004044130f4400444c00034070d1000300003400000740401300004000d330000000300403c40001100c040000c0000fc1000000000000003c414103000c0441010000f30030043100000000c0010030c530000033c000c0307400c4cc704030c03c40003c70015000f301cc00040c000135000c001730d0110040010431040cd0035303700000030003400400003dc40053344031100000140310100c300004004007c54011d001000f000005030001c04000c000c0c4000301011000c300000f33034d00c4000f00003003000040c0c400100030000030410403c3300003000300000004f3004c0100f50000430c00040010f070000000003c0000301035f03030c10000c03010100140404cc3000c4000010000d400000000010043c00f0010013007c00c40010040c011d011000004007d0030313c01300000003c000000400000d7c0300c003307c337000c14d1c300c0000004440c003033000000003000403400f0c0000cc0040503c004f03cc3c001000011c0c03000310f00040c0000c0430400401000cc0001030033000c0040404000c430411010000300f001300410c300001000330040040c0f040130330300010040c0000030000001000340003c04300f4041000030004031c0cc3040000430c01f00003f0c0000304c0031c30c0070000000047004100040000000c03d040033d310340000003740000000000100000300003000030103c0300041000000101000100000c710700030c03000300000030c004100040c03c4003c00000000040000330004000401031041057001000000cc0000f431440040000f0304c300c41c00000c00010003040004104400003001410101c1340001013000004000c4104130030400011d00000033c0041cc300000300573004d400000d00050f0000004040c100070000101000c000000c0034070cc1000440c00004c0404f10c40041140c000500000c0400c7c1001400000cd000031440d00003530f40cc40007000c00c400010c01400030c30000f001cc047004300100d104c00c003330d0011004003005400300000000000114300010003300000c400cd00011014110c00130000cc11010c1000f400030c43000300c00500003c01000130000000400700033000000340000031000c4100430050c10141c1033403000100;
rom_uints[68] = 8192'hc040c000c0c040030003003004000004000010040c000c0c004040c314000c00000003041004000000030004030404000cc400000010c0c4110000c143c0000040004c40030000100000c0c0c400040004300f00c4c4000003040000c404001c00000c04000000000000400103004cc0005c1c4cc0c0400000300440c000c10000c3000000cf0000030000000300400400100004000000030403040000c400000000410001c40140400440000c0000000003010000ccc440c000c0cc000000300c40000000c0000c040100000005000003000000004d0000c3cc10c30c0400300400000cc07000000043c0300c10c0300300430103040000c0440c03c00000000440400401c0007040c10100004000000d403001000f00000034000c300c00040000c00000c00c400103c0000000003f0000c00c1c0cc0004030010c0fcc400c4d00c100c0300000400000c1400000cc4c00000cc330001c50340400000001c000400000cc000344004041c10cf0340cc0000000000000c040c0000c0000c301c3c0c00300001c007c4d0c0000004cd0cc0400000000c004c00300f3030004000040000300000c4100000000c0040000cc001000c00c4000c001003000010001000cc000410004000000000000000c0040040004000050000000cc004040d00001350104c000c0c000010000130f400304c0000740004c0000000000c000000c0cc000c00040000000030c0000000500000c0c4003000000000c00c00000000030c0140040cc040c000000f43040000001c10000004000c000033003010004000100c000000000400000400c000300030000010000c000cc000c40001000004444000000300000c000000301f004000030c000d103c10003c000c0000140000000000c0040000000c1040000000000037cc0f0000004ccc000000000040004c001c1000000000c07c0c740310001404005c33003c00000003040041303c000c0c0000041000000000700000000000c00004403040000c3001c00000000f00000c00000100000000c00c30003000000c010400c01005000c0000000000c104c00004000c00cc000000000c000003300004011000000000c000070c04c4407c003010000000c00000000400c0c030100c00000030100010000000000000000d000330000000045000c004001000c00000000c000c100c7000f500000000000030000000000030c040000c0001c00c304c0c000c0d11c0cc000000f000000c0000c03040041000070c0c0000001c0c0030300000400c00100000f40cf00c303403040000000000040c04000000c0401c10c0007c0007300c5000c00110000010f030100050013100f030000000000c0004cc00000c300cc00c0000004000000000100c0440340000003040000404070000000000030000cf0404004000000010430;
rom_uints[69] = 8192'hc000000000c440f0000000401000c00000d0000017cc30100033000104d400004c0100503040010043c000000c0140300c5405d050d01000100013040300100000000000400cc040400000c0c004c04400c00000404003044f40000030000c0004cc1003dc0000000c003000c3004c3034001030001043000c00430003041001c000041000c00000000433d0c00035f0cc000400000000470c005300c03000c3100000c03c000310040000c4c430d040043000300c00c00c40401437300050cff4001000000300f3003000000000000cc0140000041000dc7410001103300300040000040300001c31f000f00c77c003c50013034d4000001400030000400c00c0301404377400c000000300407000c4cc4cf0000c00c000c0000c4f00301000c000c004000c10300010c0c0000340c1c13c0530c0c0c0000010700310500000040430000c1f000030010000400000c40000c000d00050c03010034300c300704c0000073045314000403ccc10f000300300c3000040c0ff3f50c00d00000013103340004003c007c0300404cc340043400dc00c0000000000c00000cc03030c034030005000010040c05014000400c0f1000030f0404000030000c000d07030000030310c7003000310d000000030cf00c000d0000140d0040000c3c00003d4441004000301c070101331f050c001d0700014743d000c00c030004f37cc000300001410c0400004c100030003101010000c40333000301040c0c1c000c303c1300000c04010dc000500000040500040cc000000c010c000c03010c00c000010c000c0400110c000c0cd00c104f0d030c0007303f4c10c010c01000001000030c0300300f000000410000f7c00004040c040d40044c04000cc03d00700034000040000c030003000cf00400000000d0305340000004300300f000040040c03c0c4c00000100c000000c0c5f00413003000c043400cc00fc003000f700c00000c4040f0400000100c0000000000003000034340300033f44c00c04000300100c0c000400f70003000400041f0c041040000104cd0000300300000400500004100c0c00cd0c034ccc1100000000000004001100450c34033030040000000040014c4000003c44100c00000f0000030c0000000cc40c7430000c004030c000101c0400c0041007c040f0010c00c000010d0400010000c3003000000400000f000c04c10c0c0010044c00000c0c0d0010030d04010c0010000000040000c3410c3ccf0000c0c00cf0014d04104700040c030000c00400004100c40040001c0000c0c70300000034c5c00300c00c00004c3c0c140000c000010f0c000d000c00cc00000c451d00000c700c00304cf0c00000000003c00000001504040000c000004100037000000000c00013004004003c00700000040c0c000303340fc410000000;
rom_uints[70] = 8192'hc7010c00c75005000001000070000134c5500f34000c000000c31000040000000001001000100f030000001c0000300c03400c040030000310c00000c000001300000100000003c070010c0fc00c31001100111c0100000fc01c00c3000351003041000050000010c000000c001000304c0003f170c004103301000cc53030c300f00030000c01000c00010000000000300000000c0d0c10041000000007010c04031003cc0103011c04000400004f30000140000c0000c74400030c0c0000140c10000d100413030300033030110000f0f0000501040000000000cc0400040c004000000330c00000300c0f0d00100c10073c300000000c00000c0c100000cc0030144300c010114000c010000003030013400cc00000000040000ccc0100010000000035000c0c000d00c40540dd0f3c000310f40d0000040c3c0000311fc030cc0010011004003cc40000300000000cd0000400c00f00040303300c0010c000c0054330030431344100040030cc070c00f40c00040000010c03000c01014f0000030c7c034c0cd000000d010c103000000cc1000cf1110f0c11040c0304170100115000c0000310104cc433030004101040147c0d0000040c0000000300100300000101000d1000070004001c00031c00003f300000100f300007000004000c1c0000c0311c010cc00c50040400cd0c0003044000010033010c3100300c1c400000300000c30c1c04c003000ccd01010c0c0300314c400304034100c033130cc000c0dfc000c01003c004100cc00104433001004c01000c000030d0000310f1131f000c010000030cc10dc4001000001000c00c04300c0cc00410330430000c03040400000000030100044700040c03330d3c1c0c30001001000c00005d0000cc00c0000004f01003003000003000cc00303100030cc00740000000100001c330013c40333401d00d00011040030c00001400000fc10c0c001000130c00000cf00cc30000d0001000001403300000c10c0d07d00c0001000430001400000c000c13030c00010001d310003f000f073000f0d001000000c040000c1730140410000c041110410fc0031000c4000144044c000000c0101000000000cc0c11300300000107000400040fc417000000000301541c00000c0000004c100c044144300c14033000010103cc040453c703040c00040c0004040c40004000054c0303d00004003c0000030030430c5003c003045300103030300c0d30003ccc00000010030400c000000c0000c00304000400010310010150c30030c43c10c40030000f0dc00c0400300004f003100d0c0000007304f1d0000c00c000000000430000003503404c30005000000450000300000003300000100c0c01000311044c10014c00040700000010c00000000007000301000cd400000300040111043000030;
rom_uints[71] = 8192'hc5000001034d030cc004030500004001330000cc0001c0000000c0004f1c01c00000330000000d000f000f000003000d0c1140cc0347003d000c0c04004000040407040041c0000c0007c004000000310005450c33c04c0500c30000030c00000003cc010000003004070004040040000041c0700c0d010000001d04000c0f000000d010c0400f1400000c00000030010d000c000003000c404f40010000c3100000310003004c000040010f403001f00c0000000300000c0000040404c0030000dc00000000f300043c00040404300c0cc500000cc401c1c0400c4c17400c004000003d0c0c00cf004501330d300000c4c0cc0040c0010100000c0040000340c00c0f0040c101030001440707000104403000001130000c07c00000c147700000403000140c05c50d00001f0c14cc000d1cc0714400000000010c443c43c11007003f0003d43001c40300c0c000c00044000c0044001d100c03d040c0330040000040000300004011d0df00040003d440504000000000c0fc0000040c00300d0000000dd70140010c00000d0d030400c0000300000f000c003334030c700004c1000c040c0004004c0310c010f00304c00c04700340cc0000c5034003000fc300003f00000004004f003c0c3000300d3300000110004c0403c0000c340c47001f1dc30105004c0040d134c0730004030000413703000c33430100010040410d1000df440303d10000c4000501070010001d4003400400114c0401cc4003400441003040c1001104001730007c403000000c000400d0000000370f30000c4005034d0703000d0c0007030c4303304004003000000d0700cc0000000054304c3101030300000c00c003c007100003004cc04c011040050c04cc0f001010c000c3031303c300000073430114400cc300c3700d0f000000003003d3010f04cfc3303f00440000310000000010c3000f0300110000c00c300304100300300033000430070003c00c0303403300f0000030c4000c4000010f0000000300c0c307000000030103f0c70c000004c73004c411030000000000c0000c040500011c04c031c000300505000dc40c1000000303030000411d000303030000c00307c4c01405c400000044c4000404040d30000001000f0c030003000d10c140010c0d03030000fc010000000c400000000c01cfcc00000003010d000000c003c00400000cc003cc03000040001313700d031040450c0100010d100c0d00000000100000c500cc000c030000f0000c070440070000000d03c4044004100c00004d03130007c40c30031430001000100c00001004004004010334000d430c000000004c0c00000df31c530f4c40100000c400303000010d00053004000104001c0c000c1004101300004100cf0f300701000c000c4003330004c100003043c0000f310003000;
rom_uints[72] = 8192'hc4004040040000301004010c1030410470010040000c000c00000000000000c000040c70000100c0000000300c4033c0104104c000404171300000003f00c0007003c03410c00000c00040003c00d0004040000c4c0c14001074000c00101500001001c11030400f340011340330fc100000004000000000c04c00030070003003330000c0000070c000000010000100403000000000c131300c000040c0004100d000003040000030400000030c1010003000700030400010c400004cc000000001000001001000747010c000100030c0000000c0d00c000000004011c0c0030014000013030100300000033035c000c0103073000c0000000000300000104010030030f00f300011c00011403000003000000040100000000000003000004000d000001030c0c0700000030001000300c40000300c00000000403040030100d000000500100000000130c4c0f040c0000100c0300010c0003050040c40004000003000001030c0401111344130030070004310010000000000030000014410f01c03701000003030400004ff04c0410f0000000000c300103c00100030004047c400004004000130300000100030c00000c0005000c44000000010c00f01000000300010001000004c0400000000004000c0011030c17c0000007000000040111000003003000d00c10c01c00c000040c00070514000043d0c0c10004304c5100000001c10000030cc100001d4001010d000003030c004000010004340c00000007040010030c300110000300000001030c7000000c113000370f330404001034000000110007043000c0300c0430000400c003cc0c0c0c03330303000007000004040d3000000c0c0000d1171c00c0010003040c0c00300434000c0400104c03c00c0035440d0304000d3c0d000003c3414014010000000c04014053040003314c000100440004040000000c0004cc00cc0044030000000700000c0000030000030c01000300040040000405050144010100f710333001000000c0c00030c0000f300100000340000000400001100c004030030c000000010000000c0c300000000c00050007001104000fc3040400f10011003700c3000c0000000031010c0030000000000000301c3400c100010c00000000040000030001004c0047000004000130000cc0004d00000003050000000000300030ccf044cd000300040c0000100000000401441100000cd0c00000040cc01004040c004030000001c0003300040c0c04003c00000004f0030740040540000d3403c00c733000030c000004000304040c01440c10000004100c0000043c0733300c070033c040000c000003000111000403040004000c0040010000000000000040030031004dc31540010500310000c0000507030000040cc0000c04000000030c0000740003000000000;
rom_uints[73] = 8192'hcd31c0cd10300c0d013000c130010c1cf000fd003300000000003000014013c0cd0300fc30100040c0f0c010c007cc0031001043c000c0f35f0003001000000170c01c400c000000300030c01000f0c0030004450403c35141330000100d417001fcf0c3310130000103c10000f00d03000043c00c30033000010c11300000c4df0c34d0000001304030c001330c00f340000000000071004000004105130c1043c000035034d04c0c003003c000ff010001010001000500300004cc300100c703000000c003403011050000000033dc300d1333030c0c4fc31000000cd0003cc0d007000300100000003757001440333303771000100c010000730cf0000000c0003003d41003001c51d30001f0cc0f0d3033000c300c10140c01000050c0401510300cf0303340404100304300c000703030400001300103f1100033003ccc00c01100c0c1000f400105000001004100401c400c0c00333c001000003000cd30d05000dc077c50000c0043401c00000003cc001410d0000030d100704d00030400003c000010440700300f50c0c00cf001013000001c01d0110103c003403c0451000d30431c004c0030f010d004c0c0c00f30c11d340300341000004403f0c40430c43c00043300030000010100030c10c04000c300404030c00f0c5071f0000000300d001000cf31d034044c4141cc3c003401f00003d03c000f4c00010304c010c3f4cc10000001300dd3701030ccc05d0c40010cc0403333c010130040104070000cc3000fc010d30d000030000dcc1000ff74100003001010d00d000004000fc04114000003c17001c400c31003cd33000050c30c00c000c410411c03007000100000310000c00510c1141300314300dd0cfc1000c40310004000000003000044310100cf000014c0c301d007d10f0000f00305c0000d0305c04c007033c00410030030003cff100040400c001c05d000000005c10001cd4000000010fc0040110000034101000001000100c03004c3c003003c0c30014030c0303cc00000000300010c4000100410440044404300147cf03c4000c030c0c00c0440014010c04f0c0c4f11100f0101004030cc1000000000040c3004c4000d0001110000c0c00313100014c0130050307303030cfc0703c7c3000010103c70444040c0310dc0400403c0010071000000403000c04003030cc000000000300c00001c304003570c0f10007c10000f035001c030cd3c01104010c00dc0100f0401014007f30c00110004c010414c0c104d30000000c144c0000300001c001000004c00c130c0c334c00011001000044d00300300043c01c4d000000000004000c00370400c31fd0000103c0033c00cf0d00003fc0c0300010000c3000000034c1c01030f3000010c40304d41100c10c00010700700c10400444430077c00500c00010c0;
rom_uints[74] = 8192'h35101000d0c0344010c0130c11000440c0340004304dc03000c0c400cc001c10000030c3c037400000100070f0000cc4cc000034001f40cc040003107d0000303000c003cc3300f00300c0f07cc00350300c005113c00100140d047cc0d004d1305fd4d00000fc000010c0404050cc004c0010f30010034000c030300cd0f100003c000504000010003410400000c730000000c4000000dc01c000143c50100403c034c050c0433410c1c00000c004000c4cccc000103040300400013c040c130334c00c0400c010034c0007c0c0034c007400000035003000043040c4350cd00334000030300400000c010c10f030c000000350017010c300030c000c00001000003043400030c4107004c0301000300c04340c0ccc1000f0c000300410031400311300040cc1107001310f30300010033330fc4d0350000cd03000fc01404000000314d0040100d040040100000071333c000010300500c47414c3c000f00000440310700300f000c0340dc00003d4005000d0040cc03000ccc0100c301000d300133074004070f01000c0fcc00c45cc0030c01c00013030f30001003cc0104cd344000c3040c0004cc700c5300d0010000c0cf0144cc0131c1c011031177c30400004c10000f300d00000dc00cc0404330000007000d0c110000cf01cc05cc474010000034004c00cd03c01cc40fc1c30ccf300c00007f0c030c1300c54f034001500cc04000c730c000014c5043100340400c000501000fcd704f30c03401000f0105c3040000045f10000000010400404000cc300004040530cf00000140f507400cf0440c00000cc10300c01143ccc000000300000303000d050011000100c0c10f0ccfc000014c030050010c033f40070c00031004010340000000433000035dc100000cc4c103400143304305d4404cc1300c4100005c00040cc07c0fc0d3010340c0030d00c4440433000504003f01010300c0073300fc0300c0000d0c000300400000003cc04000000f0000000c0000000f007d14c00c03000ccc00000003c107310030004005c100404000c04cc370030000000c0d0000300f03cfc40c0100f03404700040010000c000c00043435001cfc0031507104300c3430cc3d000c5010004050531000c0103405cc30003000440030c0dc00c074000000cc00f040c040015000c0c304c070c000000cc0000034000150000000000010300f045410cc030005040c00704500c4c100c010440074040070540070000444cc400030301c00d01c00fc001044000030f040c0100c5045000040417044000004c0fc3000c00447c01c10c00000c0340000c0000031005013c0cc04000000333c400c307f30000cc000000000c474000c3000cc010c40001100d400035404f0300000f0ccd30cc0dc00c1000f1000fc0ccc0034100070fc30301404c300000000;
rom_uints[75] = 8192'h30300000f0c100130000c00001014007010000040000010c0000c000704043033000000003d0000040000300c0000340c30500c000d0f100000000400003040030000003c000000000000000130000100070000000403301000001000033110000c03030100001000040000000040cfc4040104010d040001c00003c00f1000033030100014300000004000000304100100000000000000003c00430d3c711d00001400000001c01000001000c0000c00000c0c000000300000000030c010c044000c030c0003100010d00310030000300300000003c0110000000c010c00000300000000300000000740003f070003400001003500d1000000000300000003000004030300c300110f0c000305000c0cc511c0000014004c350010050030010001f000000400000000030004c0040001d000000c0c0340040040c0cc0f00c030000000004c03000031000004000000310003010010304101004c405004000000005000041300c41031000000100403000d0c300004000000030f000000c000000310000c011100c0030000000001000070000000000c0000c0040440000000000745c0030000030700c00d3c0004070c01000000011030000044000c033071000000c0050500050300100d03c0001000f0300000130400c001000000050c00300c000370000333000400110cc400000c0000040003c003000000300100040c0000030c1c040c01300003c0000f00050100000001d040100c0000501000000c3c430000c10dc00130000c000f1000030c03d100000010300c0c00000110031c4c0dcd000000040300c03701c3070000000000030000000300c0c00000000003001300033000c000030030d10f00043303f010c5c003c0c30030000031c0300f4000410004004c00cc3c0040101300300700000433030c000000001000303f4000010f01000f410431d00c0100000303000c0300001010400001033c010c004004030c10000003000003000001400300300041f40c00000300000330c5c00300cc300301030005000000100104100010030103040000034003010c030c0307000404000004cf00001340010f40c40100c4c001030044000c00047000004300030540700000003013cc0c400c000000010000010000000003030000000c013300f004400003000000300000010c10000000003f03000cd00cc10000100004c000000c0403030000010043000001400f0000000c0c0d0010000d007033003c000005d000000000070c0c3313000000101c300150001f000c300000cc00003307070c0001300317400c000300000100000100000f430300007330c010c00007010003000000033d030cc0000c0f000c30000000001c000d403f330c030000005410f0000000000031000101d000050004000730001040050fc0040c0d074c00f0000;
rom_uints[76] = 8192'hc30c400003000c000c03003c1140d3c0c00303000000cc0033304530c000003030304000000f0010037c000040300f03dc0303f0440c100301c00c13000000030403003c000c00000c0003001000133011000013c0530c40000d0c1003c10100c045c300430000400300c3014000001440010001007400040051330f40c01000d0c3133000100071d0c003040000000000430000004030130f003010014c050001033c00000000100010000000f0030303003350000003c0c0100000c3100f13410d000c13000cc4010100401c001140d00c001103d313000c3d0c31cc000034000300010050030003c300d0000c0010d3100010000000000c0d0100000100000014130030070103011000100c0000005000004001001000044400c10c03000c003003001103000111000c0d00003000000000c00000130001100033c1c300304404010003f0c00010333330f003300000041301030340110c0030000c013003003374003400000040d0010050100100000010001000000c01cfc001fc0d00001313d3011c0100013100000300000010110000df410000004003d000043010c0000c00c040044c0103f11010004001300c000500f043d3d004000c004101003430000003100300c0004000000700000030c0cc300104030010000000040101c030c00f0100131c13c0c30c00000c00c05c100310c0400000030300401040cd0d03004003001010310044100003c00c1003f0510300040330541110013d30c011000f0f1073045d0c0031c00413c0040000c31c00001c3c01530c00c004000043c10301c00030f30001d00073030100c000cc01000401300000030003310103301c0d000443000003300c70d4305000043c0cc0410d13041430010500100300000000000c0000030401401000c030f0034300000c00501000000300001030c0000110000d300010334c4c03304030013133000c434041304c0011331000c013c30f0053000000c0004f04070000000001005103c0115003073c00c31043041000300010400103000000400141403300010700001003001c0010001000300010010c00000c34010005c1000030000301400004c000010001000000001000000304c1f033003c000400000310010300030000d00000005303000040004c41000c000c00314003003401003c0d0033003030043000c3000700000d000001033450c0030c100103304014030c100413000003000000c001000000014f000ccc0000030100000f030040004f1c1000000040074c00005f5031010000303c41100300c03000c00c0d33700c10000000001c0000000000c0c0000100113001000330000c0d00cf45300f04010001040010000001000c000330710f4140c01010354410c30000c0000f3100d04300000400f0000001000040010114cc0050004030010400;
rom_uints[77] = 8192'hc00100004c00400000c0000000010000004030000000000000c03000d0000c74004070c000000000104300c0c000c0403000000cc400c003cc0040030000c000414000c4cf0c00d00000c0f0c0000003c011400cc3c050000300340cccc04d0300c100c04000c3c040d0c001d0041007010d401c4010030000d0c140cc0110c013c00040000c007010000033000400c03000000000c0500043c040000000004003c040c04000400d040c00c0704000c000040040000c014030000000c0c003010c001000c1000013c04311d001c303c000001d000010c0400141701500440000c0100000c30c000004010040003c00c000300000c3c00000001c0003000000000dc003c700c300054000c001c00000000440d0cc00300cc1c3c0441c703141004040000001400f004d0000cc13430c0c7000000343d44003000040000300015045c0f4300007000030000000000300410cc0014000c00001110cc0d4f440004010c000400700000d0c4c4c430000f4000c40c000c050300044c004001c00c0007400100cf30c0030000011c0001341c3100105000300040000001c00c500003001f010c050c300010000044cc04014400cf0f000f34000c0000000004000dc3303d000c040c3000c0040410143000000c00040c0fcc30173000000000040300000c07cc000004000c00141c000c000000c0040c100c3014c0300cc10ff4100c50c00003307007000c4f303040001c00000d3c037c7d013000000c0cc7100c03031700003f30001000001010043100300001c03000000c0000000c0000000c300404301000300300000c0c070c040440110004000d0000030410301004d10000170000140c3400000010001000040c0c0c1cc00400000400400c003304000000000c1400000c3001730330004340c1001000050030000300f0000000cc10cd0000c0c0000c010c0010f00000100c141330d003344c340c0004000300c11c100004000c00000000303c01000000000d00103000cc05000c3d04c301010000cc0004c00c0000d001040004300040100400dc1000011040000401000030030c0d10031000000147011010440c000000300c004001000040000030000f00000cc0cc0505000c300c100000004033cf3c00000c0007f0c30fd0400c03000003c40000000034000004041c040d03d0001400c0c1100000400070040500000d0030c033030004c001040001cd0040c0003c000003000414c00000400400c3040000c700730330100000000003400004fc701100071300140404143c007030440000400d0703c000000400000000000c440c0000c00004051c7003000030000000010cc00004400c0033005c3000001c00c45c00000f00300001131000000c0004000001004400000000000c000c7cf0400000310c000000000500000c0cc40030140c501;
rom_uints[78] = 8192'hc0400045f4c0004c44000c004000000c000000100fc1f040000dc0040c1000000030040003000c004000000000434041c070c0c03034f40cc00c00441000000500070700000404c0000701c43000004c4cd4c0000000cc0000c0000050c00000c0103c0000c07400f003d0c004000000000c5014030030000c000404041c4000c3700000c030000000000cdc400c004c41700c000033c0cc000000004cf0041c03ccc00c030030d004400c1300300140c073c0d000000000dc0000c00000030041000004000000c01cc30d4c00300000303000c00cd00c0170d00c0dc770000f301000fc30c01004003400f4c0c0400c030c004c7c40070000000fc00010001d730100400cccc11000703010c40331c00000cd30000000c00030007c0434000000043001100cc0c4cc003000401003cc0c0001c0000000ccc0c0d0c47c00043004c400004000c00cf00040010000003000300c0344c000cd10dc30040300300030300c30cc3c005f015510c01005d00000c004c000000100000000c00c14044f000c33c105c00c303c0000fc100055cc00004000740000401404f40c000c0404d0fc1c000dc30004000030001c10cc000c00345000c43c033000c00c03c0fc0004d4c03c000034c00030cccc3000c0c040000011501c704000f0cc0c0c3c00c110ccc010044000c0010d740c0000103440c0343c440c1070c430000c0010003dd0c003c00000c00300313014cc00300c0300c000c0c4000040c40c0000c00ddc0304000000100330000440c40000f001071c00004c00031c300003c000000004c40dc0f000001000c470304033c04c0100000c000d1000ccd030d0cc3007100040c00010c3c01c00d000404000003c5010504f10044400000310003c030000334c1c000034f001030000033cc147304000fc30c47c7c00000c0300030413f7cc0c000401c00010414c0000500003070011c100040c300030100474c00c4033000100300c000000007c34c000c41040c434401340c10cf7c000000cc0035040300000f0fc03040040f0d000d0c5044c000010c010040000130413000410c0000000c04c003030c030100000400340104001c41c0003c01000003010f43001001c00400000d4100000400401c043000100030000c000400c1c043005fd00c0d00003c000000004c0c00300c00c01000c000cc14cdc043010c040cc4004000c30c03100c0c030c000044044d1d0d000000c440311c10030400d0000404cccc0000cc03010c03c000c0300400000000004414104c000fc14c00000f3cc0c1f00444440000040000c001c400004c40100004003000700300c103000dd000300400000100050000d50c0000c0cc400001000000c000400c40000003040701000500040000c30cc0000cc70d1c40c10040c100c30000733c013c0c40030003040000cc;
rom_uints[79] = 8192'h101000c35000031000000f0c000cdc00400300c000007000fd04c3c3c43110003701c00070000300040004717104c03f0413c000400c00c0700013c010c330000040400300407000030c1000cc05000003010c01011103d0000000000477d00310f100c00c00000c01704004000000404001c007c0c0000000c0000c50000300407030000c03c0000000110003330003c0c00000414340000400004000c04011300000000c04034100c0c1003004300440d0400000c070c0c30003400000400c040c0c001c3010000000004130440c03f033000000430100c030543100000045000045017dcc00000000441c40c0004003300001f00c33000003c0c00000504040010103c0000c003000433010000001050c000f0330c0c13004d540400300013040010735014043c1030005014410c3c00004c703d0000010c030050c304d0040000010d0c30340000003c0313005c01000034d7700f17404111d3301000001001000031040034cc0375f000100c0050003030c31710c300d14004000000d03cc03014073030041500040c01004440000300000050100c34003c00010030c434fc10041010000330000440000010040030c0105114013c003013404f1c4cd003040cf00f1003001400000c00c03000000110000c33000000500050000c410cc40f0000000c0301ccc3340c300034034d0f0400c00f01c0040005330ccc101011400000f10000000430c1fc0000df00010c007ccc14c07000041ff000133d00cd13000c70014000035404fc0004fd0003d10000070300313104005004040d33040f004cc01040030430400030014d3000c0030400c0c0005401037000cc1011c000007000001000cc30100c00c711000f00c0001014004400000000000c15000c13c4f01c040000004c0c1dcc140005400103f1f0000c000c0401c0100104001035c401c13c4c4000001c1c100000c310000d0031013c000007040330003017003407000000003000034001003c0d00f30f0c4c0300303c00000000c030d31300c0330500000c100fc0000005c007345003f000070000c1000410030c100000010300000100f0c0000000400c0c3fc0c0001004c7000040c000c004043030100300001cc7f33df00440fc000400104403fc0343d00c3000000040cf0070044d00c300301f0001004004000c001100403cdd0d00100000143f3d000000000d1400300500010c07303d0030000000040104003430001cc00c4100100d3c0c0f1c0100570000f300000034c00c400004034c0f5100cc13303c00000c031040d104d040c4c700d70cc70c100000300003c0170003d000c0030044c70001003c0c00c00cc000000d4c00d3440401000400000cf0044004004d004c04ccc05d04143004cc0300c043001030c0001c000c4c100003000c400000040000cc00000401;
rom_uints[80] = 8192'h43000c0103c004c000000400044c0130000fc00005cc000007034003703700dc03000f0300003030001c0304040304140004c00c404f0400004dc13d0c0001000c330c03400c3400001cfc00003f04310001c0000400040cc04000c0cc04c430350d030c043104445f0030030701410f0c33f00c0407c1040c300c40043150c01c34053c013f4400003cc400c7f4043c000000000f0c0f0700001c03f00c000f4000000dcc0000010004043104040033700d000d400f01030cf444000300300c000c0000c50413004013000400c004000c03c30c0000300cc030301000000c030504044dc000000004cf040f0401c4005400d4040c000000c00401000400c30c0004000400140001340c0c00310043ff4404400100037c03003cf004010703f00000400000000f0c010f0034f13f011000040f440c0c000130043f3cf3c0010104000003000003c00c040301130c0001010004cc0cc0df00474c0cc00c0510340440041cc50400130dcc00f00c0f0500303c00400005c0000c400500030ccc00000310300cc0c000100c3c30030341001c05000c0f0c05001c03000001043c0f0050003c0c01003041300504fc047000114c014fcc010c0030f5000140c01000000c34001f0d0004000010c00114c10c00034103140100003c00000004010000013170010c004cc50100044400043c400000030c010000013c00040d40010400043534030c00000c000700040c00c3c00f4154010300100045c50070cc05003000400c070d0c003cc4030030000400051c0000c000300c0c40040f00010c040cc4c00003040130f000ff03003040c47104c0010000053c0f0035340040c314040c1c0314003040300000000c0004011015f300010d1c0d003004040c700c1c4c000441000030c0d04c53040400143ff314004000cc3c004010000d00040c0140404c0c51000130570f00004000cf0000c444070030110401000c100113000c000100000000040c7000000010010c400fc0040400000435044034030031300000c0c100c0400c00c500f300071004010c0c340003400000000c3070c040c1003000c00c0c000c300001100c0300000c50443404f00100c00f0000003001000400010030001c040f000431000000440cc1330403004cc00000030c00c0030c400cdc054000043c00044000050450040c0f01c3000cc044130d04000040400cc000030c143c00130100030cc3003113315cc03c0f0cc4c0130c00300034c371f0000c010c0000000114004c40000401040c403343003000030330003f1400400c013d0313040d0100010001d00c0f0000100000ff003c340c00040000540400000031f30f0410000c0c07004d00030000040400001d003c10400c3d0c44c004401c000401cc101400003fc00f330431340c0044000004400505000040030050;
rom_uints[81] = 8192'h7047300000000f00143c340cd40000031310040c0040070000400d004f113f0003000d4c33cf000030000000030c1000331c03050c0100c10400c4004000100d3000100c000030740400300f0000fc0000400d750f01400d0300030c0c00004100c100070130100100300d303c170107d00000f000310003110d000401330f007c0f0000010004c3000300040100dc10100dc000003c0700450007110100c400c1110503300000043c0000000c04000c000cf00300000c070c0000300c0dc03cc40430000c00d003cc0433dc0000c03f04000c3f00001c000c500d0401070000c00c00050304c0c000030135003700000435100f5cc0010000300000030001c03110000c070cc400cc00303100010c0007010cc500100c004c0c10140033031000400d00c4003033310d303030c03c3110000c04431c03303400451000403c70100fc40000307130050110f103040f00300030f0113d4d301330313001373400000100001301340dcc00004401300000000333000c00003400300000001000c014cfc40007010004334004300c30c00c10000003010071003030300c0c01140000fc3f01303300000000d0030c030100340c0400c055030000043431000000101f03000c0c0c00c001403d030330d01001000f10c30c0c0340030000000001000c0144f40000370c00c310110fc3000dfc00000cdc1114000c003c0000411441f1007310c0fd3d30f00d07003343cd0100f03c0010000d000500d003c0000100300400000000000c000031000d03050000000400001c0d400300fc03c100000c0007000c000d000004000c0d0c0300001300100c0504010000440f0c3f400f3f0414400c00030000000010430c05000cf310340341fc400cf0040f00010c010c01014030f0c0340d013c0d10030403033133d400c3300d33000c053300f000003400000030031003010400c010cc00c30c000000d03131c0fc0030400c100c0c1c00013000003503030001000030003703f00c40040000cf71340130cc40013300000d01353c0c143431c0c00400133404110d03003c140000004c00f30c0d0071c003440301040c000100030001300c03d0000c030cc0014cc0010c0dc0000cf4753000340140003d1443c400013c0003350104003f000c0000c3070c000f00dc0001cc003c410c0307c3000001c070000d00010401004100d711000f343404000c0f37104d000000400c0c41300040c7041131300c0f00c40c003101030dcc000c31010400000000310000001d0c3f0ccd0c1000300100000050007c1c03000d0000010110c30001000001c0300130003c0404710004c30411c000000404000310043d001f303400030001f30c00300303100000000071300c04c4130100300300c1000334000d0d50310001000003400c1000000003f00f0d00cd00000100;
rom_uints[82] = 8192'hd0d0100d10001000100001c13000c00003c0cd07000103070330c040000000d3cc1030000070ccc0100301f0f0f0010ccc0437c1300011f00000400003001000301000101000f0500101404100300301300043c03131d040c7c00040c03041f30030303300400300f07cc0d0000400f0c433003000f00d030110c7fd41c100005430c000034000000dc040f0300000f000001001c031000d0030110130400001c4c00011000cc0f0401c30403300f0100030310000340005d0000c00055030f0000c4070f0c0001500114c000443f4000070403440100044005050010000000050d0000004d000c00cc401010f30c04000004031004300040000010410030c00c0140000000c0014001001010c0000d5f503c0003010070300c030303100300013000010003c7340400c00f0c40010c0401030000400dc300340001c0403000100000001d000f0f01300100157004c04411140331005000100c0d0000340f04c10030311415c100c33c11104f7400000c30000c111c030030000c071c0104000d010303034c000c074004050c00100c0300c404011c0000000c000041404c04c70c0013000f00400c0004013cc0c0540400100c0c003c000003403100303c033103004000000000310c001000dc103c030c041c000000c00c51373c0400003510cc0c40300d040407300000057c00d104c700c7010d00040c4c040d0140040c0f000c010c03000001c4c0c013070000c703410004c004c04000001f40100d4377c400004005c00010040c0c400c4d001c1133030043cc000c0040000c0450043100cc0c4c04030f100713300c4f01cc4d5f04000001003d0004330c11003050140313111c004000330314c00c0000cc37400d10004303f01c030040c000001103040330130f0010000100004000000000000003300f1c000400441c0f40330100040000444d14000d4c0004000c000000404004000300004c03000c0c01000c0000000c0703300c0cc003000005cc030c350100000c334c004100000000000000030403c0000003300001300351135f0030000004410010030070000cc00c0c104c00030403001cc00007051c10cc0053d003030305004c0c030d00413400000035000f03400c0f70f3000c00c30c0c0013000c4f300c10030307003013040300c00d030001030000c04503040303441c34030004000404003010010d000000013000050000040004030c00030c070c0f051431403700110303000c3f0405c3410cc003030000410704000000457044004f0000c4d1400c1403c0400c037c101100001d00000000301100130004000110000000304000001300030c0000c51f001f70d404003030040f37100710000030000314043000c503531d041040300f040c0004000c3040d13410000d00c44c00000c4d00000c0440000040;
rom_uints[83] = 8192'hc000000105c100c003c0444f0043000f4300431304f00703c00c10000300010003330c03330c033fc100440403f000c0001073c000030001c00103070d00037001440011c303000000140300000000000000c01c3100010d310003000f100000013001c1d0070000003000330403001435005413100003000400140040d3300103000000c0000100030c010004c0000c01000000c0d000d300c0c034010d303011350030000037340303f04000010000f33c0100000000300c000710000000c00c003c40003c50007000c10104403000300c0000111330031c7000f35100000000000403350301033000d40030c304c7dfc000c00f004c330004c03000004fd3400004100370c413103c003043005c30351000c01cc003103000100030403400340700cc03c315003000f330000000314c0031040fc00030010330000c100440c0004000010040000344dfc1330c0035330050003000001000301c0370074000c0c01c000cf0c4f01d3041051010c033130f000014303c0c440300740530100c000000c044003f34000000111004737000473700000c001f00000fc403000040050c000000053c0000000c030101000c3040005cd010dc0004c400004030111000000c30000430170404000c003030340700c0001013c1c030104041000f4c4017cc003010c0000c0430001c0704340f00100300000000530700d0f34000cd0000011343030f0050f000c100140ff0c0003c013030d0001300314c44000f4004003030c40c00300000040340050001001c0c00000040c0f0cc0700500000cd0003700353040400001700d00000000004001000c01d40000030143430311c0001013000070434f5cc0000cf0c33141004033313cf030d300fc403030c000d0c003444440000014430300f4001000000300c50370303033d040c301100000330017730c41c4113f043d001003030013100000c0d0300c0cf10c4f4c00333000c003c30000000043033400c000003000d00431c0f3c00c000c0003700c01c31f14c00000cdc1003150003000104443f0d000030070c0330c00c1040300c040700f10030f0011000c03030101c03c7030c014c01f440050300040003030407140f01140040040010310010073c1c0000000070cc03300000333c1010034c00300410054000334d000c050400c101004101030c0d00f10005300130c305300300030540030100000c0533107400d333f0000040430c4001c300000000440300c0303dc434003000f00030d730333070c003003100010d0143007c00130d300704300004000007101130130c013413000030010c0044070000000004340000c533303000c11143d0000400440151100003350030000343c030300013c1f0010d13100c1000703510040400cd03000c173400cf0303000030003040300003c0100500;
rom_uints[84] = 8192'h10030000001331003700f104c4400cd5c00010001c0000000003000c031f3c0100303000fc35000c4c1000340001150c33000074c0f00c0140000030003000000050103c30700040000000c0300040040030cf40fc000040c00f0030003030000c003c340003000030cc0130c100005040013000000f33c0000401000100000050cc0d1441430103400f000c00040040000130000004110003c0050000143c00340010004000400fc3c000000040003c50cc000c00c040c030000010400030040c7000303000c10003031c004c30f00000003000000df0c031404430001cc040040100101033c00000400c000c04000000c0430000010030c03000000c0000c33044040004104000041003000000c1300c501004300cc0000001004cc13c00030014c000400000f4000400000c053003300100300c0d0c0000300001300c0000cc0c30000000000033001c50010c4410d0040003c0003c3050004710f0040000450c000c310700001c0c3001f010c0f00c01c040001410103114133cf4001d000f3c04000000300004f00304033000010000010000001004413400030110000000704100f00c1000003cf43017013d100000300ccc13c00010043f430050f030c073035c13c00501000c300c030000003c300c0034fd3130100c01000c0d10cf003011013000403c00341034000f04c300301c0c00c000c4c0000c00003010df70400cc003100004000033113c10c044044030000c30100000000034dc0300040c100300c33c100c00101004c0040044400c3400003c00500033c004000031030f1070300004503033cfc0300013c00000450000004400005044000c70100c3cc0040000043000400001410d00001000300033014000140010040001010c000314400504043000dc0330130001301570040fd1d0f5c010c30000f000543033001400300003c37c1000703470040300c300fc0030c07000d0100037000c0c00d00104400003000000c0c1000000300000cc000d50cc000400000f003c040040c000000301003000301004304303d000110000f0c0303000000000300033f4d300000440000030403dcc140100000000c00c0374100330100010401f0004004101011100c40d000003503fc4c00c04031000407c04700fd0000330007c0030500033700050000011c00444cf00403d0000007000004017031400ff0000004130000400101331040000340c4000040000043c00400003300c01454300370000c03f33010c0301d0030000000010403034003c30001c304110000300d54400c0000ccc05d007c0c0334c000c0050c0c00000041030000000c0010c00040000444c0f00cc117c05c0c033030401000300040330003c1000010034c000100010003300000030000001000370dcfc000310c00144001d000000504701c010fc00004400;
rom_uints[85] = 8192'hcc10000c5f000000000c00cc00000000010030c00cd04c000ccd40000114000c0c0010100cf000400400004070c0000c003410c40cc00133000f30031400440f0000cc0000d00000c00030004000340000dcccd0f070f0004130c0000013001404c003000c000034000d00000000c00404000000f411000000000010c1004003010004040c030000000030000100c4c004c100400041000c100d0003030c45000c03c30000003340010000001c0000100d000000003004c00040040d030130c031700c000c0c300f00c00cc0c0c0000000000c0c030000000540101415000000ccc0000c4f4c400f0c000c070cc10000000334004030000c0040003000000c0cd000400404c0f005300740030c00030404c4c0010c010c0304300f00f000400001c100007c000cc0c0003000c40c30130f0c00c0d30000000000000c0010c00070000101001010c131c0c0f1000c3004cc0f0c3c0d011f0030155140003131000c01000c0143c000000040c0030001000000000043f030033000c000f001003c033c300c40003000c00000040004310030000001000010400100010f001070003004010040440000430c0000430f440033001f304110000c00003000001535110304f004300403f000d000010403004000000c0040c04000400000000c3c1300010c0cc00c0400700000040c04000300300c1c03030304000c04001040100c104cc00f103531540000c030c0000070304140000c000cc07c43003300000d00000d033000000040c004001000001005400fc4100f0c03c40011000004010004003003c000143000400f11000c04310000000000030f7c0000c00400c4000d400040000500000000dc00005c0000053030fc4cc441510c00040c040303000d0000071000040d000c00000c00d003005004003000010d03c470007100044000003c0c3000f0004f00045c040c34000000004100c071000003f4000cfc40cc0c010c0000f00000000c0c0001000000300000003d000c00000d0c000c00013c00c03100003cccccc00000014c37c303000000000c01400c40400fc000000500010000040030c301300003000f0530000c40000000700400030100c030000000c004c04cd004000f0c03013044000000003000cc0000104040000130000000000400c00000c40c00000000000c040430010000c00c0d1c05c000c03300000000cd00400004030c0110000d00130000100d001c00000c0010010c0305000150401cc030c4004301c000300000000c0000dcc0c0045004004504400010c0d0000004040d0c140103000030c000c000c1003011000c0c34c1d00304300003400030030c00403340110c740c0000c3030030c000100000030003c4051c000341000c00d1303000000f0c001000000c040004504000110000c004000000fc0c3c300000000;
rom_uints[86] = 8192'h1c0040000c00000000004011000000c01430010000ccc0003c04303004000003c01000c0470000000c00040303003c004c40c50001001c4000c103c010000000000500000031c00000c00130000c4400340c0c7c3041103c004440000000c000710010d4000c00d0300300300c0f5d544c003340170041001c00470004c3303cc300000000001000000040fc00ccc1001c1c000000c000370c000c1c40374401c0340011000c00040004010400c13303040c0000c00300c0c30447010c10000cc0000c100003c00001000c030c4c7034030005030f3f0ccfc0c44034ccf300c0000c00c3f00030310c30f0303c10000100004d070c0c00300000030000000000c0df0330300400033c0c14010000000035000c040cc3c01d400031000000000043340030f70c1000100034d4143c040001100010011000f000040035043f04430000c4401330000c010400130c0000300000440003100405c4d4333c413000003040c000c000f00300c0310c0c330300130301c00030c43cc43f000000001c001c7cc7f70004030030000103000040c0000c004000040000c0c110000c300101113300000144300005c5010707000030000310cd00000c30004c0400c000040c0100040c000010000010001000000030f30100400cc00000010404003c0411c0c00001000001070d3c3c1140340c017c00f0044c01001130000000c0c40c71c00040000033140c03000001cc00000003140001070c0f0cc1050c0c0300374c0004d40307c10000044004000700001c100c0000000003400104000003400c000c0330030400d0000000000430dc04000000400300100000343000cc4000107300043400f004c30c0f00cf030000430000cfcc0000030c0c0031040004774000c000c3314c000000040403400000c30030434d3400701c4000c00c000c00c0d4c0170d3d004d0000c0001440c0c0410dc3300050001c300343000074c0000041004c000000000040100d00040c03f0003c3c03c0003d00403040f0000f01c13c30007c3cf1043c10f0073040350000010c0c300000003000410040000700030c0c40100004c010130010c30c0ccc04004000c3001040c300340004040040004400c1005c0000c0500000f030003000c0000010f0001c0004130000100c0005001010f30c0c7fd0500000314400003c1000000134000000c040fc0000140050010000040531000000000400030030000040c0d14105000c00014000043000400c4000d30004004c0c0000c00f0000150000dccfcc0c0403004400100c4734004000300004313040cf003c0000f00c000400f010400300510400c01000500cc0003130cc04c00cd4070000c000001000000c0000000010004000003d0c5000c0c010c3c04c0000c0c000cc00003000f700c1000c400004c0c00000040c00040000;
rom_uints[87] = 8192'h34c0c10010000c13c04000400500311ccc300340003030004150c140c134403040000040000000c0407000130c0000cc4c03000703c0f000000031355000c030c00000104000000301000003000010c03044533040f00f073000c4c00030c704c03070330c0040100001c40cd00c00430cc00c1000004000400001133001c040c1c0f0c430004000c040000070c010404000000000000044c3000000c0003103f0f000c00c30c00000c4004004c0000000d0c01000010004400000c0cc0000c050c400000000000000c0013f4000054000c0400c0c3400c1000000000510c00c305740000030f00040d400f33cc0c44040c000000030c1000000c00040000041f3c4f043c00010dc04d004f404004003c0c10cf0004300c1400000410331100300c00000051000c3c01400c00043ccc010000000107c0000047c40031000300c044000540000c000f030103f0043403010001500f0c000033000c711c4c0c043c00040000410cc100000100cc000c007300000f0301000301c430031cc300c01400010d004f010c0c334c003c400d0f1f0001000003010c0530343f14000f030430f30300043c01fc00c00001053000000000040000030400c000c000000c1000c4c407010001000c000c0c0030000004cf000103400d53c000030c000c1047c00c04070001040310003c540404000f015f00003c0040000040040000000c100f030300000c500300000f100c030c4f0330000001031fc0001c03430100cc40030d430c00cd4c0cc00001000003000c01444f0c0c0004c501010d000050004400f75f0cc000003c0000403c000031010307000003003010000c05c4cc01c1000c130100000000040003000313c070000400100000034004000100000c40c000cf000c00030004000104d000070001300700040000504c000c00cc000c3cc000003dc0cd1c440dc00003400000000d010c1074000004000010000c0000c0c304c340000100000c000f00c000cc0c0014100053044040030c00003403310403d0003000000c0c0c10000c0c000c0cc0030c1c013f04c00000043c040000340d0100f3000400cc4c0d303000100c00cc140000030000000000000f001c030c0c004c000000000c040c40010005004c4c0f00000303000400000f0003000c0004130000000403040c0c0000cc1007000010000fc0000f00c4c000044000010014004000001c003d30030030501c3c0044c000400f004100405c0304001c30170d00d0c3fc010410000300f01000100f1c31c40300000c13000c100c0734003dc00fc000043f0d3007441d000400f00c0c00000c00040100000000000040000c03140400104c000100c0c300c0c004110c0c00c000000000100f0c05140300cd1041000004c0011c30000c0400000d01003310400054c0030c0c00c04000100000000;
rom_uints[88] = 8192'hc30000000100430003000c1dc303400f04044f010cc400c0044cc0c5c107003c000000007000000f0000005d000c04003013030000030000400004000000c30c0cc0c00c00000414000300300000430000040403c50fc400c40001cc0700004000f7c10c00000c040c000000000d000fc0000c4c0cc007000500033000c5040d43c04c000000c004c4c00000000c4c010c000d00000000c40103c400030cc7d0030c0000004c450000030103013f070c400540400040c04cc000000fddc000030340070c0007003c04030c40c0040dcc004d00000300c000c0030c000fc0000003c0000100110000000000753441450400070500400000c10405004000400ccc0c04010f0c07c000054c400000000004440c0104100fccc107000400003c40000700000c03000c000401030004000004c40304000f03000c050c000c00300c4c00c000cc03c0000000003cc0c4ccc00c410003c070000340004f0c4c030400c0c000031c4cc031000c0404c07c000f700003000101000000401f304c01000004340000010c0c0001404cc00507000041000000400000000c400500c000050700c140014004000300030000404100000040000ccc4030c4c3040101010c00000c000303010c00c3340c000c0c003140040000040150014004000000c3000c4c00cc0470000010040c010c0cc000000000c00040400c00030f003003004cc7000003000c00c00c000001c00c0c030c040000010005410c0ccd00030000c000440d00040700100000c00c000403cc000003c00003000303c03000c100000404000004c000c4011100000c000000000003000500000cc00c000c03f5030c0c0c000000000005ffc1010c00000003c050001000170c4c000400000100010043430c0c0cc30040000101000f0d0005c01cc1000f00c4000fc00000ccc0c401010340414cc00000404414004c03c043c0044c400040030d0103031001c304c0c0cc0cc005400000400004030c000000000c40c00c0f50040d00cc1370343134030cf5070000004c3347040000000c01c0c0014d400f040c00110040000cc134010040044f00040000044f100400000001410c040d04000100000400cfc00c0f0700400d0f7303c00c07040d0004c703070c0007070004000d54000007000440014000400004000fcc0cc000040d000301714c00000cccf10cc000cd00004000c30400050405c04c0000cc03c0304144000c040000030400030f400c0300000000440000c0040040c00c040000030f030000c30c00400330000f00030003f54c000101030c0000ccc00c0000400405c00000040000c0ccf30001400001000004010001010cc00d4f015cc004c00f0c0003f001000000400003000f00034004400c000003c34100c04400040000cc0d0044c100000c034cc03400000000030000000c000;
rom_uints[89] = 8192'h1000400f103300c3c00303c01000000c041043f30300403400c70043000000000d301c40340000340010005c40004410f334000c004000f0000000004c01000c403044103330004040004000400011011040030001c040403c315c0004c1000100000c410000c0100000000003110015400040700374004010c0001c00000003c0034cc0030c00340c5000001c0000d0000000000c001000001cc0301cd0040304051040001010473c0004000c0001d00300c000030c00103030000344c0303c0c030c00000cc100300010d033c31040004c103041001030005cc00040d010004010000010010000f4c00cc01c30c000147001004010c003000c00330000cc00000030000000c4350cd010330510c013014000c0c030403334000303400000300040000c00304f0004011f07703030401cdc00f303ccc400400050c07004c07500000030004000000cc0354f343004000000147730013c010c10103000d01000001300041004040055c00000000000c010001340c7000530133003033000040073f114313d330c000000300c400000f00001c0c100000c3030c014c0030007004440100d3c00100000400d001003000300000340d00000c3c0447040000ccc0d000001c43401100003000000c000d100000000000000f0000030041c40303cf4300300107c00cf000004c000003000001c00000010007c00c000000430c003300c00704000003000100c0004c050103011300700fc13c13004003111100000f0003033001040044000005103c00c10d0031000300000300c004050cd100303500310330434c401403000f03000c01000f00000000030000000400cc10030100540fc10403100044004c0c01c0001401030000100c4c00000003040000004000030100400013340404c3c30111ccc00004145d4f0c43001000c403101d430000c11000000f1010cc0d000000cc003000c10170100000000151033c0000430003000000000000000330c00c00031303c000400140c0400c0003033f070100031500004003040c00c0011c030300400c030350040f300c00003c0043004f04070300013d04030c0c350700030d00330400030c130010c30000001013000c44f031c10d00c0cc4000c0403004000c03040c07004003010005100c0c00040c0403400c001003000d010000040000c04400340000100c0001000010003c00000c0c0031000100440300d300cc000443003000000000010f00000000430010000c004305100c400100500c33400300030c00000f010000000c140c0000300fd40300000c10c003030014030000104001000443001000044400300c000003000041700f00351100013303170400004310000c1004000c00000304430031c100003f00000cc3100040000340034c0000100103000100001001004c131030030003040100;
rom_uints[90] = 8192'h71f5000310500c0071004043c5010c11144c71cc031070000000d000000c010100c30c05334d00104c100314130c0000c0cfc0410000110000013001d1003101c44003c0431c0300340013c000c050000004d014f07004c0c000c3443010d7000030040004074001410014030c005074c0130c1c301040d40700d000cc004000103d030001c10010110001d00030c110d0c10000000300301700030010001030010010000033100001c0c001031300c1001c310000001000000c0c0043000000cd0400057300100010040040340cf5c035c14c1c3141070030df001c31c40030007c3003441d4001000500010310cd304500310003000000c00f030c0300500f04c0443c303f1071c50330101c000c3003015040c30fc1d303fd000500033c3cc0004c000304040300040f173070c00130000005c7cc30000000700c103430d300000d000040d0c17570c04f4105c0c11503f0d000c040df11f00310f000157300701d0103014503050453f4c1001c040000010c40000301000c000730011c0001013dc3c31010c4710100030040341f30007104c40014030303010d100cc00d43cd0010c003c1c000d0c030733010007000d3105f100714cc04000c04d101003303100d410c503503d451c71000000c0c13c0300300d001413d4131d4001c3f0040703c41030030c003f00054011000f40001dc040ff50411130007300f1000343304014d11000f0100c5cc0301d04c41430c03d3000cf3141101051cd01c003101301003c7c700000050711110c3404007440001f540c40000c1000100400c7300d003040071010000013031c000003045d300d040f3d103040cc0007013f1310c433ccd300040c04003004f000130401dc00011014cc041534c0314d3500003c0c00401000000d0c0101030314c334110003000d300300000150003fc30c00011307047f0d003f7054073cd00c003f10f33010c00314040d4000001017000cc5000c0000004c100030010f1341c400305c05000c4011303f43141400440000c000000c10301300040404100000c3300003041000f0100405000000f331501c000c001d033001300000044000000c01010414030f0100c40300d100000030044d3001051dc14004040000d0100014d0003d01cc003010431cd10050c30cc003c03dc030d00071c00341750000013c7010c333005030001d3c004001015c4c40030c140000f000c40101010410d03443d000350000003c314050031003c3000050d3df0c53130300f0040d0d000333fc301d040053140004100440f100f000003f31300500400c004c005c0433500550005d00031c0c0f0040003004040f1c0030471cf10c3007cc4000350007c10543030070c000400c0000400c5c04307701d0000c0c0300004c0744d000310c00130300000010100513111100530030000;
rom_uints[91] = 8192'hd100100014400003c0000000000c0000030040000000700000c00000040c003000000040303f00c00040c0000000000043033040300c000400000010c330d00000c1f070003c000000000034c030001000cfc03375c0c001000130c100000000c30d0030110030c30010300000000011001000030000110000c30000000100510300d0f030000010c40000000030000100300030000010003f00000030031040000000f001003043000000010033000c000000000003c00000100000040030300050003300301300000000c00030431000030101100013c000d10c001f00000000000000ccc0000040030000300c030f400010000000000003000030000000c10000c03300c000011033010c00030000004f100c4000cc00303000450c31000100d30f005007003000c0c00c1c0043030000507301000000c000004000d050c0c301015000413000000100c1d00000100300001c0000300c1000c010004003000c000040000000d4c3c040450001030c00030030003000017040d0001300d000303340c300cf000000301004c033030303000100c0000000000000050001000000305000000100000070404100f0c03043c0c3ccf4c00d040010c4000fd0f0cd330040000010001030110c000d00c00001030110c000000000c07040c0330000303c0000003010030030000000130300004000000030003000000d0040c3d3743000043000c3000000f04010100c03c000000c050300c30000000300f4c3c0c0014003130330403004103000000000f3000001001300001000004330110010010310000040c00c031003300c030010010014300c300c4000034400000000f04030300010c00003503004000030000000000300c003c4f00400000000f0000140300c033000070001000d0df40404c040c0c3001303000000c0010000f40010d150003000433400001040300c100d003003004004030000301f0030301c40000101c0c1004000431110004000141010c1040003f000c00000030017010000c10000000040300010000043400c0000401000133044040000000000c00011f000103000d110704000c1c0000000000010c00500000040000010c030c140c0c04000cc3300c00000c03c0000000300030f0c000c1000000000c05040c0710040c000000000000040010d0300000101c0c401100c000100f1000000030000015c543130400c0004300030301033dcf0000000c000304000c301000000000000001000400000030000c300030340c0c0c3003004100004001cd00005001010c330c0c4400304003004fc1400000d0000003c10000000c04000c0001300c000003050001040140c40c1404304031c400001000c010100c4000c3000f01000030001000000000000031c00030001000050000310700003040010030f53101c4334000000;
rom_uints[92] = 8192'h1003c001c010013043010000040000010500000130000d00003c030001cf30070100071c0001000003c0001007004330c00000110040000c703000000400c00c4003301300c000c1c100301500014410c13131007100030f00403c300cc304d30300400d03000410031c40100001070003300301000c1303010cc434cf00040003000000110000440000300300000000c011000300003003c0030000001c030c01c0c00000007fc011c100000001040000f0430000014030cc10000705004003c0110100144001100041034100300130003003070304103005f3c003c0c00c00000500c0d5f00300000c01700d03c00003030c00030000011003140430030000cc0310c7530001c000040444301c000000c7031011000303c00300013c304340033d030007000010300100000300010c003101c00001000000003100000700040400d00001101d0003003011340d000034010001405000f1c3f040133040d1030303c300070300030f00101d000cf00c3030000101c00000c114000c0100030001f0110007001000000000017c007000050001301000c000040010000101030c30df000000d1003010110000040401c100000131300303c0c000003430000c000034000c040000000004000043000030010c00003003030c1441011c31c4f30000c001003034000130300300030100014000c000304001c000000003c000301000003c0430000031114c100003440300f40000000000041f03000c04c1000c30330000330010000000303cc0010300400040cc000010031000cc17000040c400310335001c00000000031003c0070c010011c50401011310003007003004c0cc0000010000370003000000000000030000000140c3003010400330004000001c00003411101c03001c0000050401c000300033c0300c0d00000c30004040000011000c0410131000050043730000000c0001d000300000000401005003110100001000c00000c3000f000010000034000010030100000003040cc00c00d10100c0001cc0cc300c1000000001040300303001031043101003000100000030130011100040100010013040001030070100400111000100003c000f3d011c30c00007030330073000000330073100030300c301d10000c40000f0c7301001400300004001040f00004310c0000301070d00030000030011004140fdc0030104000c011ccc0303000040030300300300f00000014000003330c0431300340307440050c040d010005300cc00000404f0074033d00c00004370000300c3010f0c0040c0c50000030733310f00010037004300004000331c00300000007400c100010104370403100311f001350014000003010700f331001300403011000c00001104003cc000c0040c0dc00000000000c000d0000000010043c1c1cc001000030100;
rom_uints[93] = 8192'hf30000000103000000000000330000704c00003c13000300000041c3030100030c04013c333000001300030f0300000c301c03071030d0d173000100700003000300f134014503030000c0003300c00100000033d3130c000337070c00c043400313f001010003000d0c000071cc00c00040000403313103310103010300000300140331000100400304030031000c14300400000030000001000303000101017110050001c14000010000030030c3330001c0000033c003431000030f0300040170000000000103cc00000133007030040300000d001100000d0043370101000303000337010130040000310300010003c003040103300030300000300000303503001103030301030000310300314000030c070101004f10000103330100310000000000c00000000004300d000000000001100000030000cc41000400030311d0000300c343003000d0c1cfc3070d0400000000010340010103430000c00001d000000000000dc0013104000140001003000000000000410300400f0000c00003010370730077300000000000000c00004c00000001004130071c01000c3000451c03000000010000030300000001300f04c0c00100010303400030700510010000cc00cd00310001c003d0000300300000000340c01003330300100000cf400000c07c0001000000000300000300f103c100001000f000c0000030010f00300313130d104c0730030003c003000001f0430100c33300c070034741000070000001300103c00000000100cc033303c7cf300033000001000503100100f00301c34301001003000100030104000131430040000174000003f04103000fd00c014c00010f01303310c0300cd30000000303000043c041100004014001000000000703300000030031030cd00301300033005130c3010004000dc00003070000700100000313cc3000c374000300013103013410000000cc404003c10100c00c0000c30703000000030300030000430003313000000300110d00010000c403000000045700c0c300c3010000004301430030014f000000010003c0000300c0400d0003300000300000004300000100c0401300000701000303043004000300cc313500033400130001030040d303010d300330030033000000000310403000000003010000001001000f410031430300004000d043d3010140010300010400403000003303000030131100400f00000030000c0344030f13033c00033003010004001100c5001000300003010000c1070d000cc1c000050301041c70c0110300010301014101440000000004030000f000040000c70000010000400000010c000003c35c000d030011003303301103000030c000030d004303400701010c000100000003000100100c03110335070130d1010000c10110c0ccf0400310010000;
rom_uints[94] = 8192'h103004005101000c300010131c03403005040000c000c4500103014000010004003300105f1000c000310000c0f07001550300334f10004000000404c143c000c4740cc340030c050000030411000f00c0c4d1050c5030c30157cc00c0000000cc4c1303004300001401d000014010c30005c3000300040100c000003451c044030c03010030003000000000000c0070c33004030010011300000000d00371030044c03000307f04c0000010000d00fc400053110000c0043100003107c00400014403031700f300005d000004010344000c43300034d0d0c5f0000004c1001c3704400000c10403000700c0411403011000c0d300d000c0000010010000003d31400000430001000fc100100c0033000044c100d431010d730c03c70011440c00f0000000010004c0c0c030c0c000100000c073c030070011000043c00303300f054410fc304100014cc004fc00f3c04510c50000c0007017400f0040f0400300c030033f0030c03cc0074713f0c104c030050004001501fc5100530003c100044000cdc00100cd4034001000030410010410000000c000c0470041040000410117cfd00043043f10041003307071300140010070c1d0c003001000043c00004001000040030045c3110400434050007413300004010cc0c04c000030000077d0034401001cc0004300504044014111030130000c03c000010104001cc10154c3300004c000d3310000000c133037000040c00011431100c0c14000111004f10c40000400cc0007003301000001410004c0d30000c30000400400300c0000440cc1010010100000003110030030040000f401004d30c0003143c05133010003c030000001c001040000c00033000c0000c000f00100d4d3f000300013cc1403034cc0000043704414050100d00005d044c1300034ccc14700054f000f43cc0044c3100c004701000d00c703000000700010000005434440f0c1c001c0c00010400000c34300010df04300000050c1c100d153c34413c1030001c00400003004030000ccf44144c000000474040500004311031143d0c300040010000d0004001043d0030310403c3043010400000400d500100300030500455c00340000700330cd0030010000c311010000f04103000500c31c0307001d300040f4031300000031c03c030001000430044070314000c1574000000101010040030010341301d00444013304000d03c100c01000000000c0f3d1c340f00343c700c04040d3104700d0c000001304030040cd030c013c01150f451000cc30000300003cc0c0cc00310001cc40f331003303c10000301000ff0d00d000000000450c00040cc003000770050c131d0000004001c43003000040030110f0330041c007507317000431450441003041d10000c00010c05d00330003c044040f00c000c100f3010040;
rom_uints[95] = 8192'h1d000000174110003c0c0003f3000c400100410d0303400fc00035c0400f4001030000040f40000007740704f10000330301107fc000413300030004000300c0000051c000d0004003000004c34003000000410c0d33c1000003033300c30010c3004001000000400c010300003c0f0d010301000001f000100f00530f000000004f00c400c30000c403040000004043004c00040001000040034030030cf00043004000000300050d0300c00077c11f004343400000030000010010c30103004f0c000000c14103c44c000c0c433001000307000000034300c0000300c00001304000003100340000400043434c030001c007c30c01003000044440030300c103000000100f000c0000044300033310044c00430c4100000d3003000003c7ccc31100003000c000c141310d00003c43034000001d70004040c30f00cd010010cc0f03410304040000c00001001103035030010d040001410000f005030340c00001c001c7f4c0c0dd01774101004300000c440003030000030104000d000001c00100000543000f4003c0004700000c7000400000001100010701c00040050000d0c441400000f000010000d5c403400c03404c30c00f03000000003703040f00ccccc3330004f500030000c000000d04000000c003104004cf0000000001c300004173000f0010033300000033400f000300040001003100400300c3000110c040000d014cc040001303c0000dc54301010c4033004c00c040030c0500004c0c51030307c1010340c044c1010003f0140140000133000100010400030003c10010500c40cd00c0400030030d050000404c034c4343c00d0311004cc000074c01c4070c0d4130000300c30101040700333143c1c00700c103c0cc0c004c34c40700000131010000000d0403110014003f0f0103f700413000f103013c0f3d0074c000000001c300cd03c1037cc30003c0000031310101000000004003410107430047c30100010003c000c34000c00300c0000004000000c04004c00040000000003053f1030d004005000c05000043c3c0cd03c0003400000001000400000c00c30300013000010c01010003ff000043c070010100040341000010000100c30414004001c01c01c0000040004300044341000000c0040000400c110043c400030c00110000c0000000c400400001010000c1c401000d4101c00030000034044000007100040000010300400104c44d00503000d00fc3000305c000d1c041000c0010000000700000c3c0400300f700c01d0300300c00041010144ccccc000704400301c305c100c0000340c403000700c303c0100000030300000004007307c0c301f4c003073043400300c1c30047010000430340000c0017103000050f000dc000000400073d0000c00301d0730403c0c0001000075070404130c0c00503;
rom_uints[96] = 8192'h31c003000104c10d1303030003003103c3304711110f73000000030000d00030030fcc00c000010001000101c0000000047041404307331040300343000300000300100304730070470000d03003c301130000003303fd30337310000041c0310013003303330300c0033c00001300000000c041100033000003003000433070f0c0c00500010011007000c0c0101003001000000030cd4071c00100c0d40001d4c0c100000314410433000301f0000003d010000004d010d00c073133f07303c053c0000330400000000000000034c13c110003100030c300c00011711003300c00000000c00000000c0371407700433333010c0c100000000000c000000040c34033cc0030403030004103c000c0044001c140000000000003c0010030010300440000d01d343000030103100c30d000c0000000010000400cc100000043001f003043c3303100430001430170000301c00000770003033300f13100304050034c000f0000f0f041c300310000c34010c0000000413003c0040000d0c33101430fc3c03c1304c0004c00300c0047000000d100000001c01140c00cf0c30c101003cc00000000c00333c30001f1000177000004100dc0000140310500050000c000f0000700f0c003cc0000f00004c011000000130031f30010003000443c130403430000f001431043040000d001d74000470414430031c1c4000c030c1f003300cd3340334000001347c000004043003f01300c03c00c3cc00003c0000c000310300300034000000000000000313345c1730010c01100c073043030000c43030100030003f0000c050300110144000000c00000000000103c01c00030100100300100c0f00cc0100030030c0100c00f100044010f00c0000011c0000100c303000133f3000040000103dfc000010c00c1000c0c30303000300c0303000c030033000007c0d0000c3f0040000003441000433f0400031300330174000700330300c000400070000000413000010000004700014000c100041040fc4003c00050000310300c031000113010000d0000730000c0c00003000f04c0404c004000403001c0f30370c100000041f0c00010f0d00371130f0000414000070000f410c4740010c00000403004705100400340000cc30400100c000340000f1140d10100000d0100100303300dc000010103c010073300333000c1c050030004013000010051050c0000c000c00100400000300030c040001100000000100c30003c4700c0c30544000000703307c40000cc0cd101c0010000000001010d00000c00030000d03300300000440000004143000000330010010010000000030000300003000c11c001c3c0000000110033100043c300430000c000dcc0040043c0c00030c3c003010100003040c0000000710f03400010c000033330c300000313300000;
rom_uints[97] = 8192'h30c0000100300001400000000004000c010f170000c00c000c1cc010400c0003003500001000001c40304410033c00370030040400300c100000000030403031000000340000000d0c000000441c300c0c00d0c40344030c000c00c01334c4c0140c030c000033000c45c01000c100c00000000f01cf400000745c003c7010070000003c0000000c00000d4040300040001010004c00031000304c00000000000403403031cfc40000c004073c01300000cc0000303100f7030c0001dc0400005400041c0dc000c103d0c00c50003300014001000401000c0704013043000000430c04104000005dc034d00fc000fc4001010000000c00000c3403341300101010300715000004c4c00c300c1400001303000c000100300c000004040c0403000000d00c3000000c510400c00000c41c3c30400000004c0100430000000c0004000430001004000403c0000cc7000dc0c1010400c0153003000003403045cf104d0001000010440c0c70ccc0c4003001000cc00400044cc000000050000001cf103c0c4c141c00c000c3003c030000010000c001000c0c07cc000000003c4c0047140004000c440047043c000330cc0000c4000333cf0017000fc0cc010c01300f3c00c003fd0000000000040c0c00003050004c1314040cc140344f00000000100fdc043c440500040c000000000007003000000c000000003304c7010300330430040f00330c000cc440071544c0000d00340004cc03c3000cc0333414c4000c0140000004471400001c30403d4000001000000030400c04000f045404c4700c00041000001c0c000d300013c003000c130c00001c40c0010440cc1cc70433fc0100503000030007c04010c0303c40c4003300004c4c00d40c37400000304c0c0000c0403f040017004500000c0000000034400c40c00470000000000003f0400c0000cc000400c400000040c440000100c00c01c00004040040000c000cc00c0000034c040403000f0c0400040000c0000c0005000f0404000010f40000330d400c0300c504050cc704040000005f0004030000000404c30110c0004c10104d34004030140f00000c004013301404700d0cc00003c004000c00c05c330000140300004c34d004000c00140c0c0cc00c430030c3c0001003430d0cc3030f0300400000030f00000400041c453c000010340007070d4c0c000c0c0d000410000c3000130410003107000707c00c0430040c740c030000040403f003050c401c00000c10c700004c300c3c300000c0d04033000300403000c7000c030f00c13c0001440f00c40003370000000000000c17000c00000c40001305dc0c4c40443c403f04000c0000000c05033440000004010c00cc0000010000440054300c000000100c00f410000300040d0c1c4101003c0013c011c4c40000000000;
rom_uints[98] = 8192'h530000001c001410430c10037040000101000330430000100d1703300000040400333430cc00030c00100ccdc0d10100004011053301c000f31304130400010000030700000c0d030000710f00030017040f0000f13004c0c1145300033c003017710400000d00000040c000404310041c0700c07743003c00700ccc3503000fd401100044000340c0c003d000300000073000000c030d0cc40c000c74000510303010040000100713000400cc0500000c150f100000034534d0000c110001043d1004f00c01c3300c3010000000c0d0f000040003c31f00370337010043000000c0003cc0c50c0003513c310000000000334c17c04000010c00030000300003100003d010304c100c31030f03003f30c130003c44370300010f474f0000d400c04000000000030303c4000400dcc303404030031000030c040f440307040313c0040500303f00043d1400401140004cc030c41410d001000000d0d0333f000c05c40c031310030503cd003000cff5004300f0010000300f000c0010000f00077300c33c4334000c0700cd03c101110c40004c43300300c31d000c433f0c000f07005cf0030410000400040110300d0d153cc3c00f0010f13030000c00411334004300030ff30c003f040000004c10007c00003033301300c404103730c03000010040730c44410700c00430000ccf30300100fc04004ccccc0000403f3001743000700d0001100c0303070c1f01c003d0c1030314cc1330000f003f1c000c3413000010c3700000041f4d0c030c0400cc075c1003044000c714c0cc000f310c00c0310cc50014000010730100c00c01014c0030440030337d0410001c000040cd00c0d000000340030004010115d0c00003000003000000370000040005000000000c000103103304014003103c104fc410000c0001d1c004c0041d10f0030cc014030007c0303ff075113445f00f0300113431c0000d0c003c0f100300001030003400000c0010440103f00000000f0031c0f10730fd0034040100c4333301400c003c3000040c0c000704010010400c1c07103100c0010c00c00110d410004c14c0403c00000041000d0004c300c303010105100101c50510050c04cf0d13cc70000011fc14001cd00f03400410000307003310000010003004c0000410030c03400000000000c07c041373c00c0004c007c010d0101cd4c30003000f373ccd00030f00000001130c030100054c04cf000c03045d30fc101000c0000c03300700c344000d040100470f371f403f03001000c304010c0310100c041430010c00c4300c00c5100400300d01141c00d001030000100c3003030300001f0f0f000731000000f441c00003c000c4403c0004050d00041407300c000030001c00c40340fd0fdc0c000001c004010110130030d111070410cc1400011f0440dc03c;
rom_uints[99] = 8192'h143040004300c1c40000400040000440300040f03010504c0100d040401070c0007cc44c30000000033071330000d0cc4000c140f0400303c00030300073000000c441000100400c000001cc00043331400050000013d0c31fc03fc0014430001cc00000010010000013400000000003d3000030c4001000030c40c0f400500000700004c300000401003700c000c03000c0010000000000d040000cc1c04000fcc110017343400010400000000111d100c37000004f0070100030dc1010300004c03030300000013000c00705003c11c00c4000c34000c1c0100030d37000043130300000000041000011d100d3c00110001c70340000f040030000f000c035d0030300f011d0131313337fc41c10303310d04000f3c001001300d15c007c0000dc000000101001001001c00000700cc0c0c031c0c0f004404070040310c003c0000d03c100100041c000dc044030100c301000030305c30000c0d0700000001d0431cc70001053040d3003004000000c000040001410110174300010000fcc03010013003000330c0c003f300700331030004000000030307000143107d044003333347c0010000000000010c000111040004c0000030c00004010030c0c00000100d010f0001000007cc0300000d1c330300000430330133000400040d343010000300050703370404000c00044700000057300000030000040000035c3c030300401400003c10300000304107317dcf010000c040300c000fcf4034000cc30000000040c040300104004c000000c03453000403014d0c0c040c000007030734010c0101c0000004000701741700001000000003000400105c000c00c04c70c003044d304001f004cf030c0104000c01000003410100040000c10403c0033300001004000c045c750000740cd300d0707c0103013433000100c03cc00c0004000307000c04000ccc03c34c010004c44c3c0d00000c0ccc000111c00d0030010334000d000000330cc03030040dc404c433000530330c0d000500017307001000c0001c0c0d00001c011c1001430c0070074c0301000000030d031c0401000000f70100001c000000400300003407040001010037400c003401000401d0300f000043d101c40000c0010003400010014104003003100100040c030c33100000510001c310c140311010000f013c000003cc304000010d43000c0000d0fc43011004030cc3003c0c000c04cd00030104330c01130300000f31000000000df4d10c3405040cc00000010034dc00003030700000430df10300100d30f44100c00040030000030044300c001dc4003c0301070014000034000005400003017d070004300c1334030400000000000300000300001000100c000010300300fc0cf001043040c41044050001070c1ccc410001000001000103cc0440005c0c000100;
rom_uints[100] = 8192'hc003100000010000f0000300f340000c1110400300f34c00004401000540300140c04c11007000333001000030400d1030c3000043004004013c5010f030d3000110fcc140000040000010d00000d3003040c000d0000040403510000033300030f300c440c000000010c0c0c01033031c000c500f00c00003d00000004c1400c0c013041100000011c000c00300003070cfc0000000d00040704350000d1000cdcc01c03000c30c00034000c00100c000403040001000000c0500c033d00000d000c04000005030c0f000c0000cd0c0c00c000000000000130100c00103000000f0000010404000c00c0031c0405400000010744000000030010000334000f0d0000010c40001400c4303c013c100300011c104400c50c1000000030040400040c3010050c50043003300c00040443140c00033f300000000003003000000c303c071c00031c0000000c401c000001c40c01130300000704000c011700104001050100034d00000ccc041c0f000000010100c0000f00000030001303000010043f300c010c00cc0040131000140504c00000030c00000001000c000c0001d70044d1c0011000000000005000011c0404000000330c0f7007000414040c0f404f33330c10300001000cc00003000c00001c0300040c0003011f0003040000d0430c443300053c00030300c0000c000c00c0004d031d04040c10040037c301000000013437010003f01c007c000301100104000400cc400c001d1414400000000c0007041000300d10000000005c0c0f0347300004035000300c1d13030400fd0330d00004000004000f00040001041010000c00030003000f0004000c0003050100cc0c0f0004010c0c0c040c0001000000c330101d05011c0f00030000001d400731000c1d00030010000c0cd03101301f0000c0000000000104300c030c0007400c0c0c0d0c340c0cc407000400cf000304010114010d040107440004cc00030004004c0003040100000001040104100300070433700004c031c0001000030100000000134111000111030c0000330000030310010510000d0100101c001c07c0040cc400040c0c003100000001030c0f04070c040c10004100014010c003031f050c00031330040000040c05070410040cc0400010030000000011100f0110704c010f03000415000c0000c00d03014c104f100403030d330500000d000c0437d0d013cc100d0073010c040003003f00cd03000d0400000410040305c1040f0d05000540030004000c0000100f033cc10c0dc000c3004c1f01000f00000c14cd30041c15010c00c330000c3c0007000d1000031000040c000c00050441130030003313c43c140c0c0c0c141d0c4f04000000030c00010d04010000040c04030d000c040401000000303c00074404070004000c0107005111001d500000400;
rom_uints[101] = 8192'h140400c0c13cf0400c00400400003c0c1ccc005440143c00c1000004000400c00000300070000040c1000c0c0c4c03fd100c0c000000340000000041000c300000403000000030c0000c0c4000d03004ccc104300c1c0000c10c0c301000000040000c0cf050000c0030c01c44000040000000003430300040103cfc300f000040301d00140c00000c000c005004130401000000000d040030500004010c40000c00c0041304c0000314041c100030f003003000c0c0104c3c0000400c3c0c00000c04c00000c0f0040c300401f31c001c100c3c0c000000c300000c4000000c3000000f0c00043c40500000fc0000000003d0c1d100000000007000c00040000004304f0c0c4000031003031000fcc0c1000010400d3cc001001cd1040c440f1d4000001030c4c0110c0c4c0cc010030c30000c403d0401001c470010303c04c00030100d01004c000c0d300030f0c410104f00c010c030107ccd040c104400c000dc7300000003340fccc500c03043c40c3c00043001000100004040011c0000cc0c000d0010003000001f0000300fd0001000040000000030c13f0c0000c000403000c000100100cc0c00030011000cc03700004c040000140d001cfc0c0cc010c004003c0c000300000000000000000000c0414717000000000cc43034000100dc0c07003000140040344404100400000040c0c04000410000001003cdc300000f100000400000003000f000d00cc0c40007c03010340c0003111c04103400d00044030c00300d00113c0000030030c300c010003c0c401c0c0c0003c040000c3c0000100c0c5400c00d00100050c00000004cc00c00004c010f11041cf44000004d4c00c4c000001c0c0000334404100d0c10f000000c4c000000000c03000c10c0c0043400301c000400315300c00f10100f0410d0cf040040f00c00c1000000cc0c4010cc470fc040000014000c0dc0004000000c0010014c030c0c0100470d4000000c000c313c00c70cf003303100c0040c37c044000c001c0c0103000100c40f3000c0003305000d00000000c04f10c4000000004ccc03470100000c040010cc1000000000300000c3051440cc0c40040cc401f0010c0c100c440c4d00401d04000000000c0c500040100c00007c40100000100000000c004cc300000c404004cc000c4000001c040c403c000c4f34040c3c0c1300000000c000100c10d0430300301c330c00cc001030003000f10c000cc0333cc013000f30103c0030003c00000004000c44300f0f4004c40000c4304c000c0c4c10c0010000000010000c000cc00040fc010003000c00003c00110400400100400010000000ccc4d5f00c4004340000d13000c0000040140701004c1c1c003cc0dd0013000c00300c0117c13030000300000c0d030c01300001000040fc0c3040cd400100c0;
rom_uints[102] = 8192'hc30000000040c3c3001000004130540004c3010134000004001030010031000c000f0c4c300400c00011000c3fc00c0000f71f41001100c000000004050001011000f44010c000dc100040131c00c0130001004c4503c00c040303050000cc30c01103710c4c00300000004c0400400331c30c4c3104100c30c3030000440340cc3731c0c0c0000c0000003d0000011d03131300001000c000007000040045303f00f0000c0300330000300cc00c00d310c033000000c31104300010140000310f0c00304000001001430111000330010130003000cc103000100c017c0000003c0100100c3030014007045d00d01001000030050004000004000333100000101c4300c0ccd340c13530000000030010300113431413c000c00f00700d00c003c0f050000130000c01050301350001300c040c001d0000100500003cc1414c0030000340004313c430cc04d00f000c00010c017000c0c30000c10f0044004001003cc1c0401433c031c44c4003001041400001050055000f0f050c700030137434c000040303034330000000f0dc01030300003400c03010033443030000000000cd3000045f0000000c0031170cc0000100340c40001000000133d0cd0040dfc30c40c3040400131001340014001000c3f000000101110c00000004010513050000005cf0010303411000cc10000000000010c7010030001000c0104000000c300000010000c40300cc0304300c0400000000c003400c311103c000003704000005f304000540f00000010000000000000103000031c001c3000503d00001300c341000000030000005c30100053510004303000f0c4000300fc0f0ccc050cf35330c001f04100100101004c303400000000401030300010041f500c00c4cc0f0313c100f00001501130001c3c30133011035000403304404f300000330041410003000400713010340c14d34100001c1004c0000010cdf000300000c4300000410c1403000003c041000130474000003355c04c00003c03100351c0f0134000300403c010100000003000c00cf000cc433c130c01c00000140010c00051100c000010000434c01010c0040000040c1fd100300447010000030c040003400c1d00d00d00004004000700c5101300c001c0c437c00010000003400d000000000010003303000000140014150c0001300010c105040131100c0300000d0000310c0034504000c00c0fc1100000040030040040000410004030cfc440c1001300340f034f100004000004c40fc00f00d000c3000000040f1400103f01fc1c0000704000345130130144104011304000d14007f03045000050300003000140003000171f7501fd4130000000c5100000c40300c0003000fc03010101140000000d000000100014000c40000c50040510000000400400403f03f7313f040f0010300;
rom_uints[103] = 8192'h4000000100f01003000000044001c400400100000000f01000040003cc10004010000001030000130030001c004001000340c0504000000000c00101d000400c04000130c000300000000c4000c41040430d0fc3fc14cc00c00041400000300043c003450000c0004040400c0405d370c00103c00cf0cc41000304030c00400c005341030c0000000300004040010300040300000000000cc03c10c0010000004fccc00000454000c1cf000d410003c00c0150000100011f0c000000d0000000f3000100000400000340030003f043000300c0c000000000f000004051700000000000014fc0000004000d0c00c0cf3c4cc3c0004344000003000000003000030c0005140d4c044000001050400000303003030000c30000c0c00c00c10500c00013000c3030400000000300c4034300400000000004400003040000c03300040000c040c111400f50404103100401040000400004515c340c00400003c30000004c0000c01300fc000c044000400710050c000c04c03304c0330004c300cc4c03430f035010c304c300000001050c130001030300003014c0000f000003400041c34003040000c00000005001300c01000301000c005f00c000c0110cd350001cc3cf00103000c30300000440003000c010000cc0003301000003404100f30c030143f0cd04000407410000f0c00000c301c40001c00043000100000000010000000c000000c0000100103040004011010c010cd00d0300c30fc300c000d0430000c0c000000110000100000c0f00c00c4340030300c1c000c00001000c10000103033f00000000c00c0100014100000000000005c4070f00000004400400000c000f0fc300c0000700014000001c03c0c0010cc40100000cc1400100c0030000010303004000c1000130003f010300007040c00f0040400c00000000cc40c30dc04000030301033f005100010001044c000f000000000000cd0100c0300000c3c000c00000004f040043c0030c00cc0354004103030041c0000fc1000f00cc000c000fc07000100000c3c30000030304400c4000c00000cc03000c0100d0c0c000300300400000000303400000140c00001c4300110f030040000003c0405041f00401000c0101c33000c30c000000c00f03501c00000f003307c005004000cc0301c0000400001c000f0c00003000410001000c3001074000c000000f03700c004300c100030050300000000301000c034400c005000441000440400000c7c00050000000c00c00030d0ccc0c00c00003c00047000003d001c00c00041f00000100103040400000001ccc0010011003000001000000c400c50000c0430003c0005f0050000c10000440ff00030000030000c000c10040000000000300c100c110c00000300c004331c0003c03000c004000cc000000074000cf0c00c0000;
rom_uints[104] = 8192'h44c440c05010cc00c440c00c400050c040000f0470c0c4001c0040c30cc0c000400000000030410000d00d00410cf000c000cc0000d40f0cf0000c0400040000003730c00000d4000001cc50000c4040c4d401c010c4000401c000c0004004c0030340c04000f040004400000300010300100043000000005cc10000c000c00fc03c40d000000030c0004c0cd0c30dcc00c00000000000050041c0c1c3040033cf30000c00cc404030000000510004400014c0400c0044c0c440c0c01000040c0cc0c40c41c050107000030f000000000341000040400000004040c403404040f04000004400100c00300c0000414400cc0f40000c0003000000704000000010c010000035404000310000c00000c040000c1300c004144c003000033005030001c0000c41100cc005c01000400000000cc040c77300300500000f04144f444040100040d504000000c040034000000000d040040404011c4341c04400c0d00040433c4040c010c400c010000010033004040c1030f04000041f001c00040000030c10c000c0004030d000004000700010000000000040004000c01010c004ccd30001500c1000000000c0cd0054c0c10074c00004704c000700000040cc004c0c40cc10c0000050c44401000000400070c0001030044040c0c0f03001c040c030c0c01000c0003000c300004f0030c70000000334004c0050d0004001c0030c00040100fc00c30040300c5034c000cc00000c00004300000c400c0c0400401c1010004074004000003400c540c10cc0434000404003344c0d30c0014000c0000400040400f0c0000440c00000440000c001c0c00c040400004c00504007400c04c010c0c0000000f0c4100000004c0f00f000400c14c00010010001100000c0c443000c0000000001017410c0d4c0040143c3c000d004000044f300c130054400500c00000040004000f17c0040c40100c0001010cc030030c0013000cc0040001cc0010004c040000000000700000003000050100cd0310000dcc0400cc0004000c0cc004c03300c00ccc04000c0f00004cdd40100f040030000043741703000cc000cc0cc504000004c000000404dcf303100c0004d34c0c1001d0000000c140010c0c14000c00c00c00000010000000c00000040100c0040000000004c0001c4c0300334c1c004f000405000000000004440004040030040c000404c10dd000400c000400d01c0d04001c00c000000000000f040300c403000404030400c4cc000000004000c00c0c01c440304030dc00343dcf100004040f0c1c000000004405500c050c3000040400500010000c3c00010f00000c0434c0000404c401044004d04100051f0400c00005000c0030f300000007000c4040000cc0c00c31007400000400300c00005c10044000004100000000c40000000cc00000400000;
rom_uints[105] = 8192'hc1400100310cc003000003033700004040cc000570030d041000040001000100400c3040f4f400f00070303000030044c110000c001d040401000140037003001c1004d000f0010c3f000d10300000043000cd30403044004113c000000dd00400700000f0c30041fc5001f00043c30014000503c5110001003300030003000040000c00010300d3010000cc3001030f00000000000000000000000103070000300010000c0000c010030000c00f303c0030000000010307410001000400000103c00010000000000010000300001010010000030040300040150cc010f3000c000000000301000003c0000c00c403000dcc3103400300010040100000c0003cc0003103430344c004cf00000c0030400100000f0743c10004100000c3f000030404300070430003350000cc0c300c001c1400310000440d0000f4000d01c0540740c0103004010cc003000003101340000000003d001100c00c0d1c350101c000500c0003110cc040c4031d10003300000300003413c0000430000001053cc40373137104c31000010104c03c4057300000000000400100350710310c00450100c1000000030040004100c10004400f100040003000007c0c00d50c0001030c001f0100d30300400000c100310000001cc0410144300301010f00011300430004c030400003300400330070000000014400007f0003410dcccc0004010050c10f105045000c0400303000c0c35000c0000404100303c3103400000f0c010340430400000440010000040d313c0000330300000000c1004130000d0340000050d3400c0301040c000003440000004100000004000fd414003000c00d00000000050100030c0440040000000400030070000000000d3000000cc0710304300401c0df00000000000301035303000c30050000000040000000005c4000171001400c0051c00c00000c140000030010003101c0cf100100000004400c0410501031000300c313000c0070100000100101030007003104004000000ccd0f03300d00000000100d00131100001c000c0000070c000dc400c30100010c0400103010001000001011c0110003000103013010c0300031001300400c0c13101cc4010070c00000003310011000070d0031c00100004c0003000301070000001c00d0000001000c00003300401000011041001f004100104c01300010d7003000030f03010000000000000010000c00000100000c00c3000014003030d3400030000400000c3010c00c0003000100000300304030cf030040000c100001003403030000400000c000030014400000001dc004000300100330f1003403100003000c00010000310110000700010003000001330cc0010040c300400030400d00000311341400130400003f0000c03d010033c043400c03c044000000df0300140001440003;
rom_uints[106] = 8192'h300c0013000004330004f170300000401040303000110000c11030000ccc400c00330003100530cf10017100000033c000007030001cc010000014100000c00c04000000000c44100c1011000c400000100c1c040c001c00000113040340000f0000c410034000011000001301513000703103c3010103043c3140300140043030301c40300000000000030403c0100000300005000113111c000003cd43000f30100001010414014c00c0000000f0144c000000013040003c1c110c1c00000140300000c70101040c003300c15000000f11400155301c7c41700c050101003310000170100130000001100c100000500400053000001000100000000001310c000000011010f00440044c000000001010c1003010c10c00f00303111c07f00000100170100410000303000010c3c7000000140000f00300014013003c0040300c0c000c140005d0000001000031010000c013100100d30001311c1043c000000c30303037341000c11003c01c4fc10030000003c113130030c41034030c30003c040140400400101010000c00007050030000300c10000c0d301304100c1f0cf030ccfd000030000003000070500c00001050001501103000c000000100050030030c00000c040140f01330040c00000014003004303044fc0000c110410040c04040105100010005100030c0050c0500001400000000010000001c00310140030040001cc0010034000d31000c030c00001400010000101c703c100c040000031000d1040c100000100000001400101000000700c0040c00c0011000014000001004c01c000300103c00cc1c00040c01440040134000000110040430c41c03100000c704004c000043cc0c40000304340010004c5030030c0003001003c00c0000000000300010000d0c430c4430100d000031301030011000043c14fc03004010300000300c74000c10040703100310100003c3c31303010000000000001030c00000000400f000000000c30c0000400c001001300c30d0c00c0c010c030000000dc01c00000f0003d000140c04401c07000c0103100d400c0c1003d000001c00c0300003300000101104000c00050c100000300c30d0c0031c100000310c1c003c4300000007005c1000101c00000001100100000330500030c00000000c1003c00c0300300001000743000403300c304c10c4001447c0040c0f100c03100000003c41000c0100500c0000000c000c00000134000000c030400c000c0cd0d00000000300030010005c07043c0f000c301000cc400f340c000c7400330000000004401c00000005001d400301100400400cd00170000011400010040000004c3d00047003d0100000000030040037c3000003003030001c0000303110d00000c0040cc014c0040c00005c04000010000003040c0c11c00010000000100;
rom_uints[107] = 8192'h1f1100000041003000c0c0f4300000000c0c30001ccc3f0000400105300000003000034530000000343000350c00f303c043c0041cdd40f30c00340ccc0400000103001100300000030004000c00000300c00c43300311000704d04000c1010000c1d000d0000003c00430000c00010311dd000c00c104300c0ff7c0f00000c03c3000104004c04104dd00001c000000000040000000c0040c00000000d0001000341f0003c01033050000041c3000f40011cf0000070c00771010d034000001700400c001001000300c030c0300cdd000c031031c0030cc0311005010101c0000010040000c0000300000dd3f031f00c030000c10c00030000100c01000000c1d0040335c51011c04000000c0010441000f00500444cc0400000c07cc3c1c00000ccc00001d000cdd0c00010040011100040c000d00c000003c041f1cc004000f010001c4043400c0040cc01c030d001ccd0041cc4cc00c001cd47c00004300001c000000c0c0001d0104001cc01004c001cc3007054c0304000c01000334043c030c30000001005c01000cd0cc5c343300c0300000dc01300fc0c051000030000c70000103dc400000c000010cc0003dc000c073030c00c000071440004c050340000301000000040dc0001c000c00030000000c001d03c00033000000047c040003400000443c04000cc4303700000f0310004100cfd003c0000034010c305003c0314030010340d10000000000000c0c00c430400c0001330c0c003004030000033000cd400404010100010000001dfc000040000c5d40510000d000300c00cf00c400400000000d0400031100000000030001040000001c000cc0c00010c0303c400f0043000403fd0400001104f73c00500400cc0c00000300d03c00000001c0034000c00011440c043c03c0000f11d0701c0700000000000c0041404000010cc00103740c4c04514c13040000c000000000100c0000000370cd00c0300330c40010000000040c0034000034000034cc3010c0300c40c004040c4000003c004000c00c404000c030003d30010300000c03000030003c000000000c450000c0400004010001c11034000007010033c00300410040400000001000c4001c010000000031cc00000dcc4070000c10001074300000004003cc03040301c0044130000c0000001103c0314003000030d0001404c0000dcd000c00000c1040070c040f03031c0040d0013040070000c00c34cc001d0d0c04c40000d30000cc0303000003d00043000334000c0101c1000340444400005000000000075d03303c41000001cd100047000c00153500000000c10400c000000000030000001f73003c313340c4c3c10430c0000103073400dc000003000110110004fc000c00ccd1070300000f00440041033c040c0c73001000cc05010040000000004043040100;
rom_uints[108] = 8192'h70010005011070045d101000f301101c11100c001000111004103000fc5f00000cf3001f31100007f0cc0000300f000c040c0030cd1c1c000434000c0c10041cc30500c300330040000031c000400c0003011004c033cc44174c3fc4000dcc440cc01043000c1000d4053000000013007c0c45f0040c13c00070c00c3410000340007304300030000c000c50700130c070100000000c00030043c0003047004130f0300c4304c1000330004c301030001c031140000300d003000f13740000010c3310c00c01030410000150040cfc171c33d00004304000001c0c1105c1003f7400001c307030003c0000d010f0d00007000010000040300c0030fc040000013030004f0310c5400c173c3030000c433c0041c0000f0000000731cc110fc040050cc0003fd00040000c30c010010000441400000c0030000034fd00c3f07300003000c003110000400001c0340f00101d0034000130c53c400f3300c0dd000000001001300330413071040d040111003c100414301440400353301c0d4000c00010100f310cc03c0ffc000040000000000440000007c0040070f3f7101040100d1405311700430c033d31330c343011c00000350410f0030000444c0300000d030c040004c0000010000030100110040c311f0c0c0c3c0007000304000003c07c340cc34030404401010c300c400d0c0c00c0c50c0000010000000034100000740000c010c4100c104c00003c70d0014f40030d530d4070c04d3f700c14000030c0000c330000d0003034045c0c31000030c00000f30700131d1004000c330300f0000c00731c00010c0f000c01d0000505c000400c0c003c40100c10001f410000000d1470430000100000044014140d5c00141d11000034000c0000003c0c303c3040000c44d00010040705300070c1110c4c103033003030000500043007cf0c100c0c000c01f0c043d00000401c4111c40000003c3010403003300033003c057c0040000c0013c0d001030c040304fc0430043073f4d330c4400304303c000003c4c3c101000cd4c410003000300400d4530000000405003c0fc4cf103740043340c1dc0044100403f00004d0c00000000c00001000000011043430c00400c000c0400c4c10001c1410000030c000003c3c44f0310100100010c1d00000d0110c003404c01300000404000c000c000437004030010d4c7cf00cc00034c04c511f5f0000035c300030000010001dc000c1044010130ccf401043c0377c0010433343000c0000000c0130c000030150130cc11000d013cc000400000040040004041d100f411014003000d030040000300431c0001c00df00400310007c0407343010c3000013300700f0c400c513710004000fc010100000cc000400040100000010400001443530d0050c004c0400c014040040000c000100040004303;
rom_uints[109] = 8192'hc04000c000000300000004c1000000004040c000fc00000001c40040000040000370000cc0400cc30000000c404040fc0400000000404000c04040c000000044c0cc0c0000c0070000044034000140000000043001c00400740c00000fc3cc00c00004400004000c0004000004400400d00c04c00000000000000303444000400cc4000000003c000000000440d100000f000000c40000004030c0c4c400c0000c40c00000c00000cc4000c330000c00030cc0004400c000400c00c00400000000c00000000c000011000400c0c00c0c00cc00400f00004c0004004c4000c00404000000c04000000c004c004004040100c00c00c00000000000c00c004000030704c0043c405000400000cc0000004051400cc10000c43001c0000c0c00000004400000000004000000300040c30c004044c00000000000000c000c4000c30c04030000300000000400400000005014004000000c40005fc3c014c0cc50400540c000c04000c10000004000fc00000000000000000040d3c0040cc1010c00004000c00010000c00000004404000044400000cc00000000000000400c00000d000030c00000040c00000430007c1000cc00c0000c000c0c0000c0000c0c00c14004000c000045000c00c00c010c0000c0000043100010000004cc000c4c0000030000400040304c0c0100000100400014000c0c1000c4040004c04cccc00000300c030404000c0000010c01000004000400c000000c00000000100000c4c00040ccc00c003300c0000004000c0004400c00000000c0c0000000c004000c0000c0000300000000000c0c00040010c000100c430004c0c000c00000c10100c0040000000100c00000030034000c4004000004cc00040401000c0000004c000000400c4c0004000004000f400404004000c0c403004c00070000001000cc0c300c03000fc30040c00dc0f400c0c0c000400c000404000044003c00000400c04c00001000c000000000000000000c00440000c0000010000000c00014c04444c4c0000c0100000000100734010000cc000101cc03c00440000c4000010c0014400c000c0c0c3400000c4000000000040c0c0c10c4040c0040c40044040040000c04404000000c0004c0400c000030000400014000000c000cc0000504c0000cc0c100000c00c0c0000001004000c0000c0000040000014000000c00404004000430040004000000004044000dc050004000000c00000100c000c1300000c00c00c4c0300004000c000000000cc00c0c1040040c410400000000ccc0c000000000004c01004c0403000c500001004000000000c00c70100f0cc0cc00000400010000000000000cc000c00c004004043000c40c0000000c0c0c034f0c000c004c04000040cc0010000000001000c0c00c000004c10000040034070000cc000000000;
rom_uints[110] = 8192'h3d03100440000013c0330100c100030044000d04003301004047303045c10701010c1fd100041300014110c0001031137500c04101440f17cc0d41470c13f300000033f0010003004d0004433d000c10300c0f010d010300c013130000000fd700cc031101c0c00f000fc0010000013c00330300003001034c01504d00140001000300134003000c400000400f000071000c000000cc0010d104100000c37014c30043000d430c00f00c0000000031440c034500000000c00c01003c000c440030041000c0004c010100001c0004df0101000c000531000000003c000403000c000000011070450000c000dd45fd037040010c010cc0000301000001000000330f003dc0f0430001040001443007133370d14001034d00f00100001f11cdc3000c3010004010010c0c4c0f43111400c00c0313413c43c100104400c00c31040f300f3104431417c4003003c303004c03000dd03f11030430c0c13330000040c3c000400f03430c3dff035507c34f3cd34100400c013c00003c013c01000703004101cd0304400c00c30100000051fc1500000001030003c000015303333307001031000000000003000f0405010f3d0001cf377d00000300000001040c0c40300f000310f0c0000330030130c0000f077500100000d30400443005043c00fc0d3400014f0c011300c0010d00010000001354030f0010300340400dc0300f04000140c000050004100000101ccc000030c0040441000dc7031440003c3f04c4303c40010003cf00d047303c014fc1df1400dc3300300000034330c700410441100013000c00000105400100c130cc0040000033004f41000d1c0cd300c33103c0000304003700030c01410c0000070005cc073013044300ff00d3c0000dc1554f00310c013100004cc0000100007c1c07cc100f03100c33d000000300fcc0c40010305440003f0300130003c1f40000110054410c0300001dc0000011004d3000007d40fcc000c403001c043004d000410001400047fc4310c04030310c037105d300010c0dc5c0001005303c0c00c00030c01d0400300040014100000044c4030c3010000c1700030c0000c70003000010010731c00d03031313407000000d13417c00000100c313030430300304003100001f3c0ccc500307300040f304d4140010030303d041c0d00100f0701d033003003307c1131004031f00040000007001140404cc300000170c03c0f5003100c00f130000c304000301000dc000000cc00101017c000cc00400354d000c00cf3000030013c400403500040530000100174c4331d0310303c0430133d410c0000001440cc70000110000040010000300010104f3103001c4000c11000001000000000300000311140f4410703f070c040300331330400341000101d00000000040000300000300440c43470101c30d00;
rom_uints[111] = 8192'hc50000000400000000004000400000c3003d3000c010c1400070000c000cc000000340cd7071000000c0400000000c33c0c3c4010040c04c000000c00c0013000000033c00d30010000000101303c00000000330f01003000740005000104300c04d00440c0010d010030011cf4040040000c00000c0300340d000101c300c3003005000100000001000300304005330000004000010cc00f00041004740f03410dc4030700040003cc001004033011c00cf0000000010030000c0c1dc330000400100000100404000400003c0131000c03000cc00000303c0c31007c13400400300000040c03100c0c0c0c000d400c0400000003044000cc0c050303030000010404003470c4cc100000003c010000430cdc00400d0c300004100dc00f0303c0031c0003c40044000c30003300030d3404001c0030c00c000000040cf0f000077c0030100cd00000041304144001000304000003c000441c0c04437c0cc10045434000c000000c0000401d14000070000000c4c000c04010001c33010c0cc0000c0f03f7414004300000000031010401000040000000400f00003000c13300003d33c03070000004000010001c003010040030304c4003000703001531000501700d0004d00400000030000c0004001cf03000c04430474000cc101400003c0000001001c0003100c01300c130f0000f000300000c000000c400003310310140100030331000110404070000700f0104041c10043000f0400031d00c70030000001cc00700000c3000100c073000000c14314000000400010d3cd000000c0000000c100c0000c00000c0000c0c0c0c00001030000110dc00010000c430c70d0001000c0100310000405304001040000c000300100c000f400c3c0003103704004c100140013004000c0c404040100400c07003000f3040000c00000410030d0c00c0cf00143000000000031000000033c10c000c000d0000c13701400c014031040430000000000030c00101043cfc00030440070041300f000f0000400c0c00c000050c000040004f100014f0501017004c043000000300f0007044000c010001034c003000d431301430400030030400011d114000300000030cd04d30dcc3003c050c14c00303c03100cc030cc0113414344000c0000cc000010100003c0c0000000c001703000100071400f400f00100000010400005770000000f13400003100001c03000041030003110cc010304440001053300040cf000cc0030cc01000c00c000003400000000f000cc3000c04470000000100d0c1c143000000f1c0c04010c004c0c040c000010000104010d00000c100730c0043500000410c00c01304304000000c00000000c0c010400f400010001000c30300c000c0440041400c00000c0003031030cf4334d003c00100c0000000f001d0000000c0000000;
rom_uints[112] = 8192'hc0041047c4cc0c00401c0073700500c0004000c0c00000010c0c4433d00000300c00c00100f04075c100010000403100cdcc00c0c0c0d0cf0044c30300c0c0030004c010c10007d1f001c4f0400c404003cc144350d000401410000030f01000333f73000000c00c00430000515040c030400301c31040400cc50110004fc000403ff000370004c004c000000003cc44c4c000c000441040ccf1c0c0fcc0304c0cc0000041004470400000fc10c00dc01000c000054340c13000c0cc00c00005000010d040cf00f0100040c0c0c35130cc41300000c0300c0f40300c01c04000c00000c103000100d000c00000c440c3c007000030700040c1004030c000405c40c3000c007040000cc0c00cc000cc0d04c70f3c40c3cc4dc4400400f0000000f0c400004510003c0fc0c0cc00000c0033000000c0000000c0c0c04c13c470c0700037c03000c000f0441040c4c0044430035000035313405ccd0350c4400300501003cc30f303f3d0000410c00000c30040c0ccf4c0000103cc400000000000c0d40c0000c400700000000c30075c0110030040000cc400003010c0000030ccddd4c01c10d00c40004030c0c54cc00000000100c0410000dc0033cc40c7544000047007c410c050c0000c3c0000cc000000c040c00f00000001000444cf0d00c000c1ccc1c14050c3300ccc004c400c40400c030400010040d03100fc4050dcf0c01fc0474cc1040334000000003740404000004403cc30c04103fc57135c3045c000413fc301000330c00151010300c0c00c400cc07300f0400100000cc4d0c00300740030c00040c00030d30c4000c3000c000c00c0700011140140c0cc00cc40000000c040f0f00cc10d004000fc0400f0cccd43c0d10010000cf0000010400300100010033c4100d03c30c0d0c7007c31400c7307000c404413c010cf00c040c100fc1440c010c04df0400130c43000001004005140c000031000c4dc00c00330ccc00040000000013010c010c010c003fc00ccc00c10c4c30070ccc3c3400000cc00005cc00070c0000d430c40c05cc0000040004cc00010c040044004d040003040007c0cc00400c0f0001c0140f4000400015015041003c00000f0003c000001401cc40007414000c500000170404cfc0140cc03050410c00cc001401dc00040c040c34400c0c00101c01100ccfc003003f0c0c05000c0cc5400d430001404c0cc00051c40304c0000c0c00030d000ccd040c07c4140004040c0c0330c4400c400c40c0c0100c3c07000c01c30000453030040000c4c0003400004101300400cc000d004f0c0c41000c3c0c003dc00c4c004c054d04d700007c440400c00c0f00cf000c0003000c10000f0000030010000400c400c00d031431003c00150415c000040f040cc0030400040040030c0c0444cc0400d1103c0c000c04;
rom_uints[113] = 8192'h34c0000404f040400440000010c00104d0404300041d1cc04030c004000430000300400410103c0000c0000050405c40300400d010c333d15000100430404100c00000000c100070d004133140010c100004310ccc130c100000101000cc0040cc303c13000c0043000c000000044c0030cc0100c30f00000013401034133c0c7004c010000000000000000c400000000030000000100030400c1001c300c13150c01401cc00c0c000103000030c000c004004c003c0000300440000c0000000c010c010001300c3001000000001101cdc400c3350c13d0c107c3c304440000c000000004014400300100c50c140f000100c0c4040000c10000000000000013100c0300000f01130005000c0c50001c4c030000c00307304cc000f1c000003001cc30000174014c0000c400340000000040c34c1030cc40000040c3400400c703400001d1c44fc001000cc30003c0030f40030050c00440303001334001c30700043f00c4440040000305c00c405cc040000003000c0300c00330000cc033c00c0cf003d11045010c500000cdc000140c00c301d000c404c30300000010c04310c0070003ccc0400003010000304c00000c407cf0040dc00c000c000c00010003030c0000f004cd44004f0d00000033fc0000c00000430000030000c013c3c300000040004144c30404c03400000f5cc1000053000000c1405100c1c00c00d4010d01c003030141c10011000fc0040443041000430100030703c1c10003d00d01004cd10404c0c7000410c04300440000001000010c004c010000010c0001004cc4d140010100000c4f0030c300003040001c00010101f007110043030f03c001000004c301c000000070cc0004c440c30ccc044440470300f0040001003000004007dd010000100000030040c100c0330003c0c1040f0000f110000700c1c05fc001410cc0030010013401c344c0000100050000010cccc000000000c0c00c01000f0100000301c000340040cc03000001000300013140070c3050c30c034100000350c000c0000004c033700040004000030d40030100030003407f430c00000c030c0001000d03050c01104700030c0c340400c403034303000c00c0010041430000400f4c00037c00050000050004030010c0c00003d00303c0c0c307400040043301004007c0c00c0030c00001000400700d1000000c43c1004c00c10000c040000d00000000403c10000000000c000c1c0000c0c1cdc000c500000300c0000c00cc00000000000c400300014004170c700004000007d033004000040103000000440000330000cd0c44c100000041015c0300c0010000010000c1cc3c0300c00001c03000110f03403100001001000cc0403000c4c001000c3c341000430000030cc330000053400c000003001d0400000003000d00f3010cc0003100;
rom_uints[114] = 8192'hc0000c00c00014010100000c0100c4131505400410001f0300450d0037047410000c15cf4305c1c0c44cf000c03cc10344003053005cf003000050033c000f000470c0cc005004031c00c0c30c0013c000003c000fc00cc4f0f0c30c40034414d0c103404cc030c0100d0301004d003c4043003400000300010011d000310f30c0cc041010400c0010c3030c40c0500d000c0000000014ccc400075000301c343003044c0c001dd401000070c00c0057000003000010c5000cc300c0100300cc40070000c0034c004c0c001000cc3cc40005f00000d0c3c000440d40c44c0cc0030500000c07d4000c13030103f40d00400153031001000000040000000100f051c3030130004040400f4513c00c00f0c3550400fc0c04000c110110c1500100c05c010010000000004cc00c4400333000170c400c000100000000c04000d000000000d30000c00000c0c0cd1000130151400000431707405000043cc00001f031c003c30113000730501401030cccc30030300c00111dc000400013c0c7f0c13010030043cc0d034000400cc3c34df400000000c0c00003050334fc10f0130cf450d0430030000500000410054000000c300c4c10411003400f044530c41010c10400f00c00000030f000004305000740300030d70153000703000100503c01040000d001013133dc0f3d00c0000103c000431c40c00400c3000040107c03f41000c4c4304c0000ccc040003307130001c40400000c40004400d0040104c300014f71004100001c00040c00f00303c0303700000013053004c0100c010000100000f0cc03c00007000107c00000300c004c00c00304cfc000fc040004000c004f0040000c01c40000100f0cc001130300000cc0000010030c30f0004c73c0dc0004014c0cc000ccc000000d10111100f0004f001000c000001d01003130c300414c074c13c3114c300c07000c4c034dd007001c0001003d000030c0400c0000c317010000000000c0010430030400d0c000d03031030fc00300130340000400c400003c50000c0410c40c04004044c000300f07003310000f1c0700343011304d014cc44cc410003004cc310301d00000430434cc000d030413d143c0f31000510d00300003c7070c0503c0c0030400000170cc000d0004040c001c00d4300000303001000503000150c1000c404000070000cc4c00c04050c31c0000100003040700c00ff30010f40c0000300040003000c33440c0130000000040c400c03030113f340c04300000cd004c010cccf00000000c50fc34000301c000f0001000000c043100dc070c004003000000040300cf3000f000c300000003000014010000000403100340440301c0000ccc030000000c03000000c70040301307f000400c0d0c30414c000301000403000044001f00c00c0004000cd3c3c70340304101;
rom_uints[115] = 8192'h40300c0040000073300000030c003c00c00044004000040000000100cd000000000040300c0000100c0000000300f33c40100444c300c013000000000000f0001000430103330c400000000cc100c0f40004400cc0c03000000403f00303c070000d04003440000000000000000004030ff00003c000004c00140004000400000f5300004000000c01400000300400043051c003000030c0004003300cc040000c004400000000000000040c0400100000d0c0000000c00c000000014f00c0cf0cc40cf00000c410000000003000300c4074000000000000f43000c134400010031400000c300300003000f40307000031cc100000c000c000f0000c000c00c0330000130411000c0cc0000100c0c041c04000030000030c100c0c0c0030000c0044c0000cc100030010043030c000000010040044103000c4c000044f7000400c000c050005400000000000000c001000000000350044043300000000c000100004c0c1cf1000013040044c00c00034050c300dc0d1c0c050400003c1000030040c30100c40000cc5003003c000c040140000000000440040c0f0c04040c10100400d003c40000cc000c0444440d10400305cc00040c40000400d0400440414001010c0c0c000c00040cc03c00000000c000000c0400300010c040004004010000304c0004c30340fcfc304400030c0ff03d410cd004030000000007c00304030c3300000c043c00000c00c3c40000000c00000c00300003003c4030c0c300000400430044f1030004000000c001cc0000c040000001c4c1cf00c00c0000c030000400c00c000003000c00000c00000000450030000000c4040000000000c47000140030c1c004c0c0c000014000c00000004d004c01400c000000004c3c00003044000c3c0001030c37f0c0f074003fc001100f00000cc00000400f0f13c0c0dc000f0703c00c00c3404d3044000f50000000000c400c0c0c003000040000c000010104c0000003000041000000040c000000004c000100000c0000000d334c400c01c0000000010040c000100c10c03f054dd0007c00000010000c1ccdd00400c00000d000c1000000000000000c00101c4040000d00000031507cc0014cc0c4000c034c01000000c3500001000070004c004003c1100000000000cc00003c1070001000350c0007c000704003c0c00c10c100403000430000c00000cc04500040c0004040000c410001045300040410c11004000f30300340c34f00c430c000300010400c00000000007cc00000c30000c000010040040340300c400000000000c00c0000700014c041c00cc000100f0d34010000d030000cc0000500cc4001c005c001c3003000c40100000000000000c0c000c00000c0000c00c0000001c00000c043c0000000c000001400c00d000000cf03cc107c000400000000400;
rom_uints[116] = 8192'hc00c00000050c00000400400000000300000140000400c0030041c00003f000010143000400000000cc00c00cc00040300500034500044033c10000ccc0000304000000004000c0004000004305000c0c4040d00043050c0301000300000100c004000000000040c000000000004331010001030001c003c003000040000f0c03c3000000040001000000c30000c000000000000000030000003000033c4000c300c01000433100010000000107c0c140043f01000300c0133040c004300000010000c010c0004400000041030c01000001c00001004c000045010f4c0d00040c3040040331c00000000004fc050cc003000cc050010000c0000000c0040040040000000000cc010c0000c000c010000003000000c000c0c50500033001001000c0440003f000c44100004043cfc00400f03001410003000c4c0130400301000500c0004000c3410000000c4000c003c004c0010c0011140130c700c0000040400d001000000740000143430014c00f404c0cc00cc001000140000000000000dd030000f1035000031c400407034c0134c00c0300000003000f0000c40300cf044100301000c1000300000041c5001304011710734cc703c40441004003d000030003000c104403004000000c3000100d4000000300c00000304040004cc00c00000000f1c40300c3040004c0430003003040040c500000000300000cc1c00100000030c3401cc70010000d0000400c40c4000003300011000004404000c3c00001c1004c00c0000000c05000100303005001cc000100014001c00400000001c100010cc300c3000030000000404000000340f00400000000c040000d004c00fc0300400c050330000044c000000000004304001f0000010f4040100104000000c000d3001000030c00c1c100c33010400c004f000504c0000d0301001700c000c000c50c0004430000004040030000c0c00101000000034c00000000043001c4c00331000003033cc00000000c000d700c010300000304f5ccc33040c107004040004000f0030040c040c00000000300000013c0040001000001044f0c000000c400cc0400040040c00303030030000f0001004f110305c001000d00c30000c30000000004d34010c0000043000100404000300c0f030c0c05004143000f000c04004001f140430c030c001301000000003000c005030301350003000001030300031345040005000c0300005300434d00070100000c00c00000c00000c100c00ccc00000001000000000dc004c0c400c0000c400300400000400331000300000000c30401051f30100040c000c10f0005030400d0030f00030040000003f00001c001c300ccc110000300410c30c447010000000100030000040401fd0103400c0000c403000f000300d00000103f03000001000f043c0003010041c000000;
rom_uints[117] = 8192'h40000000004001044500440c04000700c0000007c0c13303c01d3c400f5030000f31c0c040ff33000034070151031d040c103030303d4c04000000030400400031010131000c001300001370100015c00c400010145c0d0043cc011500014d0f34170304010050c00c00c0300007c1330d4003c407ccc104000c003c00c31c03c1401d1000100030000100c1030c001c1c330110001c40001500dcc40043d01c0003cd03140c050730310c1c030c00f00153c303003010470c0c0731c1113000030f0000000030430c7400400000c531300353030c3c05000370307403000104000100f010cd03000005043d343c100003cc01014d1f00c00000104d10000003d10000000141004d1100130f10c01000003f0001103100004410c5304434014400303100110c010040000000440f0cc00040fc31340000300003303735c103400500cd30400307000d417300400001003141c0f3301c1c0d0c0c1dc10300cc0cd003330045c0704130011330001c71073304c34c134c0c00700c0c0100403310c403cd001c33c000c101c00c510301d70003c0c100003c0c0303d00300011ccf0701010d0003330f00041c001c7370000307310011300d0c330143430504c0f170543407401001d0300437000400304303010710c00431d40c050000f0054cc1cf41000000f04400c440400074071005d7100c0d0004c7304c0d10010400f0f400cc134013c01c010004c1050340c00c100330311c040d05043003033030f100400330000035000400440c10043030040cc040c0c40107f00c000000100004134007c31c001310033341001530f0030f010000300001340c3401000c0440073130000c001f3d0357c144000c0010004c14030c030c1301003047100110010c00000c040403cc0300c00343400000000cc73301d0004c40c00c1cf0004d04003fc00d00010c00400c03315c0103d11cc31c30030c0fcc04004030304c00000c0004c000300000c3010003003c00c3030300dc0104030c0cc130040000d0000fc3c0001000f000130000c3300704307c0104003c10000010010300c0c0c304013013000cc34103500077100f0004110fc0c000dc0c3040003f0004003c010351050d010c0404305003000043030000c1100003470410d000000333403d03c0070403040000000401000c0300003044ccc10304c00c00c303007d00111001f0d300cc0003340d430c0d0f03000010000c0c304040300004c700040000430f0004f3f40c10c0c404f30700d0304100401d300f100d400033030070310300000100000d33030c0040010330300701d01000c300010f04f400140730100000d30d001004041310cc540c0cc0003400c03300001c004000040007330d00070f341f01d0000300000c000001035c073030c40c100c003300030701cd7d3300c003000000;
rom_uints[118] = 8192'h4000104c0c0000140c000434400340c0330100007001c0000c3503003c30001c00c400330000003000d0000013c3004300f3014030704010000c3f7400005000c030001c3000010000000c0d1000431000011d033c500400f0100150c000000c010c303c0013311030010c1114100144cc0004105003100c050c10400000000f33000104000000140040004c004400d4000000000110000c3000040103c030000000f0000434000000403400153000001003300000000000f010030c30f000041c50000000300004000000003cc45c10330004c3100000010c10140d505110005010000c0dc0c103103c0c30030310c03000fc400010000000011430000004103030030d4d00073300010050000000400c0c0c5047f0000c03100000cf0003105004000cc4f000cc410f04130010c10430301cc05000100000004005004050001d01014000110000700000d340c4003c00f3001730000c0c1030040c0000071100c414745030f00c43c000300c004050031c0003040cc1c503300c01fc00c010300000300450140003300df1000c131100000000100070101c003000cc00000000c000003000433000f003000400cc00000d34c00040500001043430100f304000d034d00cc010c4001003133004001d000c0cd00153030300030000003007d05003f100003400047d00310000c000305c0001040010001000010c300c400d010400c07000000c30410307017033300c100d14303014070cc0c1001003311c140144c00c0c40440000100000004130c050400300040104134000043100000c04300004340c04c0000000300f000f40000401000104c730f101170c0c4003033031c00300030000050004cf00f0100400c00f3014c00c000000d040c000f10010003000073cc0c00000011001403cc4310f43300010303c0000c030043410004d130c074010c40000104000001c0103cf0c4030c0003c10d000033c00113700c30c013cc0000000001010c0000c0003cc00400040304cdc0cd403c0f0143000c0000004000000000003d01000dcf000c00011304030c00000c0140400100c5000c030003cc31000100000c00073011004004000301011c000f404c0001d30010001000000c100000500000d0331000000000400440410cc00c304ccc40404141007d004d33000000000f00004330004000401007001010404303000000000303c30c044c03100010400040d1c0000003c400151400040400415c001403340000003c3000000000004000000c01404011310440c1f071c000c3000700d53c000400c1c1004cc0cd500740004004140103007300000000030c010c100004034cc30cc0010400c7300100000c40c370c010004c033c000d0011d004d11f0011000070100101c300000300cf1000c0c00f00d3300010000040003010030c03000000;
rom_uints[119] = 8192'hcfc41000000c0000300c0c3010c0100010c30c003cc0f40c0001d40c434c0000000f101c041500100000001c04001c03007070030c100040140004503c400000000c00010030c000000010007000500000c0f03300c4000000331c0303031c17c4300070300f0000003053c0c000003040000003030004c000c00300c00010f00f0040003010000c004c5000101051dc00cc400000000040070000c00054044c1010c500000c7004010001011010000f0031370c000010400000c004300c0f4cc05030040003051c1c04005010341000cc140010403000c40414d000001000144c1000c0100003030c3000c4057f031003cf0000000500000c0400007f0c0000c05c00003310440110400453000c00040011f50c00c5000c3f04001034034000000000001100f3001cf000133c30cc3000110c003c05000030000034000c0c000c00001000fc0000040000c34030cc0000034700100003104c00000014000000007000100040003000101ccc300c100010c0140010303c0001ccc030051000c010100c140f13c0d0f70c043c003000400400040300000c00c0433014cc040000303c00000c0300010c01100c03c000fccf140010431011100000c034441704000c0000471c0f0c0001c143030c3000100003004310001c0f0430000c3073c03cc033ccc0f00130c0304c4000304c040043005c10040f044400d0c00003cc134cd30304000114cc34c0100c1037c0500000cc040d4000d50c0c541414c1334005001cc000700000003000c4c4010040000044cc04301000cc00fc00c034007c703003c4300004f03000000c0c30000c000103c10100c41cc400fc300040c00c0040000c00c0010cc000001c033000101c301710400c400000000030301304d00c0cc517f03c0cc00040000040010c0010f40400001004000300040c00ccc0030c3003c40000001010100c3f7c1c301c73000c3000003034503300000030c40c00303031f1cc00f010403c00300413103000d00c440404c003cf3440c040c01d0003003c000010403000131034000554c40c00fcd0003c44003057000c0300c4003000133000c0c0c07c0004d003001f00f030040400400cc0c41000113004003104400001c7044000000004340000fc04401400444403f03100c0040107034000003400c00c300c3c040400303004333000000c1cd0f0000050701400cc000300f0c004f4fccc0000401110043c100cc010045f000c4c1400000000c0c31cc434f000c0000c303f30011000010c10013000303070343000100c30fdc00c500000f0533fc11000305c000103010000000300dd0100f0000030303000001001540000110400000d0334000304cc040c007430040c0530004c0f030040000c0030100400000040300010000c330000470c104c0c0c00400000f00143044f00000000;
rom_uints[120] = 8192'hc4034040c0f0300010030000000000100000c030c00040030033c3000f3003000000100d000040003cc0c0c10140100cfcc00051f04f00400100000000001000000000430003c0000000300050005100045130000050103003000043c041c003305c10c030300003054051000010003050c100500043001000001030400c00c0f00044100040000040310000300000043400403000001c00030301f044104040714c0003000c01f0430033340d1fc000400f00c000301c000301000000f0000040c101000030040000305000350041000030000c31c30cc010144111c0c000c000010000d003000001100000001300f00410003030030000314000c0d0c3003010c00000003f50030000f01c0010100100014000c0705300c343031710031037300f1000400000c040c000000041f070000150c00010010000c000c0300310031000501103c01400f300010c01004c10403000c00304400c5d30010430110010530000f010000030004000f1c0c00440301000c330004000c401301000000000c00c001004c000c1f041000000305150300057c03300f040c300400030004030f033000000f4000300100000004341cc00c03c40000000033010300c30011371013030004f100050c0400c000cf00000c000c040004003c00040000170000050c0c000100300100303c01300030000301340000000000001400c00003300400c004040004000c000d0000001d010d04c00c0c0c003000cc403105000400d70f000034c00100300f0000001003000000000c4d110043000003010000030c030000010400001030c00300000303310c0c0000000001000500351c40000d00000f0000000501000100000d0c00c005000c0003030030410f300100430001350c40000405101cf04404c000000100100d100c10504501010c0c0000cc004f000f030f15c30000403500001c0444c5c0300004001f00440c040c00004000003c0403000000040000000340040000040101000000010015c00040003330000001030105000c004000111701000c000500040303041000500001000c0004c0051c01010c30000c403c30000c000001c0000500311300cc00100100000403030c300c04c5010000010403003f00000000c000000104030504c4000000c104004c03051003000005011c0c0000005303cc04000303031001000c000c3054000000c1cf4000000300103c00053100001300030330000f00030f0c04c00410300000400c000010040c30030f30030c0f003103c000340451040045303000100c3304cc00003f350400f0f00f3300c0304005c00501000400ffc0000c000f310000000c000300050000010f04c0000010000000000010300c30000100010000304040000c10003000300100050c05004c34001001010000000000000000010040001c0030040;
rom_uints[121] = 8192'h743003003c0df4041000010c10003100cc0000140001037004c3000030d300300030c04c307400c130003044010c03d400333530030003c01c003030cd0010000134705003c00000c0000d35dcc0100c403310d1d0fc7000c040400c03307034401000004c000300f0d00c0010d00c00441074107044ff0d101f01c3cc0c3000f0333d000443000400343c00df40101c0000003c0000003ccc30000cdc5f0040101041000030007403000330740d04c400513f00000010010031403c30f0304cd074000000003c3100dc00c00030100030040c0000300030134074504400100c004000000c3040003000000000300c0030c05303700300000000010100000003013130000c0050037c1c0370f43140001014c44c00f30000710000030cccc010003f00001c00f1010310300c430030100000003703c1c00040c01000050440303000c1700001fd000cd03400c4c033d0103100703c0000404437130dc30103000013300c3c0000003370440030c1dd4010001c003070c0f0003c1030300000100c000030fc0134000cc00c0c00001001c100f00c101000400330c4301cd00f0cc117140c43304011c0c070407734000000001cc00dd03c3c000c10341031cc147510100473333ccf0310403040043150c4c0001030113c0c04100400103034103434f0f530cd10c0c070037100c4cc0110001cc00f00000c040040000000d0cc3c00043c0c0c03003c503001c0347000507010c0f10cc1000001100300cc301c100300000fc00030017470100d00010300fc00000070500040044530100000000c0ccc30300000000c3030400300000000030c0f0d70303010c004f01140c3030c0f0003007000c1000dc000340000c000f000440001c13c00404c0000004c1cf01030030c00c3005037001c35003430dc000cc00010014f003000401f0033300c730000300100c0130c40505c001c0c40000cc000001030000c003c30fc0000f0c00074000000010c03000000333130114cc3010c00f03cc000100300305d4350000c00c340d030005300101101701300dc00f000c030003c010000447330000c100000cf0c1000004300c430d100001f003f4340000100044f01400c1c010030310000c3300100100c00d0300004000040003c301c00700c40003401031401103530143010005003030c100cc00c040000d33000000c001003c0013030cc30f0004344f001040103d00001ccc004cc4c3030c044010c40d3000010c0000d0313440c0300000000500070ddc000400014ccc01010031000074030105004c4cc0f71100f3000370070f0003003000070303000000000c3140011040040040d3010d0040030f000703000155dc3033051140010c100040050c0f400004403c070000c0000c000003c10d1750c0004f0000070040c1050001f340c003107000000;
rom_uints[122] = 8192'h10000000c003003fc0100001300130d001014400f40440311c70c00003001000000000003300003400500300f0010040cc0cc010400004c3f0040004700300000000001000f4001000001101f000c0100000000300500030304004003100c0fc443030000c100030100c010407704000d00030300cc314000030011000c001003000004300f0000300100000c000000c033000c0003d1100c40003c3c3000c0000004c0000030004000c0014054104301100300004000000c0000000c0000f0400d0c000000c040c03100330f000004100301c000400000000c000c00000000cc1100044d43c000c0440410431c0000000040c400f0000000010100c300c0401f0000001000000100400000031014300014003c010c00000075011c00401130000050000f11030c030010000011040300c000000000000004100c100f0fc0003040000043c500007000130400c10000c0c00c000304f000010c003000d0050000f3cc00303034000300100d0040010403000400040400440101000040000c00003c1300000c003005100000030c30305000010000000c001c300044000000400000c000c10000c0043d0000471040c47303004011cf100100403000404034001cfc0044350000011c00c30000305001000c0000003000f0410003000033cf1f0f0010000c001d0000d0c40cf0cc4c300000d0000450400100400000400c0cd140040003f0040c4004330400c00c0000303d000100031000cf001c000c0334300314000001f30c0040030700003000c4000c104000c3000c000000104000c030000000c3d000c500000c00030010000040c00f104000041030c111003c043300030000000c00c000030000040000054001430004f015103010cdc300c03005040043f00000000c00003c0004400015001030cdd100d0403000003000f0c04d0cc0000300310d0c00ff11c0000001000000000101500040000400c10f00430000d1000004c00000700f10c000000c43110000034030000d33c34040c000100000c1000000c000000114c0043000000300c330100104004fc000430300fd1cc4000000c001c300000000003c0000c000003500730005c00000c4310704c10c000040040001003030000000530c4000030700c33c0000400001301010000000c010000000000c0000c00000000430c103300000001030000343c000000300100c0043c40014100c00100100130030030100000010000c33040c31010301000c3043054100000700000003430000ff03c010000c000000000700010010000710000400000030040301cc00034004004400300004000004000310400c00000c0000c0c000c03f1000010300340000400700030c0000040000000c00400000003310000000000040c00c50ff300c000044c00000000005030100341530000000000000;
rom_uints[123] = 8192'h30000000350d0000c000000f3100c030c030113c04430500000f3000040c00000000010400010004001c04000000d0c1000100400f1000300000001c07c004000c03041c10000130000000030400000000100d010dc303cc040c0400040c0c040003000304000000c001000c000004c003400000104c34030c03305d03c004004303030001010001000c000ccc000000c0000000000000410d0301000103000000c00f00030010c11010000c043000550370000100000700c43400001c000000cc0c000c000c010440010000c0003c0000c40000000404050444003c00c000040303000013c003000c0d0c0100100000c0c03001300000000c0400040c0000c340033f04030044041001040000000c40100d030000c40004043000cdc414033300170000444d04040040000c0000cc43000000004d00030000000000100000000000000f10c7010004000010c4300c010c3d0c00d404403000003404000c00000004000c000003001300000c00c4300c004c040000dc00000001000404c00c000030c100c0001400030c0000000c0cf5000030010c00403004010004703005c000cc0d00000c00000003300c0407400010044004004c414c000700040007073c004043c7000c00340c0d0003fc000400010000000030003c000330000000000000440d00004c00000c3000040300000501004c011000000000050000f14c00c00100340000000700000000c45d0000c4c0000400f100004000c00c0301000100001d0103004300c0000044043d030000030c340403010300000c050000000d000000070001070c0000070000c0311f00000cc00000c00000000000000030030004c400000700000c04300d100000000cc0000c1700004130030010044c000c000c040401040c10440f0c0d0c30c007c00340403c4c01000000340000000300000f0f04040001010c01000f530100001c00300c01c4010400040030010000000c000004c300000c00c0030000001000040000c000070c00040c0c0003000c00100f000c000c00000c003000030407003701010c350000000d0000000030044f04cd0000070d00000c000001130400000d3100f507330d0000130c0c003c004110075004000000000c003317000400140700000d0100c0000c00010040000f0c0c0d040c000000007c000000c401000f00000c4c070d401003000c0000000c31010c0010000c4000044010043100c10300000030004c000f0c3000000c040003000cc000001c0007040000c70304c10000f00400010000340003700004303710041003cc0000000f0100cc000d40100703001c000403004c0c00000000100101c10000c4010c1c04350004000004000000000000040000000f40140c310000011303c0000c410c0000400004001d1330010d000000c00c0c030400040d00000440;
rom_uints[124] = 8192'h3130000001333001f00c00000034310f000130c0030c4040003030030cc034000f3300000f303034000100031000301c70050cd750c010c3000d000310001440033017040010000c40003000500f131041030d40d00400c40103001301c700000c0d00014000040004001000031300000c40001000c1303000003043000c00010000f3113300000001000dc00000330000001000031c01331030001c004101d11000c000cccc313000003003000cf700031c10700dff004d04001003c400000300f0003d00007000101003000c00101033cf400730330c1003430110c307100010400400030000400030c040104030c030f13740400000100000004101300330030543440c0c000000000c4300000c00c10c300c0033030031003cfc1340cc100000000c0503000c300000c0c00011d0004331310031000c000000010401400440030c0001000000f3c00103010041003f0010010414030340d3d0003fcc0000041cc00fc0030100100c4000330370000010c04400307000003000000c000010301000074c40c007400003400000030000000004000010414c101400c0007033404010041100033001030c03003333033000000f001330000c0100f0c10000100001100071000d000050003100003001c01000000f13711000000010000c300c03003d00007dd01cc040f00030000310101c00000001000c0300103300300401103400313000000d30004cf030740c00c0007100011341004c3c00003010000c014000c040d001100f034c15f00004100030000100303000d0000c300000f71330100400000040c00000010001011d00fc0070010037103114040003d03301303f303300f000034101000300cc00000010cc33033103770c00013330000004cf00d0c0007400030d1034041003030004441101001100340000f0040c5c1ccd0dcc000300043c0c140000cc00c44003100310740000001003000445300d000d0340000003000000c0d00001000000f04014430c00030f37003031c1f00031c043d000100040001d00000000101030c073000001050701330003040003d310700d100031c5034007c00000000c00000003533c4034144dc0f104500000000140034300030000430030041033300030c3c040ccdf030fc00000314345003040c010c4300300d0000c00013c330d000700c5000400c004000014401030010c000c33703441400c000f3000000001000100410033cc0d0c00103004100110001c300110001005100443000030030000d00313000cc0000d03d005c0f00073130000c0c003100f3707400073c00130c0000c0c005c000100000f0000130000107030311c000c0300301c0c1000007401c00043000000001fc0001430000d30000400000c0404010001d00000c00010011000000000040c000c3f1070300531110000c;
rom_uints[125] = 8192'h450030040400000010100005f001001101000010000010000301f000030000100000111130d00000000030100030000530304300000400f00010100c70003000000310d0403004403000000010000000317300301cc05030000030300330000000311000300000c1004500113010031010003300030000300c40000013003000000030004c0000000030003010000101000100000000100330040300003001003300c0010000333013000010300000000001300000003030300000404010000c00f000300031030310000c001010c04c030030000310013c7c000033300000000010031303000003100003300100c00300c00000003000c00300000000103010000030003010c0c0c30715c30010000000f000300d01030301000030013010010050000030400000000030c11103c000c110040040c000000130050c00713050001004000013700fd0000000000010000130000331c040c0c401034000c0c130000c0133c001000010c0c00030110330300000003031100c010000000000c0030000f031c303000000703000300000003001403000001030f0301030111030001c00000100003010001030300100030330000030c0400000000000003070300013000003300000f0c0103031c030003c40001000303001000000000044104407030030d01f00000000040000400030003000301030013c0003000044f30001033000043103310000c0143004cc40003100003010300000c00000c0f1000300310034c0003f043000004340101040000303300000001000010c330303000300c301003030310001713001003000c300300033000000c0c00033101101300031400110001cd01000170000000010041000053431c00133401dc043f0013000010003000010c1c0033000000c40130050007000010000000c0005000003c0000013f0300104f010300030010300001000054030010000011030c000143000001001100000000000300131300001003134d415c00000000c10013030030003001001300000c0c01030c01130000300d001c4303001301000300c00c100000000300000000050d100c030000c0010000000300400c000000c000000100400c0103000f0000004330040310000400003330000100dc0000300c000f00c3150f000000000400000000030000350f3030003001030300030000c4c0d04303303000000131000001300000000000030040030405000003410133000003c10000001000031001107000000c000c0001c0f00330051000000000103000053005030300000001000000000301000010300c1c000000001d0000c4001f0000000c000c30d303001001431000040000000100001430300000000100100003100000431d03033010000100400f030000000300c000030330100000301000000107111c00000003;
rom_uints[126] = 8192'h3003000300001000c3d000c74040c000c0000c0c000004f001030004cc001004000c0400cc500000000004114c00c05f400000500cccf40040c340c000000000c031c010301cc030000d000c0007000000003c03c1303400340000fcf0000cc0304004000454040c0400d044000c0430007c0410000400000033300000ccc001c003cc34d00007100010001000000c0000400000000040300c300c10010004001c013000000c0054d0c0c000c0400c1040f0c00000003c3c0400010300000c000c5000000000010000000000ccc41400030034f033f0c070043c0400c04000000000013003c0000000000c00c04df0ccc00c4400c040040041040000000000ccc0000400c5404c01d030fcc0f00c70400c4c340cc00c0004010000d10001000c0d00c00c4000004c000cf004c00403000f40c0040040100100cc0030df005033f0f0004004d0d000c4000d0030404d3130c0c0400003f3404007003c000010c003000000f4c0f0f0030014500c0340100000000c05c000c010000000000300c03000cc00c00000400c000033000030c04000000400070c003c43d1c00f40400040105004f05000f0001cc00cf400c14c000343000c00c0c0f00000cc0c04c4400030d001c33010f000300000300000000c00c030300033001000005001f0c040c04f00000c000130000dc000f0c00031df0000d100f04c00cc4c0cc300f3c7030004c03f0100c0414030c400030cc10c0c370000c0303400c00050413070c000034c04cc030040c0c000cc00c00044000334000000c1340007d40cc0c00c04c00c004cc0500d4000c000c3000d00d0c0004000010c00040043044cf44030c31030000401c0000000040030000000000c000c3140d0cc0001000c00000003000c000d0004000000300304040f70c1c00400000011070034c003f000353040c000403000c354fc1c3303540c304cc0c533030c5710c00001cc400c43ccc0401000400cf404c0040400000c04100000c000c0dc0141340c3cf3c00000cc4cc004c40004c00c4c40000c0c000c4171004c70cc004700341000400007f0040001c000400cf0041fc047303c0040500000000400c04005140d00c00500c00000104cc031400000443cc0c0c4c000000c000cf00c370d4004f0c000c04000dc4c04f00033cc0440040c030040c0000c0044c300cf04c0c00444403300000000004300c0c0511003000000f0c300304ccc001000000003034000000043c004400030000010000c00000010704010c0340c3c043000000c03f0403004000c0040f00000c00000c0010004c001c0c40103001000100710100110004c0cc0403003004040007040f30000f00330d07c001c1000040f370001c00040340df0d0401040000cf04000c0c3330000cc00c0f00001000000300001c00040003003f034100000400;
rom_uints[127] = 8192'h140cc0010105101010cc007011000c100c0000030030330300303700c0073400000ccf40030cc101d0051c10c3000013407000c3030c3c0301000004110c1000cc000307c030001d1f0000000303110001300c103741c44304f0440c440c0c000700013000000cc000040704c0410c030400000c0f3c04000071100f010401000403340104d40000000000300000030c40c000000040000c04300c000004007f001cc000700c0c440c100c450fcd01c03c0330010000010c301000057504cc0cdc1c300400003c4c000c0000040000140413340c03d10070d003cf10001c0c00000d00c1c0c414cc00000010c11d4c0c000003134c74000047c30c40000000000c00004c140131541f0f040301c10000c01001c04c01030c044700c3440ccc530000c00013100030100c00301700ccd000c0cc3000000003000110700cc05410c400000000015000073c133dc010c0c300010000001000055700000310000c0c430040700300340007001000331410031c0c030105f001014000c33400400400cd00000fc71d7c00fc0c300c000dcc13c000000c1000c74c40fc00033130150c0c004435c3c1100d003034000503000c0104000c0c07000c30c0c4310011343c5f300305cd004001000fc0f077000c000503000c041307c30000cc000c000dc1030c00cd15330033c11103000040400f0000c0030001400f000c000c34f0001000c00314f30000c000c00f040700170c00cc34003c01300005d0730100000c0100100c0077cc00040000c0440000d001d134c0030051003103010440000003f40077c50f334374030000013cc003c030000150000c31c0031007100334000100034401100d430004100000400000043400440f11004d11c01c0c0303003705c003300070013003fc31001404c5c01000c0141303300400c40c340c003dff00003d0c3507c404d40c0437303c1300070f04040f050730c40c0040cf40000010340c0130cc000000030330f03000cf04c10007001c70cc1047c1000701400d000d0300040400c30c0c00401c0100c340337c03000431c01003c30100cc3300341c0d0040040001c0310100c01003100101030000040003300000c7013530041040ddfc000005c40c0004035c01400303001f00051c00003004010c0d150500470030011d70040001c3031c01310d57300c0301c0c040700001c043c1000c0000c0000004d044d30c000c3c0c0137000d0000001015001343003fc40403040044000c000f00c100c0303044c040000c000d03000103050dc000d404c1010500400503dd0003cf1cc734003dc0300000003c000ff0100400c00000300400c144000c000304340030310c331100000410000d00043010303f000000303004333000fc3370c00000c130013030000100c00000cd030cc4000077301405030000000000;
rom_uints[128] = 8192'h14000010040403300504300c0010fc050044c00130040000110430000c5c00104444cf100400100341100003043030040000f00c011cd000000000100000000003d00000000404100030100000001000300051300c3300000400d003c070000f30103000000010100c0300300000040c3003001c30303c04001043cc0400000000000030c000000000000334004034300030c0003010c010341000700000c4003c0000030033d004000c0c0004cc0300300000001003400000000c3c030c000000001400000451000400403000000c0030001034030004300000001c0400c030030050004cc40000003010004140c03431cf03c0400000000c0014000000c400010110300430001c4010000040041100dc300c337035105c0c00cc3c1000f03000c00000c0304300041044301004300030071000000c00103c000000030310300c3dc43000d5303d100000030100005cc011340cc400740c1df411150000300404000130c57300300f140010300400300cf000005c040c040004000000010c0c300410040c0c44400f0000330040d0f000040030040000100500c03040040134430050030c001410c3000040033000000004131000040550700ccc05d03c00c0fccc000cc403030cc3c0500000540c10340c0c7c001003003300000340033f14000140400010c43000c00000334d00cc001c0504000000000000003c404010c0000310004c30300004301c1004c00c00000c44140c0c000c40003004110047c0401c3704300100300c1030c300003c0000000000144c0030300414000000340cd3400010141c0400c0103c015030c0303004300404000000f500013014d0c1004400003c00000c3c0000cc0cc0d0000010f310110034043311c400733040c005c1000400000030004000304014100000003000000400c410c303000000c01001335c4c001430000030f47c34c1041000311404004c00c40c0401100330040000100000000010000030000c00001010001440c3000034005000c03300410c10300000300c00000f000c0000004f007000000150000400000400c0d03010410011303300300003041000000700100010033000300010004010cc0cc034f00500401004031010c0000030700000010c30001070300c00300034010c040000030c1c0014000310c00004300c00144c1000000c301000c400c007cc0000000010144400005430c0004cc00000440c0031000041d35000cc30103300003001030f003400d011000000007700305400c000c40710cc00100c000010003040c0c04030011030043100000101440003300c000c003310c0100040005000300004150c003003044c007c030000004000c40c000000c00000000f0000041014040c00004c000000001103000c000411030010000000c0000031000c003c00000000300000;
rom_uints[129] = 8192'h1173cc00500c0040c30c1000300030000c0000c03000c0300101500000000050003103004c3c00c0030000300c303030501304110000f00cc00000005400003001000000001000010400400003000c00000010c0c0007004000c440c3000c0100c53c0003000c0c101c07000303430f0300100114c104000000f0030103014013000c3030030000030c04000d3000c034033300000000130543000000cc34030c004100000104341000000400030401000304000000cc0000040000040f000c00c01000c0000c0cf00c00c0030c00340410470140040300001040001d1300000f10030c0c01d0c030000001f1cf00c100003c03370f3c01c3300004000000000c3003140013c144030fc5400141000c00001100100043310030c00c00c3000407370c0000000004004000cd050000c004033f00044000000000040301030000430000034c00043000cc0003014003000d10040c0040000103dd0030000000d0000100cc1000000000c0c00044c430030043414f04c0c000040700d43000144000000c030071000000dc0000000c0ccc73001000030007400044ccc0000000c4070013410304000d7c0350033404100c00c00c41000c0344000c03c340cd31000c00000c000c0001dc0c300103c000d10413f03c10c3000730030003000c004f04310d3005500d03073010000c00000001c000104d3f0000cc00030404c00c140510000c4c0c000cc403030103c03110000000000301100300000300c00c0000000000d140077043000000140431000d0c0731500c0030c0000011c0000400000000401d4700c14c04000300010f0000130c014c0401c0c0000c140c3c40003c0304001c3c00c000007004000c000001030c0310c10c13000f1113400004070c0001cc00010d000c0000370c01000040010c00030cdc0001d00000000c3cd0100d140001010303070110000c00c00400c404c00ccc03000f3fc30f004400000347000300c000000000000c04400301000cc430f04c0c3c037030300003000cc0100000c000330d1c000113c100000c0c040d00c0000040000100c00000314410c30113000700000c3d00000104000000fc400301010000000007f4001303000705c4f0000d14c03004f0010040400000400000003041f00404c70ccc003301000000000f0300030c33c00d300c04000404000004010000333c133c0000301c0003070105c7001000cc7000d14030350f000030714000030c10104003051700f001cc030c03000fc30000400d00030c04300c40711d00003c0500500c000c1000c57000000000003001c10003c74700040000c10101130030000410c00cd0031401000d340f043500000c1100000000010000010700010040000d0c04d3cd03040400c40c030d000030000100011100000c304000c000100110d007c0100300030;
rom_uints[130] = 8192'hc0000000c004d0c0000300000c00044c030c00000003c0f000f04c00f10040100cd00054c000c00c07c000030000030fc04fc1010c40134c103003403d074c000d00cf0c4000c0c50400040c33c4000cc10400004000dc4300d044030004cc0c0f30400403014000000343000f10c0cf440007040303c000cc740cc10cdc130043000c104c00000f0700404000000c04040000000000040c00300004401dc00000007400000c7100010f03005d000f10030c04c00003000d0310404043035000040000000100153001cc00004304433f0003c30000703d00c5000013f3000c00400400c00040400000700300c11070040c004003cccf04000c0000c4100000c0000300c0043010001003c0cf00010f01000f03000c740300000c0010710403000c414000c340005001001c400f0c1303000c0010010343000100c40017100f01cdc0070113c01c034003000344007410000034c03c1cc1c103c304030034c00c030c040010100c7c0c0d10c1003011000414030040c100000040001c4d0c001004001c000130c00110000001400100f00000010000000000c10000cc0000000000400001c1c1400300010ccc00d4400c040000400c00cf0004000000013003c314cf30000010000001dc04103104c000045000003000044401001040c04000000070c10c00c044300301730ccc0304cd1f000330404c00040cc3f30000c104c300c0000c130000000f05005c0f010cc00313c3c0cc114440404004c4400cd3010000400000f00000003c0c00000003000040fc044070431400045c00f00300100400001cc00040000041cc43000c4004000504000400cc03000c00030c037031100304074470000c4000c033030030004003f00134000003001000004007000c50000000441c04cc410cd01010d1c0030300130113c030d0000000104001c00cd030c00001cc000403004d410030400c0c0fd31000c0c00c000133c0040404003700000c00000c0053cc00000000000c000c77000401400f10c00334040030000c0000444c0300100010ccc04c4000000c0010410000000043003444010000000c0000000c401000f00103d0000300000000c0000c0003000003000000000343030cc00f400310410304050000000300c0c0404c00434c0c0300040000051410cc0440d7400c000c00c04f00000cdf000f44c0104003d0000d00c000003000cc300c00001311000c040000000c0000314030c0f000010301c4440001c1140000cc00000d0000dd0000030004040f0cc407c0044c05040d00030101000d4000044000c00c0300000c0000000000300c7000430c0cf0000000c0033000004004000c030c034c4cc5140c000300c400000004000000000450c0c007000d0034c0000000c00004000300d00000100dcc0c000000001c010043370c00700003005400;
rom_uints[131] = 8192'h4c434000c300000f004c0400011000700000031004ccc70041f43410330d004c0310100400070004000300043010030000dc00130040330304104033010303101000343000c0cc04000004705004c01003d000110f0c000c044004010c04c0300c100403000d0030cf30c00035140000400000f000c10000000000000007004c3000d00003100010000030040f10303000000000000404000000040001000000030734001001470000310000d0310c001030703000000103cc0010400c31004030d00043000104000047411300033040001034010030030400040110cc700000100004003000313000001c410340000c000104400c17003c403007010034000c0100000c4000003000f0030500c40004c04c3030cc040110cc7c0000c0c0303f0300000004400cc0040030d000003c100000300310001000000030074c1c100030000304300004403d1000f0173c00c140cc0003040001c50010d0f104170004311f0000010000304000c00003303504010000000000f3c0f100f40310000013405100c004045000300000000400301f0c0000c00000c40000000c0001003500004cc3c0041c000000400d0030300000000003c03431c10011003000040c4c40005c500c0c00303000cc10c003003110730413014301f030010c0305c00100dcc001030100050c00c30c41000c300004f3000d0400100333000000010f30c733c000c0c11330c3000040000c047533110003c0043000c700c004000cc440300040400c00f00010430010c1300010010000d0000000c0033010431c00000001c300f00400040c4010d3000f01131400000cc0300040000c40c01000401001c4010700003cf700300d0000c0141fc00c40110040400cf03500000c0000c0c430434040cc30410c0000344331000f0c40c40f50103004303071000d00105c301c04c07c00000004f0043003d4040401000400030c000000000443003304004340300000000d000001001000101000f4004003300400007000d43010300100300cf0c4003f0000050100310030134001d4011300501000050000d0000c00c40070004c130000001300d510000100000c300c1000400041003404334000001400000031cd0000000405100044040403c40c300000c000040c330c000300430040000c031c0000000000004040c100000c0000140330340000040007000c00054030000100004040c4000113c000000100100440c00010400013c4c050001300000000535353c050003300c00150340000403cf30300100350000001c40700503c14400000031c010c41304013037004000004000c00510f00c0030300f4003044f10000001013001c000000c0410d0c4000f00000000004c0100035c40300000030f00000f00304100400c00c000c0440310003100040040030004000c33010000000;
rom_uints[132] = 8192'hd000000005000030d100000000cc000000000c000000c1000400000100400705000f030000300000c00000001cc4004100cc0001000000000000040000404c0400000000000030c304000400000c0fc000c04000c3c0c14100c00d4d00050f0000000100c0040000c0003000400100473000410000000001c003c000c007c001000c000300000000000040000c0000030004cc000000000004040000c00d400000c0014040000300c00001000000cd0300c3c04c00000000000401001c0d00000000100c030c0003303000030007c303000d4c0cc00004000000000004000040c00000000004c00c0c30c00000c304000000000004000000000000000005011000000c0043cc010c0400c000014c00c5c000c3300000f0003ccc100004d00100ccc04d0c0d00000300010000000300505000c10010c003c30f004000410311cc300000000400000c01000500440000000300300c4d03c5000cc0000000000004c0400c34004d400103f3000100000000050010000005000c000103413fc0000304140c004c0c0000000140c0c00000c00000c030d01000010c000000cc000040004c0000000000ccc130010000c5034f014000000000304000044100040f0c0040000344004000000c00000c0000000010005400000c0d01404000c0014000c40000004c010001c040000003000c00004000000300000c001000000c0cc0010430440300000010001041300140cc0c000300004400004401f70000c00000000c403103000001053030000c000030c3000070040303d000000040c701400000050004c04c0c00000c000cc40000c000003fc10000004f400c000003c400000000000000c005c30000000004000004c00000c00304c003c0000d040000004000000400000000000000000000307cc03103040400c0003300000501c000400c00004d00c003c0070c0100410050050f0030000c000400000c0c0000c0000d0040440c0040000300000400c10000004000000343c0c0cc000000000305410f0000c00000c00000c0000303000001000100cd0010040030010040004043000007300c0f0103000300f01101c0001370410300000003000070004c04c0000c0d0000004d40000300c00001000001000003000d0010c000c00c00430000000000f0130300000000014501000000400000c0c00c0000000044130304000004000000000030c00003f3c0000c4cc000400001cc010000000401000004000cc00c0f44cd30004000c00000004c00000f000300340050c10d000300c0000000000000030c0000c05dc047000000c700000d00050100300011000000110004000c00030d050c00010c0f0c04000100000000000000000000004100410300000000000000400343000004000000c304400004c0000000101c014c010404f300000000;
rom_uints[133] = 8192'h31d0000040f04000fc040000103004c0c000300043cc00000c70001505103040104010000c400c0003f00070dc0070000c0000d0100050000030000710014000c00000f00000c37000040c0010040c4310c0cf3c40c070014343c4c030100c0005c0501000c000304040003003c0103104fcc33007d04304073007000030000133c014104000000000c00310c30000f0cc0040000040c01301000310c0440303040700000400100004c000c0703014004140d0000c44c030705414c03c700050c0f000040000503300f030c03c0c300c1c4040cc000100c040470c100000030010300c0003f0001c31f1c0f0cc70c010c17100004000000000c0001000400034104040034000f0c000000300c4340430c04300000c01c01c0014fc3000001cf041000004100c00300c3000c1100f0001c1003040f430000000003000c0dc000004c000c000cf00033000c3104000c0c0011000010010d000301c5000050f3330005050c040410500c0000cc0014030300003f300504c000c0c1c7c01f1000f00d000400c14000c0300c00c00d0c40c400001c0000000004030100500f034000033f03c0000c000101cc11044070000000d0304c0003000301000c0c0100700c040c0c0000040000003f0400c3000300c031030c0030140d0030030c0c34c30c43000740d4770003050003100c03401c30000100030011f0cc000004037000030300cd510c0000004c10000f010144010104c403300c3301040f031f040c030c3f4c000c30400d0000010c0c010100000c0104000000cd0010030100100000f00c001f050c000d0100001100c0070c001c0004334c00070401c0000000000013000300341f03000000c040000100c000c004d000000043c01c0c31004f04300104400300400403000cf1040000307c17300530000cc0000000c0040c0440c10c0c0c0c070d00d040030f014c00310c3f040cc400030000c0000000340c000003070400000000000001100104000300010040c40000033f44c00c04cc0107100300000400040100010400c01f0d0000c00404000d01c0000000400c014f4335000000000c4c0050cd4c0c03000c300c044c4d00004f000333f10040c3310c4000700000004044d01340001c501000410000000300007030000c0000ccc300110014cd00000434c000000c4c0004003000150343400c000c0003010400000c0000300040cc03f40430014003034030000f0c040d0c00100100000000010c4d5030cf000100010cf40d0c04104700003c000005000401000000c4c047c04104030f0000400043040100370c044c0000004c00574000c004050c000040000c033f100040414030415c310030014c33330000100404001003000000c00c0000000c0000330f00343d0003000304010044030c300000030ccc103c0034000007440c04;
rom_uints[134] = 8192'hc00010c000710410100003000000c0000d50000030000c300c000c0c004c00000000010300f4c1c00000c00000004310fc3334730ccc5447000c3010c00000000c0000000001c400030000ccc004c3d0c100301d04043c300c0000c00103c044f0035000410033c0c0000000c10050cc400c043034304041000010400044c000010cf30030c0000030c0000000000470000000000000d04110500300fc1c40100c003100030f013400c3400030c000c3d040100000c00010317010000330004000c40c501000403000400003330011cc000c0000401340c0030cc00cc0c000400f74400030f00000000f0015fc30f104000140c3c044000003000004c0000000c1330d0430011101000c0cc13f00c1303015f0100030000000440011d41000000000100074410003c300300d4c1035c030c0000000410401003fd3003003103f5000c3000031304003034110130c300010cc0030401400c1c14c307300c0c100c000304000030c03000410107000000003100030c0000000c0300000c330110434030400f30000c0c1004000cc041d3440000030c0000f0d000000044010304444c00d00c0c0c0101c0d10100c07cf0001010cfc00d010400000c300f0fc3111000100f10050c000001040004000d400003030c4c310040c30c00000000000440700c0300c03d01000c30d0103010000c7000100110030000c4c010000100cc135000c0c4014001000c01001000003030044000c00c0140040017434104ccd010000040011cc0000001cf3c4500c103000700300000c003000004000000000000f1131c4400314100074f01000401130000100000cf10340dccd50501030400333cd0054700000d0000001400000040cf00400c300f00300c00414000030400c007cc00c0c00004c0003310c33c00003100c1340000073010004300010717300c1000017c0033c430d010cc01100010000000c000000c1d1c4c000010030030000c030cc000000300d0000000034c0c04104f0013330c000110043fc0031f033d000010001f000010014000000c000c143000040410444034004c04300331140310001017d100003ff000c001c50c0451100c003001001000000c001030001c1cc00000003743050105500404010c00000301170c00030300d401531000004005033015100004000003ccc4c013034c07000000000104410c0500300014100f00004c00070000000400c30001400fd11300103f0003003050c330010c0c0df0000014000030044000103000001004400000400114054c330103c1fc1cf04000010ccdc10c700030d100000010010cc000000c343110000d00010cc000cc40001000f137000c300701000004000f0300014c0000000c10010300000f01070c13040d03011301401001001400040c03030001700303001303c0073000040000000;
rom_uints[135] = 8192'hcc0003000454c000f0300130100000300301100cc0c01330f3300d0004cd040303400070040000dc00f00cc07c3000fc00c1130c33c40043d00400044000c4c340004445001c00130c004c0c40d07040000454033330cf004000000400f01110001033c000003f0300034c00030d04303000000000f10c1004f33000000730f07030f0011c0000c040000000300010400000000000007070c40305000000003110300050000010c045340000c4300c0c0010c41300330c13c00000d000700033400c001041c0000000000c0c000c43000ccc00000000440cc034c1c4c14400c0c0000040c0130130300540130003f030c0344c000110000000040000f0000000c0c00031100cdc1030001000114000100403c000c1d0c04cc07c00300c00400f400430000134001340ccc001f0f070c000d0330300400c00c00014f053003010104007000c014030103c000301000d0c037000c0070d0dd033c03d0710540330c03000001430530401701100000004313030040000003000100003c3403007c0c1003330110004d15cc0000304c033000c0010300000c4041400300130c010000300c40040c0047d301040d0011cc0f04000c04400040100000040300f01cd00000043c0c0300c43303400000c0003d0f000000010c0500000cc3000030cc040c0000c00d0407031c03c033c003c0044f00000530003300000400000d0040303ccc00cc4400001000043033100004c01000dd00430004000040c500004c00311101003000d00400000c0004c70c50000150cc40040000c00010400c000c0c40050c4d03004300ccc00743c04330c05300030140000d00000c1c0300001c0000003110401c300c04cc07fc40040f040030c003101447047f04030c4000000007f0400c03c300f3300010010001c0c4000031110f03000000c4030000000703d0300f30340d0001c700030f1103c001004000104c000cf03f07c00770000000000000003000000c00030033c300000030040c5003004100001400030337050340000007010730c700000004000404c50d003001410040c0100301300001dc40c00c0043010034d00dc0400301c00000c00410041c01030430014004030c14c004013040000c3040000001040100000300001c0cc0c40c0c0001100000fd0d00c00003cf3000c0000c4030c1000c010c000030000000c0000300c003c00000330cfdf00c10f0c30001c310440d00000000c00100010d0d0c0310c500001c0014c504cc000003000000c000040440070c040401000034031050010c404d001f0004f3403c00157000103c000cc0000004c00004000304000c1000000d00004000000300c01c100c4c00033c00c000c00000700c3c050404000cd4300c03301040040f0c300f014000000c00004040010f0000000004310000004700c30ff10c03000;
rom_uints[136] = 8192'h10004000c0f01070c010c100d10040007d00001003fc0300000100c05000000404000c3014d50000000000300000000030d1073df010504000300000330000303000cc3400c000d0c000c0c40300000401003000400000000041c00c00001400000000c000004030000000003000c0c0304004704300c010c070000050400000034cc10004010040000000000040c0000004000c0000c1000000104000001100400c3000f0500001000011004300f010000000000030443040043033400000001c013070d1000000300000d40000003003100100c4f030130050000000c0000040000000000f0100303000c30010c00c00003043f00000704c7000034c100044c300300437703500000330141030403c30ff00004000000030c000c03300000000cc4c001c4000000100000000040000000010c030005c00004000c0c1100000c03c3331003c0040c0cc70d0030001c03cc0000000110000000045441c3c00403000c0001401301c40c001000133000300004300000000100c3c57000000405cc000044004004000c04030003300031000000c000040030000410010000c00104307000000303015003c00d4c000c0c0400000001100004010000000034001300000300010000030000000000000041c004000100000007c0000047430c0007411c00044004c044c31033000000030c0110000000c4d400100000000000070c0c00000011c00110001c0304011101010101000400400000003000c410343c30010000000001c000300000300344010000c05300040c0c01000334100300000040c500050001000004c4c0030c0c04000007c030000cc1400c0c7340075044070d411004000040000c0300c1000f10430034030000400031000000410c003c00400000003005700000c0010d7d5d40311333404004000c3100000000051300000c340f000011440005c4005c00430004c000c140400c000004000f010000c000043f0f000000000004000c00030504004401d0040300c40d010c000f030cf030c010000c3d3c0000030d0004000300003c044030040d00100000000401100c3000000300000513100133040003000000040010c0c0440000000d070004030003cc00310000000c0000010f00100d000130300000000400000000000f400c04040004000044440d01004d001400403150000000007000c0003004cc00000000014034000030000001014000003000000000000040c0133000030c00000101000003cc00100f00000000010000c000044400c40010000400100c730000001000c4c0c0c30404000c440000000300000d10c00401003300000400000c100400400000000c441004000404000000d003010000000110030004013041000c000440000110300003cd100000100000070100030d04000c001300033374000c400100040;
rom_uints[137] = 8192'h101000050cc4000010000c030003300c000004cc30300400003c3d4004004000000000c4c500040c0300004c100c0003d100c030c00140f4010003000c0000100c0d1400c0000c0000000350c0031c00300540034300001550000000c01403000cc0000300001300cfc003cf00041c0001040f10c000030c141cc04030c0005cccc40c300730c00040c03110300000000000000000040004040400d44c3cd000304f40001d0107040c00040d0f030450d3101000100001100000000330000033f000c300100441001400300000043000030c0000300330c0f110cc101d0000c0003030000430000010007771007c0030150400071d0000100000001300000c030100343070c00410c501c001c00000c0400737cf010000cc400dc704040c340c010c00340030040030400004c0000c34030000c000d30300030500f0001100300c100000030400001000cfc340c0405c300010001100c00304cd300000301c104d0400cd0033c441000004754130c000033c0000410c00c00f00011414d400301033000110100430700300f1c011f400000040000030cc0d101003cdc0340001011001040401f00000000c0d0d410c00000cf00c0c13000440c0004000733c004d40031000000f00fc000033101c00000103c710c7f30033f300c00c0c00030001537c01d0001c0d0300004f0410041cc014030c4c00003c1c101c00dcc403050f0310010031010c3303001c000cc3cc1400d0c403d3c00403330c110033044c0c003100cfc0d030040c400101040031d0010000304000003100000c0014000310001c031040c0300000041c400f00043c10013c001c0030cc0410000c00103105000130100010cc0333010f001030c7040041000f0040f000300c30003010104130004010100030100c0c4cf30dc0000cf1070fc0344c0000c70050140730400f0000c030cf00ccc3f0340030310100010c0f33300c001300400303040030c303000401000034d0100000000c0410001010cc043070c0030014c3000000c3c0000700440c00000030c440455004044c000d340034c4000000000010dc40000400000430c300f0510030000004300fc430000000004000000c0400013010000c1d000c750004040c4c4504c04400343000c03430007000310103f330070000000010000c100c001c000c000000c00001330c01300031001000c0000000040fc711007c303100040400303104c00c030014000004003c00d00d00f001130400400001101c004c04c0140000051d000c0000c00f000131000dc40c340134c07c013c03cd000c040301100c400c004df30003004d40000c00000c34000c3337004c0311100cc10000003c00000f0c0030d100300000f000cf0c01403000000fc40d00c410000017c00104c001004d03003f0c105030040f3007140133c00c0003;
rom_uints[138] = 8192'h35100000c00000400300101c4f40f400c33400133d00d04c0c040303f00000000013300dcc000033cc1000403c003000d03401340cd34000004400c07c1070303c3cc000303000f0330033c00100ff1400100c1014c001445031503c00003001f030c0d0c030303000c0c340c0541c0c505500f00c1c404000003c307410300000300451c0c00010003400500030103000c00c000030043c0dc0dd003c10103003100100000040f010c0300001c00000703c0c000014044c300400413c140000c0340cdf3000d00c00000000d0100030c00504c000f1c0000015001004750c0c004000f030c004005050500c01c0f000000043103034000000c300000c000000fc0ccc0410003034ff00040c710c00400cc4f0cc0003033030040c0354d1f0cc1030c00000c000c07000700c4030001413c33c000c30440000c03000c3300030c03c0014300c3100d0400040000c003110c0400010343014d77504c0c0033000005431044013003f4100c7000cf01c100004ccc0140dc0010330d0100000d44010541000300000300c1000c0003c0c043c00300c0000113030c040010c300010301000003c3c0004007cc3000400353010301c0cf01173c000001c004071340cf04c000010c000fc001cc300dc000005141300300000170c00c00df030043440303400fc00030044000cd0c0300c033c003c30031300000300000030000d10c03000f0000000040c7c00f0100030134000001010cf100013003c1f0000d003700000c0041000000030443c303011100030341c0010c340104040100c04103000cc1c700030004000dc003010303c0c04000003c01c3033004c4c30105130c0041000c010f4c0000030100c3100f411c034305004f0fc30003cd030000c004303104040cc0003cc004c10f40000c330071d544030c3df04030c000000030c34003c1c001cf41000c0c4cc5030100003100400f0d3143c0c50030000100cc310c1df10cc4004003110430035000000f300cc7c1c000c000344cc400030000c1ccc10000000c0400c0330003050104004300c001c34c0c013001700f0c000003130301000501c040040340000000c03000c03030c004c1000d43054003070000074343d00335100701000c00100c0000040003010d00013c03004d000f0341cf0000000c00000003c1030f014000030000003dc00dc0c3100001000040000300ff3300c40000c0000000400005001c000c000040474000404407c040000003540cc703040000c000f33cc301000440040003c3507d0d04431c0000571004134000004303c00c00004f010c03040040c040010d370307d00000300cc7700f010f400d013040400003c00000003301430000c301300000c00000100d000030004300c0000c00cc030000304c0000cd004f000cc040400c0300c3c330034300004c000;
rom_uints[139] = 8192'h740400c0c100010000f0004500017310c140000000040c00d10300700043003000000043c000004000000000000050c0c500f400c004c0001000000c00040400000007000000370000300004003000300000104030130c00c000000030dc00001c31f0003034030004100000c03cc040501404100c400310f03300c33100000030d000000000100450000c00004dc0400400000013000013cc0000c0140d140001000000031001000000001030000310000f00000007000030001c1c0100301000000400003040000000f00100105000000c3000330d00044000c000c00000303000c0c0000000004400c3004000300040010330101000000000300c300030c03000303330c40040cc001c07100000dc510000c0000004f37000c10c0300c030cc300005d000c0c00430003070530001c0000cc03000000000000c00c04c00100c03c0000cc0001003011040000000500004100137001f1030d7143000000010040c1000740c3003000004003000000000c3300c400000100104400000000400c00401d70100101f0010003f300400040010000000c0000000044100300400c03710003000000000c001c0003410000003004cc01110001000403000331410f00c100070004050f00000000d0000300c0001010030410000030000c04000c0c030000704003017303000dcf0404000c00040000000000407000c0000130cc0c00333f00054c0300000003410f000401000000007001000301005c5000000330410000010c0005c0010100001000c00fcf10010301050f0c0c304301d003104031c030000004000003c001fcc01040300000030000300341c00000010c0333101033033c140000000f001c0001040000c03304c003000340c0c00001c4000f40c00100030c4000c00000000000000004000044100003040000000004033f5000000040000001000d1c030c000c0004003000034000007500c0030300030000000400c03c000000330300004000307c000001340f00030c0d00c703c0c00304c04000010f40010003000005c4c1c00004010375c00073400c00010c0004040010000000000c004003330030000710000700c0000304f0410d0400c0000040010f0c000000070010000c000f0000370001000001010130c0003c00000c01f307000f43100040c001000300010c10c34000c070000000d300c14100100000c3010cc00400c04340010040000004003c000c00034ccd010004010100030000311005c000530303070004030300c0401c1330015c41130000c00f400f0031331407000301c0301004003400000400040031f000000701c003000300000003041040c300030c0c0f0303c0000cff104c0000000001000001400c30003000040000130300000004030003010103000103070140000015000100cdf50000cc500000400;
rom_uints[140] = 8192'hc313000d0f000c000047c0301400033dc00303000c040c0003004400000430430040500cf0130001034fc03f03000c03d11000004030d0130dc0001001000c040533033c000c0c00c000030c000000404100001013004c0000000fd00400000000403f0007003c5d7c73400c4c4044d330413033000730300411004f3cc400330350010000c0c07110c013000000dd050000000c0000300003040701c10d540001134010010c3000400001004030300c0c340410000c000001000040c04000030000c40d00001f171001004c1c03103d03103000f70350d00c0c4d4000030030300300400000400f00000303100000c00010000c03c00000cc300500c00000300003430303003100300030100d40c0000001400001001400c40030f0cd10100043d0f0001033c03001000c0dc73430000104000000010f00cc10c0000c00000074047c030000c0c0d330307300c3f14010070300134c43054c304c3010013000000304dc34005000001100f015330dc30040100113c00000010c700030010100c3010000cfc10001300000030100401004000cc00101304000d00c0034001000014c41cc400440cd07f11710044000f003000007c4300710c10040c3003ccc453300000c00c700034c740000700000043000c0c00d04030003000000040341f500f0000301100c0c001003f0103c001010d10711c0f0103000030000017c413c300040c3004140071310140013100f05000005000c104040014d511d4d30101d000cc0410304010f03007003170004000000000c000c00cc070d00000700c043f00011000033000311c000000000c300100301400301030105330303400403c0100105044033001000c07300340c0300c01f0001c01000430000c4341003110cc0c001c0404301c4000c01431c30f3400c0470fc001f001f0010030001330000c044000f3c0010330c3c0dcc4c3301c0430400430000734c011c030300c10000cc10133101000100503007000c000c0007100000100100043300c704030010c071004000010300100050004040430001170000100340ccc41001000031c00001017d000c040130040040043000004000000400c0c00300000003400030700011c4c00000031004400000130103003000005400001c00c0000c44003f0100003000000040330104013300cd1300034c00073d00c7100400504d140c00c03553000000103c007c001043004004c000000010c001d100001c05c10c007c0c0100c0017000c0030040000f101300010003054c034013500100010c300d0111030c03f1c1f3300000300c03000300000004c0000000f0f400000000700100000010000d003301000c14500001000040400030030c10030040105c40000010300400001110000400c0001311c4040000c30cc0070000300040c3000c13104000000400;
rom_uints[141] = 8192'h100100000c310040000004440041c040c000000000c0f00000c30701c0030c70014141c110c003c0044c0000d00140003cc00001f0c4c0cc0c003003400000004000003400cc0000300000c0c0030c430c01400c0300404f03404050000d0cc000f500c00000c00c4c00400000440703404c001c100003303011c003c0051000c0403000311c0070c0000000110400c44303000000000030cf00f00c04010040430004000140304004034000000cc0dc01100040001c3d4000100040000000cccc010000300000d0c17000d0100043c00010c0000c10d4000110501113040300c00500c0100c100000000003000000d103000c400cc00000000c0000100000400cc14000c0c00d0000400450410000c01770cccc04f3cc00c040400c30c00100c050c400c0fc0000001400000040001c00c000c35400000301c04030071040500000f03001010000c00400c00430314000c000000040703c4000030000404040d0000040c0c10000000c303001c000000050d001c00034000301d000100040000000d00c330c103000c000c00010401005004101000000c000034c40c1c00000014c000000c0000000000400c0000000fcc10c0c1030003300010001000003300310303150c0000c000000410300c000cf0040003d00c10000103000000010cc1000330c40734000c01d00c0000340000cc000000000000043cc01c003400030000000330100000000c000000311c0004000004300c113030c00c04d000cc00000000c000010000d00405dc03100f30000010000003000c000cc00030300d0c0d040c051000000003cc1c0c0c00040c00400c000c0000c000103400c0c10f00003400000c0400000c00004010000000100c0011c00c14300010cc00040c0c000c0014dc0c00c40040000c14144001100000c400000d0c4c000010400450001001100cc030000c0c003000101c1c14040c0000400000cc0304c00c03c10c0040040c0040000000043d103004000001000c300000000001000fc4000000001c1504c00c0c00c00c010000c0001f03000400040404131000000000000c03c5001000d0030000000111100000000000000007410d0100400003011000000f4c0cc001d1001cf4000001c00c4c00cc0c0000cc0103f3000c1070000000000cc3c004000f000004c00c10000000cc47040000041003004000400004fc00000c700c0c0300000000000000c00000cc0030000700000010001030400434d00000003000300334000c100000000c0c003c30110310141000004510300300000000c1000c44300c35014034c0000000004300001330040404504000c0003000c000014ccc0004000410044c0ccc05000c4cc40c0c00c04000000d001c00000c0000c00000014000000c00000cc0000cf0000000001c0500340000c010001d0000000100100;
rom_uints[142] = 8192'h304000c4c0101c400400040000004fc04c000070c5c040000cc000001000c441f033dc0c000c00304000c040404000c170fcc00c30040c00cc0c44c00040040004040000000000000400343004043c4cd4d03c0033005000c7000003cd0c0000100c0040000000c007d000004dc0400c0c43000000003003000f44c00040c17c70c000c4100100000cccc0000000401070c300007410c000003c40303110c0c0c0000c000001d000001c100070c0400440c000000044400c00000400000030011000040000000010c00040500400000000100000cc0cc003cc0c0dc440300c07c0c40c040000c4040000c4c013000c004010404100040000040c000c000c107000001000dc0c000070041004c070c00400c000300030003470004c4400cc4004304000d01cc430c000313000000cc00c0000c0c00c1000c000c3c03c00c40130300ccc4414c000c4000000000c003001c03000440c0ccc100c01000750000030030030c00000000114c030c040c0400003000c01300000c0004cc4c014c14c00003c0100c000000cd0003cc4f1750000004000740c00400104c430000dc034000c00c00c100f0003050c000000073400003404310400003c10001004c0c00433c3cc00000334d04034000c0000000330cc001d10100c4000000003100c030000303000303000000130344c0c00c43470c00400403003003430000d400000cd00cc40c100000000100c3314cc04400c0040c40000c4013450c40c4030000cdccc10000cc0cc040000d030040c0000d507d0700000c0003000d400303040f100c040c00000001000c4003c4070307000cc003c000cc30000d1f0d0c00004000140c0031c30c01000d4010040c0107c00c0000300000400005c4c4000d00003300c0c000cc030c030000cc03c007730410ccc00c07c40100400103001440fc0000c30c1c0c03010410040001000c0037030d14c040c0030300004740010703004003400000000cc00400403000003000434003f50c00004c00c0c0cd000000004c000300070010040f014301004101c043100cd100400c01000000004dcc00000000440c03010000000000c400c10c00c001000c0001401000400d0c00000040007000000c0d410004040c00000000004000000d0004c0c00000004fc0000101440c40040c00000000000c00f00d01c401c100f0c0400d000140c4004000c013004040c30cc0040000034c003c0000000140010c000330730c0000c30cc0030cc0c30003030000000000004f000c007044100c0010c50030000c03c000c400004003c0c400c00c00c00c030c0010c000004000000000c7000f00d00000070cc0c0c1000030c400000000f040303d303c04c00040004c04030000000c001000040303c000c3c400c70d0443000000c101c30403030001000c40430f0c0704000c;
rom_uints[143] = 8192'hcf01f4000c0000000000c401f00000040500030040040037000fd04c003003100300340430030000000c3030000004503030410c0004d03c0c001104030110070000c4c701000410c400c4fc000cc410100300c0c1d000403c3d4401300c5300003c130c1f1c0c403f00c300001c00300400000c0041003c00d5000c00c000000004030000000000000c00711004cc0c00f04d40000014c070000004c4301c043c0010300c00010c001000000314c0030c000c0000c40c00001ff4413100000000c000c000001ff0000310100400047000c03fc40f104400504c03704c1000000400000400130c0000400400410000040001044c003f00040101050031000c00c400000050300c00004400c4d700000311145000010c00003cc3004d1041550001371400503f041404001030300c144d7000c30c00014d0010000d0c3d0c0004d004400d00040000c40300500f0010001000000100d7300c533f5d510304101c004c00cc0030040434d00431c043013c000c00003c3c001cc304100104c031000400c0330407010c07414c0441101c070000c0f0000040000c0c040000c0000004f0030f070010c003000000430c1010400300c0104d0401000030101c071c4ccf00000cf400001c01c430000c00c43c4c0501000c0c03300030000000044c010c030f0d0400300000cc0404cc3c0cf7000d00c70c000c0d04073000003f0010cc1c03cc00c44000c10434303000c0030c010c017c0004c03400c40f303d043cc03d04405c30050000071404304070304403cc4000c7c0303031c41150040040c00003c00c010000304400300034054d0110d0100010c4c00f14000f301c0c0001c3000000040cc010c00040100f040d100f3034000510c015000c0c004cccc400c3130300cd00f0c0001c101dcc0700000dc10cc0c00400000c4000c00000450dc40004c1010c4c0f0000100c5fc1040f3c00cd003000010000c73000300f30170004c40000303c000c0300004c301100f34000300010303c30c01040c0c4170000c003c4001000140c043030d40010c450f030000300010c0004103c0c00003040343004f0300000000010040df03cf340c500000400c000c00004000400331d10000050f30001304040000000040000c03003041d0000044d5cc00c0130007111000c347c1001101410000c0c0100303c0c0c10013030100c0d003010300104003014000c10003c4c030c00001c0001c300740000110010410001003cf0030c00f00400000c000c00f4c44c0000c4034c4341000003003c4c400c00000001310440c407001000c00cc33d4c30000c00c71000000001000040030001c04f00c0c000cc00000c0000c05000dc10003c0ccc00040447010007cc00fc000007040c30dc43500073c01c10fc4d40000c0c0000c00000030400040404c00000000d;
rom_uints[144] = 8192'h10103000000030d00000404040c040c0000c00c000000c0003407000c3330033c0c00030f100c00000000000307100000140c0404000043c40c000c3c00000001040c0300001000c400c01c00000c0f01c100f4dc0040c04500330c0c01dc000430340d0300440c00c3c0003c43c74040000000000f03c00100310435140430400c1c70057f000c0000000c0000003d014c040c00000ccc3fc41000dc3c040f300c440110101c00400000004101044400003000000c0103110c003074000000040f00303040050400c440000c04000000003c00c000c000704f0d30305f00010dc000000540c4040000010f00dfc401c04740071305000103000c10300000001c00443c7340c000d304440ff10c310703c00004104000030c00013cfc3404144370f30040f411000f41040037400d4f0d003f304f40003cc40d03040f0c0c4404003400000c300007130d031701000c3001001030cc0c01d00704430c301004000004000300f50003000cff050300f30001303101040c14001d400304044000c0010001140050d0cc0000003000040301000c0500000f00040c111000010400314f001404000c3c0ffc000005f030004000010c4c0fcc040c043004030d470dcc0100000400003113003c03c0000101350c0f00000f170004000c0c0c74051c5c00cd3035100f004c000001000c04c40f0430c04f0c0df40400300c07300ccc1404300404303f000cccc03f03450f0011c4000c000c1f10d30c0005000c0cc50730c330c3470c00030011100330f30000501c0000c034400c4f00000310004c440cc5104104c000300f00cf03047c30004dc00c0c0400153c0c0c050004070c1404c00c0515040c003110c1c10033040c00010f00000c51000041000000330c1f0131043c0000c0f3003f00001000040c3315040140003100000f001000050c050034400c15044400544f0400040cfc000fc0044404300030010c0c0001d00c0f00000400003c077c34000001c40d00000fd30434100d0c3c0530300c407d003c00003500cc3c000407043cc0001000001c0cf70040040300400c0004013001cd001c01313c000c300400100c430000c0440000000c01003003030c00013c710404013530005c300004043000c00c400c107c04030000003530030004030c0c0c00c0040000030c0104430031f01000303c000700400030000c04004c001100100103c7140d000404070000130071130040043c3c0df00cd30c003301310c71c10001000c000d040414005c4001c4350000003344000f003f0770000c00004c0f350c5c13140c4000000000c3000f03001310003c004000000035000c10040c000c010333041000003d000000c3003c00040000004c003c04300130cf470000440c100000cc1000000003000c3004310400c000000007040134003440c40000;
rom_uints[145] = 8192'h7103c10040040010d00c0410d000130c0013040c0014344d0c043100c301000000000c4c130f00cc3033000c0000d00f370040300c00340d04000013000000013400000c000400343000fc133010000301045105c0c17301030c3c00300d00013cc010073000100c400c0d340cd3100300000134000d00040001007030000300cc3cc500010000030100c003010010130001000c0000040c710033010013c00000140430330f00014c00040141310030c000300000c00017000030710000c030004300c00000cc0001c430100004c00330013c0040101033041c0040711f000034100c300c04d0fc004001f50437000005c5033c100000c001f01403c300010004130000300c07c01c00330044030000c0340c40100303335fcc014504733cd40c503000140d043000003c03cc0030300410300040003f30330300100f5130370000000c0f004130c00010cd33303340040d030010fc0000137031400003300004f10007cd013c310c000047d1000ccc0003f0050f050300c43000001c1040001313070100010c0030410030cc30c3110000100c0000710070f030d000440103043331303c00000400001d0700003c30300100300341c3300404fc3c0cc001151f040403001331ff00100c333c00010000f1c015c713000f000f004401fc40f00304003000c000030cc00c01000f33000003000cc00c073c003000000541507401f00013030131300f0dcc003fc0cd0001c0300700c4113c0003d00411040004017400770030400d000475001c47c40000c14303030000433040fc3c1000000cc003c40c00c071000401000c33c000000f04000034f0c0cc30740c0000350f43003400000303000031001114cc00000c3f11f0c03d034000f00410000d0c00f100350504fccc0004403d70004007041070330010c30c10c000c01100cc34303334030000301c0030014443f7000c00c40d4030f0d33c0c13fc003c400c04003c150c0d303000310303000030030f100300cc004d00003cc34d003100df00303700000104f1003f040401c01005cc13f010000d0c033c1400c0d00000330001000504c334070000003000000000000000370c0c000330103000f00c0c000d0c00303133c034010000cc010700000103140300410400f000300040c01405c0030c0000011c3313011c00c4f701043101003cc4000d05010141071010000f3730007000033c004100c030301000410004440034dd00300003340703003140530030c43300010000c000000100000000503c01400510c0003c000f4077143c1c00cc0004033511100c4c100400013000010000c3030070000c0303000c00f304100134c00001000f30f40004c0103c0401310f000000000300043c3000c1171000000f10c0500034010c30000000503103033110100c005000340300c30d00030100;
rom_uints[146] = 8192'hc0c0000300c0400c500c1001101000003000103003c30000000d004407333001010c00cd104030c401f34004cc330030c0c40500f004040130000407440440f004cc40c0005005111000c040400051050403c401000003000030031030301c000d301000c03c0033000c400431430010004430500430030010cc0c00300050c041c004001000000000100000c0c04dc00030000000331c00330040c1c33c1cc034070c00c000c31100130033705030000004c3c000043000004003c7d0c00c300550c0f00030300c3fc0001500001c300050f00c04c050c000430044005c00000c700050501c0000340000101344003dc00c0d4cc040040000300c00300000c0d403dc04c0c070cc0c53c01400400d040fd0030135c0c000c000f40c34c401710c0cc0001340000040c34050000000c004c000c00000400004071c01004c001017d301c000007000d050f0345004f07cd0100031d150003013c5040d3000d031000cf4101c400310c0c0400c00c100700701c03c0307c00d1df14cc0d1001001c00100001c14300cc4c4c30030041054c00100000100400c01000044c00c50400403003030c03d1001340000cc00c000c0000400404cd0c00000c0000047140000f030035030040000c000301004340431c1c00000d550cc0000003101d03000410303500c10f4000c00000130400000541001300040407000c0017cc0000001d40004dc100000c030f410c010310040407cc4004000100340400c00000010f40000003c7d400000004c400300005000cc040000c0cc340000300040c0000000c000f05430003000cf010cc10001300cc0000c0010304044400007c00000313d1c000000543c40c01d0400730c004cccf0500c43300c130000403000cc00f13c04c34dc4003030007fc04400d01d400410c00c010c1005c30000000470000033f444c0d03040c00055150c3004c00c3100c010c007343c4c30000300f03040001101f0c00000c30c03300c40c000701001100400c010005004f30d100300f000c00100c00040000c0050003c30d050c3001434c403005000400000003f34f01c0030c001c000013050303c500c033000c50000053c407000f01040c0003cc0c010400000c04000c0303010f0000033004c40300001f0f0c0f33000c03003700300fc100440030c00001c300000040030003070700330c0101040100037100110c0400004104003100040543c4034000c30c040c000414c04c03001013030303030c01000c00100013040c010401c01303300c414c0c0000c710300c0300c043c00330c704cc0c50000c004301040000001145010c000dc00003000013003500c0c0dc04030040d000000c100300330404100400700307c51014c3c103004101000300cf000c0400000c0c000404c50f4100040003007c4d0001004000070040;
rom_uints[147] = 8192'h30cc13300c0105c000030047430003030f10030c00c00d070000500c00100c0d010d0730c00300000c0130700000001001030173c00310c70100001c04300007300003c304c0030d0000000c03011011033f040d4c34c0010c300033033c1004003d0701f0c004333f30301003000003c01100c4c31f0c10000430c40404103313430100010000110c0303010000c10101033000003010000300300014c10d00011d0004c0044000300c00f0440040dc0104301000003000030c040c13000000043f003c00004c070140001001141f043c030cc701330f30070f0030031500400470000500300303031c0c300401031013000000c3330000400005c100c00000d70000c73c0c0514001000130000003000153103030cc00730330010c1cc0c000c07000003330015003104c433047031013c000c000c3100053c13030331c5d41003c000c00143000403c400010f3c00013f1003040403001003310c1053040003000c0400003f0400000300000300c303030c01000000c31c040c034405033340501104c4131013050c0c053100044340004304c000000000dc00040400400000c51c3c33040410000303c3400d0000000f00410010131c00453104044033011c0430c044403034c314c004d100100013000000010400f00f00000435003c0000040300000003100100310301040003c70c00034c040c304307cc0c030000fccc0fc04017040307000003000c411f30340ccf010401103000000d3c0400ff013000040d000f0400000001031400c43030310c000103300110cc0010040030cc301f701700040100000730000001340c010d10c0d14c0000700404030c003c4f1d0c030c340000310d30001040031000300303100303013c0cc4000310000c0300051300f0010537040c0304310d401031031c040307041d000100c005310f01057000f300000330030c00c4050015103c030c010c000010310033040300000c013d70040000000003000300000f000d03000c300f30000010c00700331c31350f00300301030001001f0cf1001c130c0440f05300c00100031cc0740f000300010c0400000000053340c30c00d30700454c050040c403100001c003343000030c130000043000300000000f0000040010050d00c0000c000f1301004c3c33030dc1000000014000000c0030010c01000301c0330100010001030c00301c5f0011101001103100003000170c00000c0100000300000f0f0513cc0c010cc000303cc13005040035c0400300440c440130000030010c010700334fc000000700f00c07300010000100001001010300040c003c000033000004c00000000001030c00000d0c07d00f00000500000cc00734000003000400050730130000d50403500c00000001031400000103074f0c04001000030030310034401410433000050c;
rom_uints[148] = 8192'h10100001331000c0000c4344000d003010400003c10000013000003cc0d11103ccc00c0110c300d00c400004c050dcf300030c3100c50004100c0d0000000005c00c30034004500000100004c704000000cd003140c00c310103000313030003030304300c00300cc40337030f01010003030c13c03f140000104100405001ccc3000403d003000c300300000c04f000c700000000dfc140000003114c030300c5c000c014000000c0000040530005000001000010001c000000c400330040033c0f003003c0c333f1c000c04f0c0033c300000d00c00013001300310c0403c0003c0001005030340004000041175f01000000344000410000004300000f3001d04000f403003000010c0104001c030100c45f04c001000110031043c0100cc10300001ccc1c0043c10340334340c300040cc0000300c04300ccc0c0440041c0000030004d103130ccc4c001c40011004c00010000c0450033310c0304000301f3c3041030c04100c0440001f310015010c000315d30000030ccc3000000f001034c000000c0003f0030030341fc001000d00040010c051ff00043100110050c031003300103000fc003c1701d0100003004cf0030c003c010003570cd0000000c04034c0000300003000c40001000cf00000033c05f7043f3000cc10cc400030101100c00400df04001410dc3003c4700cc05310c030c01400010c000013304000d3000003000000400003003000030c7c0000300400c40d30334010c10c5c40400c0071050c0010141400c0c000033c0000007f44003003f0c0000031cf0f0d300504001400300ccc000044c37000000500007000533c3000cc40100c41314400101030000040001c01c043140cc0003f041300140040000100013c400f000001030f0000c0000f104401340070f40ff1c500c010101030300004333f10140c00303fc07d000073303000070400c330003013300000500c57000d0c4003c0000c300000c0300cc00003c0001d0100334d00cc301130000000033040030430004440070003f01104104300d1000000030031040000400400c01000c4030000030c00f03040301300010dc01c00c330100000f73c110010140c0c000041715510000000000000131000000010000000300c0c3433100c030c40cc40301000040000403000400c00f00000000cd30c0c30c3000014000030fc3400400030000400c7510000000c3fc0003034004300cc03040340000c003c03003000cc04c03ff0c414140030c440040040700034000cccc0000c500000130005400c10040c0000c00400000010010000003034100300031000100000010c040400304401303031000c0000007c00003000300c000000003c10004d00f100400030000cc0300c1500001d400003001c0c313010c00004000010c00110401300003003047100;
rom_uints[149] = 8192'h4000c1f040c0000c303003004040104000001030001000141400c000300000300030300f0000003c00004040c04fc0c40101101003c3044c0013400040000c004c0c4c300004000000005400c310f0cc010003c3000100535d43c00100004070d43050c034004000cc000c00000c03304005c0400000000430000fcc00003710c400000000cc045000400100f0400040004000004c1c01000000400fc41c00c1003040c40300001000c00100c034034000100010000000c1005c0003c3033000300fc000c00000c000000040cfc00400000400000c403051010001404030414000c004040000003f004030cc030000013f0010000003100c00c0001000c005004000415f00000f0100c005100000134c400010fc000030030000035c0000140d100000300000000004000300cf01000010c4000413000000000000001c0000cc014010c3010cd00c004c000c03300400c4100dd300300f111551cc0c031000041000701400f00cc00400c005401c00130c070000000030c005003f03000000f003001404000c000100007004030403004cc0c00071000007001c3c0c00300074000000004000000013c0003c440000c000f300010c00f00000400005441100000000034040731440c00013000000454000c000000300004000c00010fc33f00100c000000c1c30c40c000c00000c0c0000c0003000400c000c00c00500c000c003044000110c1c001340003c14c0000000100404c00000000330110cd0c010404f0000c00030c00101003101011000fc0500c0f04c503d553f00141000c00000c010000040400000034000305040000400004003c304000d000c4004003c00000050c4040040c140011f0050000003c0000c101010000044000070fc040040004140030000300c00000c0d004000401000000300070400000000031fc0000000001c00c0000d00c00003000000c13010004300000c0003400fc00cc0c011c004001000000000400000d000c000000c00dc0c00000000c03000505300000000001c00d10c03000000d30f4c030cc00000d07000c4044000c40c01100410000001c00c30130034410000df00000330430400cc0c000004001300004100000f3005030050f0c00040d14000c000000cc00004300c4000000300004000043440034040400000c00013c300000000c4c0330010dc40100cc500000100004000000000003000410000010030300100100c0004013000c01000cc400001000000c00f0000304000c303100000f01140000cf031054c000001c000010d00d1007000d04400000cc0c0400000000c1100000000c7d07c1c00f43300000700d300f0c0000030c0000001740000c0c007c010c10000000c003c0000c0444114400410c00050c001000001070114c4400000c4730010400cc000d300030400c400000010;
rom_uints[150] = 8192'hd0000c000010000000000c414d10cc013cc33c011300fc04003340340f04000c004110341403000c010f00403004000c011005c0f3100c10010000000f0000d00c00044700043110c00004000500c0500c30004c4d0d41137c404400000000040040dc0d10000100117f07000c0c031c5400000330370401000c0c073c0100003c040000001700c701000053041400cc040c1000000cf000040cfc1d1c0300074101040000c44cc3073f000130f000334004fc0000c00ccc0c000054114d10003cc7000c000c03010001000c00030c45043f50c10c0c3f0c0014c00433fc33001100003cc0c0c000c0407c303c3007000c0c50010433000d000000030c03c001fc001f07400d0400c3f33c170010000000c5c00f003c0f0400400cc0000130105000c1003003000100cc000303070f44000c003c04000d003c1c0000cc00430040cc450001103700cc000040000000000300040400070004040735300cc53fc00c0054005000033043000000000c0403c0000c01400030003cc1713c0c0c00000c0c0d07001010030034001143007fc3cc000c00000004430f000100000c0000cc50330cf00110c1c034010c301400f4000c0311fc04000d00110c344001043400fd00144100000400c3030007000c00037000c00d00c3070c010000f033000d3c300c000d3410334d0c0d0110c40001000004043f0d0c05313cc00000070000130c000c030c0400530003100cc00001f011303cc700004c00d4000dd331c40c10000304030c0401044f0000030504cc010000000c004000404441004304c0703c0300003000500300000057000400000c0c030000013d00000447cc10001f4000040430f004c70dcf00000340c740c010fc01cc0400c00c10c00000047040044101f00000700cc0070433110d00000075534d3730750130000000003d000014cf070d0c00410000f3405450c00044cc40000140000030303f0c7400c03c1040c14c0c100c000040100000040c00f0cc0030400c03001004c01c04c40010fdc0070011fcfd4730070c000c540040004c3c400dd3010030030d0cf000070007000c411000340310d030000c0c0000000c030c00300004f0c00000040405000000033100010c30000000c004fc00000400c403143d044d000013100c000c3c05001c10c3030140000000cc3c04d4003103040100f40d100010400c000c07030c00003037030111000c0400000c3000100000001141000301440145000404000cff0000171c04007c000000000c07001450010cc030000304c00404050f04c4301c00c400400c70400000000010040000c3003c101003000c140c045000c003c0030001fc47000dc0c404000f1141000033000c14000c03500000000cc01400000c0cf3000304ccc0c0c0f00c444000c70c00040c4c040440c0001c043000041000;
rom_uints[151] = 8192'h3400c54000c00000c04010030500350c30040440c03331c00005c050010050004010c04c000000f00c4001c13c00003041c3cc03c3c001d0035030341330c000c00c10004c00000000000c40000010c00043033470f50000001000c000041374c0040003300c00c00000c00c000c00000cc000100043004c00cc05000001c040cc00c000c03f0000000000fc4400004040000000003000040400c400c30c410030c0c00000c0cc0004c440400400000001c0f000000100000c00000c0300000040c0c00144c0000000c071f330c00540003040c01030fc0000c0040cc500c0003300400040300300500c00f730f0c00043d00c00000001400300000000000040f404c0400c0c1000100400c0540040c000c17cc00c430cc0500d0004730d000c00000000310034cc00c400040000c0c0000c0030cc40000000400040f30000c0400000403450c400f044500cc0000030d5000010f40100133013c0110044c100010003301c01cc10c0c000501110d300c0040000000040000040000000000c01000004c000c00000c0300000c3c0c0c13c000000c000000010404c005030f0005c0f01040043c040c00c00040054131c00000040300c00404c403c1003c0cd1000004c401440000c0c00c0c00f004004500c000040001500000c00000010007c00c47030100040010004c004c330000415c0c0c010004030044040000000000c0000c004c1c0c000000cc10004c4c00000000c000000fc001000300017400400300330000cc0c000c000d030500030000000d000cc144c044c430130c0c034400f44c0c000000030701400000100c40c407c00000003150000c0104c00100040000010403c400070c44100014cc400104c0104c0000000400004404033c140000011f00030c040030030004373001700040f5400c50004300040000c040034c0cf0c40040040c000c004d3000000c054053c40c0300000300000c03000000c50334000100000c0c0f00c00d000d0c10000540010c3017000000301304cc071004000000cc400c00400c30030c0cc0004c4c003f00000010000c440000f44c0004c000443c304c40c100000c0c0000040dc1400001000004000c000c03000c0c0c010000030d0000000000000d0f4f00c0000030c004c00003040000c0003410000c000400041c0000030f000300000c050f00004000c43004040040000010040034004f003c3000c0004010000300cc00000041000c01000004c0003047000400c40c510000000c003100c00cc00304050410030c100d0c001dc0c0017c000c00c004004c000034000004003c0c010300000c0500000c030000c0000c0c43100400007c00013000100000000400cd0c000c00100000cc030c00140040310c0000000401000c0000110400003c0d0003034040000103cf00c4d00010000000000;
rom_uints[152] = 8192'hc000000000c3000000000c0304004000000403300cc404c0074cc3c00047c0000c1000000340011c04540303cf00000c0114030004c7cd000fc0000c0000000c0d03c00004400403400000c0c00c031100c000000500040000c3c0cc077c10000f173100c10500050c01f00c000dc50cc00001034f000300010dc44000014704c3074c01040003400000000000c04c41030000c00c04070000000401030c4304700cc40c0140000300f7050cc04c034c00040400040033000000030001100c03430100000007404d04400c4c07000c40033c00000000c0030c004cc0fcf000c10c000105010c0000030000040440000404430140030c100000000d4c04000c0c4001410003000003143000130000000505cd0101014ccccd00100700010cc0f00300c0000c000000010dc4f0c40c0004c003000ccc0c0300010440000c03030f03c340c00c0000010c00001d340500004000c3004c000140d00c0cf0000000000f0044fc0000c50f0c0404c443050c00040000c10010000c41400100c00003000cf0140010000000000f0005444c40000000000040000c03001000dc0000400000000010040004440003000c47000000440000c00000d040400100000100c700c4040000000400050f01000c1c0014074c1105440100000003c40101cc400c00300404040010000f013c000c04000f031040000300c30c00030003010c404304030000100100004000030f3cc00c000300000005c4000cdc0443004000c1004303c7c0401fc400000c0ff4000c00000c0c17000000130003c10c0000000400c1000041c0001104000c001c5000540f000400000c000c100c0335000f004000c4040000c50300000c000c03000400c0040000430c05040c000040000c0040c0010004300000c00cc00c4f0000000fc000c30c04030c1040c70d00c000c303000000000010c103c0004c0001070000004c0100000c014003000000070000010c0d740000000000040c00000700000000030f0c00c000040c0740040100117015000003000c000004c000000cc33003004c030c000c04400c0d0c000100010c00000000040400070140c00c000c00700c100c0400000000044fccc00c0000010c0d3c000c000c0400cf00040400040c01c3000007300c04c00000000440040c00000d00c00c0c1cc0000430cf0000400c00c04c0c05400400cd1f440540004400050004010004000c03033005040040040100000000430f0010000004000000c00000000003c000100400030f040c000f0c00c01030cd0fd0000000314f000000000000cccc000c000000030003040304c005ccccc4000c4000000c00004041410000700d4cc14c000001000c0c0030000000000c00030043700073040000000d104331000045070010050010c000001c0000000c0000001c004000100c0000000;
rom_uints[153] = 8192'h1310000340c00000c070d0c010c00000401013c0cc00303005013c00ccf00c0000000040013000740cd0400c400c130030300000004034f000500000400100003014741c0004000010041030000000000c40f0c7c00010703cf040000301103400d03c400030c17400701000001003c1000040440440003011f0071100c00c04000000050c0c014400100c3100000dc004004040000110700000c000d0c1343300c000300c0100404000343d40030010000c30c0004c00d03174005014000000100c003000fd1000000000100030007c1030007d00144071105cc07040c0400040000000113130040311005c00700c300000100070c0000733c03030c000100cd000f0305300f000d0c00c005000c003003c30100000403334101030001400100000100c00000015403140143431304c00d001315310c0c5000010344d00c015000c1010100030400cc0007c00011045f000400345003d11100c5170044010103d0030001740340001d11040304f40000f0c0004343001001031000430300403f0c0170101034cc40d0000334c100030c000d0c000047c0011c0003003300001574010c00c00410030403c13400cc1c3c0001003c01300c030d430400000300c000033c400000c00007100c4c1401000104000300077c0341c300c0010303cc00003ccd403d0cc30f000000c34000030003040401000300000cc00c733000430403040c00400330fc00010c0300040f01130330470c00040000000004c3100c00401734700500440010d10001c0000d0c30cd0401440000000404c10400310300300f0c0003010413034344010c44000c0c03000d070c0004c4400c1c0000cd0c3f0030d0000031010c3140c00301013c030c130f7d000001140000110c4104001c00031c0000000430d7000000014c04d04d030105430000c333000c4000c40cf4007003100d0f103d074013c1c04004300000004004c1400300030000c10301000d5000000003030003c0001000c140400140030d03333c0330c4c03ccf440c004043fc000403c04300004014000003147443004000040c0004504300430033300004401d0d3010000cc0003c0400030c07330c04000c00df041000000004111c00c0004300c0000014000d0f0400c0033c40000f400013cf00010c14174c700c0004000001070000000cc34f1f000403c00c0000000051007d0000004300c4030001700010cf03cc00003f000301043000044411043cc134004101000003140010430500440c034003c10f000740130000000013130005050100c34001407001c4030000003300000003000010000005d00001003f00000310000c00030300cc0d030107c0530400030f101000100d001301000400570401400300d300000000030340c04040030c4000517003c0c1000040c0144003310c000400034c30;
rom_uints[154] = 8192'h31f00000cc13cf0000c0454074000d10d44d413c0004000000030c10403401010003cc043331000c4c1c131051000c7010c3c435000d00400000c101010c3d01c00000c300070304040011000d031c030005d000305d00fd0c5fd0010c15c3004c3405003004000c000c1147cc040040c0c1f11000004c0103d3dc034d104c001030030110d131c0001000c0c140f10c10000000000300701700000000301c7131434300003c0410c0130000101000300c03410000010c00000c00cc30cc0c010d3404014000001450c00001f100f0c001014f403171030140c0cc1540d000c0313300c3401d5cc1040033c010000d3000113000c30c0000004c000303000000c7c45040c430543000104c140133031003310c000f3c0d1400c1003130033c310c05700043300300101000c701000301f03303c1070c30110c500003110000c34310013140d314004170000f0000000000334003014034030d30f3130d00040f0001d104d310414000005034c17fd0304000010003c040c1c0130010300ccd01c10130d3c3070000470401100d4030174001000000000100c04001010434000d10c113c0c030057001d4cc0400cc31007c01f0dc13d403100c34000c00d411c0003410c04041c00100d501300001130101041c300010d4c0014c4040040c307c007043000dc30dcc0c5c30f0400d0000000c0104c053f503c11303000c04c07430000703410c4c43030105d14001104041410c0fdc04d0f000c1c1011c103c0071010113000404410c000071c414030c03d0c700c4c101c743501d003000001f0010d043030c4d014000003c00f0300d403010031400c0000004030cc47c5007311c443cc10cd040c3040340304044000c11f0001103410130410c0007d05c35000000030001330413c010403cc7310005050c7100c3c0010003000153f0f4100f100000370cc00010074043050fd1030c033701c0f03d0c4dd00c4330c104000344000001001001c1000013013101400335c0013cc70d035030314d3cc3300c4300000cf7000501134100000400100c00d000010c030100411043104f5300c1c004c035c340400041c00cc30001cd40d30c40500c0d1d1040000cc013010f0c4cc300013011c0014c410005c040310d00c01000c07041003dd00cd10431051df00300cc0003030000304400c4cc1c00f0010341004011c1c3d30000d0c0c0c10f0001010014001c74000110000100340ddc40030301071337440030004c000dc4007d0304c00730cc003003dc0001cf1cd000300131530001074300101000030cc003fc100053ddc00001c01c000001c00000000400c001010003001301cd0040c03d13103f700dc0c00010c130101001004c3003100004c0c0000007d003011c011cc3007700d0003011040404d0013030004d00c030000d10100030003000;
rom_uints[155] = 8192'h11300000134000c0f0c040004000303003000000333c71000003000004cc3300400000003c0c0000c040c0003000011040330040000003c3000140001000c00000c1f0300000404000000304f000001000c0007001c1f00dc00100c00000400000fcd340000030c0c000f00000100c0503d00040000cc00000ff003000410340c70000000400000100c0001310004001d0030100000c10004c0000103003100013000c0000c0304300001001c43000100000c0000010010000100001d10000000040000040030f30001300c00030431c4010303100c0c00100c0c00153c40000000000330c3000004500000c300c0303404153000010000300c0c0c0010000110c300010003150000003040cc00304330043101000c0f3003000004010410001f0004c005013003000c330431c1010100300003040001000c300000340c00030c00100403001000030c00000d00040c0d300000110f4300c110000d0000443033000004000330cc030d340450000004343004001c30301003030d0c000001000c01040003040014003000000cc00cf0000000000f0001033030010f101c0c30000f70c1033011043c000540c4000c300000000c0040f4c3000000010c3c0c3103400000100140010000000000c0c10105010000000001303401100430000c013f000004fc103140330000000c010000040000003c030d303150401000000c030f00cc0000033010003c1401510fcc300d0c00c011300d00000000000f403d0003000000000004000000000001000010040c301001303000000015070d50003010300000400c040430000c00f4033101100103301010c430010010003000cc00330304010c0000000c04000400040400c000450000304f0c500400000f05fc343014c03000004000003510dc104403030cc1c000300011000000100c0c00010010f000000430410101341414f1010000000034d00403c0300030000300300000105000c000000030000300041001013010000c3000300f00003001010400001000000000300001003000000030314000c00d00010000400000413c01301301c0330011010304300010300000c000030c010c000000c00040300fc0030c1001030fcc300000000300c004000030030000001031410001000304003007000030110001013000000c10c30004c111010f4000000000140c10000c113000c015f0044cc03003f44400000034007c0f10040000c103000000311731000004001001000400001c000000000330000c310030130c4d00000c41cc00074400300c03000040004000130f0cc3400030000400000c00040c01000c000030330c000403c00004011c00c00c100030010104300c100000100000000c0300cf010000c3ccc30f030000000104f00c0000003011030001030c000f03000000c0000300030c00000;
rom_uints[156] = 8192'h107c00111150130000010014f00070003000400f0000100100330000c00cc13000343033430003000000000000003000000101000033f0040000003400000000300301300044001d100000400050010310c01004030000304400030000030043000430003104c030330051030013401137410c1c00013033531cd04c34d001033003330010100041c000000f4000440300010000000003013300c003113000011d0c1000030431000c104000031000410033000000130340c03f0030000000034c13033044350100340003033300d0313c0030000c0003101040400c0c100003c0100c0c1f004c000037070001cc7000f100c33130400000c031000000000313303000040400d0000c130103403004300d000d30d003300331300113000730043011f00000f0000301103c40300001100000003000103000100150001071c003400030001401100033c004010001300f00c00003300300013347c33004cd04700030000070f0030400504103004310c0000001130d700000103000000331000000010003704000c10031001010031303100010c10000100c5001000310000003cc31010300100501010001014040100000cc03030003310f0000030c00c300030001000000f01000000070003c004331100300030003300053c000034c10750000c0000703000000000030f000c000003001c300170000004f00000000500d410003c473c300001007c10030005033134333000cc100010430300000103c30d001540f000f400300100c000000303000034c30000c400100013034f3000c03c30703100033300c00000c00310000011000100c000110000010000304331c4c0370101000c000100101100300000d00001301d40c04c310350100100010001130cc00000cc030303031c0100c301c0000340031c0f100000000070007343000010040fc01007103035014f4300100c000071d0130100cc0c0301c0100000100000100cd00000d000000000033330000000dd07410011013307001c1d13cc0c0003001131c033001001001000000004300301331d000f10000001000140301f00011330100350100030013041000003004030000000130003001f3c0000c11c00043000000337400300550001030003300330000f03005000f00000130d4300004c0000000c10000f00c0c140000303033003000000010171300c0000011301d001c0f0c00010007c4fc03070400010407001470401033010434f0004103434001033700010005403c100003400000001c0c1531003507030100500014c0c307010f00400001303010c0300004c003400004000331000300003007400c0cd000d0043007f003311f10100c30113000f013300300100000c003c000c11100001300c00c000c311000c0001000000000d0cd000000040114cf0010c011300300000;
rom_uints[157] = 8192'h300300000c0300c000000000030000017003033003033700001540c003d0000001000d030030000300300030030001c0304f00000033031143050003310003000300050400000030000001430000c30130000033001000014030310c000373000300300cc100c0400d0f0dc7313011c0100140101300c1033000001330dc030014010100300c00000073004000000001000300000031300cc40d033041434c307fd004000005000c30c70030003000300000c0010003000013030000c000000300300c000000310000430000300307310000cc00010d104030c131033731c010cf130000c3000000070104300704300000101000c0003000300000003001003c340033003300440100000c307501000303040000400f010311010010f0000f000c0000001100000405000434000d43004000001003030f00000000007100030340c400300300300043001100c00004100400000300340c0030040c7c0c00040000c4003413000011000143040c004100000330010c01010044330c00430301000310004c4c730330300000000100304300000100000001015330031000004f31040d000000c040300000030300000100010003c00f0d0001013340000003040010c404000c00003303300300c10033103000004040000c1000f0cc00c0400c070c0000333d01c003cc003c3000c00040000004401c1300040313010000c101f101030cc301037d00000000031000000fc103100100030000000100130d030033000304310100040c00413410c0000f0c001301003070000303c540100100f00c400013001013000340000000c300000040005400004013100334000c000013cf00710003100000f11f007c100ccf030c000c000340c3011004050000000000300004033140cf3300003c00030c70071030031c00030f003700001f00cf00030130c00300040c03c100043104000d41310c00300000400303104001c00041000c00000d04000000400300000000400000c3310cdf00000013300010c1c0340000010033000003001000030004000000401030014c0c004001030f1fc3000000000d00000010400003c400007000000003401c000c0000003100043004311310007d70000030101300000700410303010c0003300000330f0040010000400000000413400000331300400004c071000f030070301c00140030401003000304034330000340100c00301300000013000100310c000500d3071000010001300c00001701011700000000700003cc00000000010001c0c00003004004117004d100070100c0114000400c30000d0003030400004000c307004c00c000400003000c000400cc11000d010000003300000503030000000000000003400c0430c140330cd000010001370000000451000000c13000000340050110040030404310000303;
rom_uints[158] = 8192'h1000400000c101c00001041000c05001410404310c03c4500077cf00c0c0040000400cd54f100000003400c0c000040141d3c3f300010001300001100040c00000001003000340c0000001041010cc000107dd040c403f0001470000c04340c0cc30d003000000d00741cc00000401c0cc3100040037040c00c1010404510044000f4333c01100300000000000c00030c0c0403000130044000000c0d03340d300400c30030c43000000001031c144004001530400050005010004f0010c4701000700470400030c000d01030404140033c0400000030000c4ccc300c0c500004000430017d0000000300cdd01d4c004c300c3c0c00300050040000100100040114350c4030cf41043c03311f30100010075110310004001400003c01040740c00ccc100010d0000f0cc0347c0c0000113000000cc00530030040340010710d0030140030031cd001f00c004cc00c330005000000dc3c07000007f01513004030d03000000c00f03000004045000d5400004440405f000000000450000000100c04444c0d300000c403000dc44040411050400000010f330c4440040000c11403007001301470403100d4000003000300040004000c000c0000070c000c0d04044c001000c300105d000010070404400744000004000ddccc000300034c43034c303c035c3d1c05044d043c3c0c11141100101010043c00440014404c3cc01d41000c0001000c30000031001413003000070c0000114d100c0c170070100040000400430103f0033010f40003541500303ccc301c0c000000033f040400000445c0001030000000003c0c003c03000310034c0040c7003000000c041000000030301300300c301d4000403344303c004c4c14c330000d0033000030013c0043043000300c000404000000034000303c310003fd030cd0044010100000f03c300470000000300013001cc07731000c00c404104f0000f004430c1cf05c30c03141d1000000000010c0d40000c000005c001dc50c040dfc0300000c0d003003010030000c0030105c700c00034000000000c1103001010c1000404c003cd13040c0043c4c3cc1730733300014400c03503d100404337000540040f0103400041c044f0003000001c03001400f0cc44310011010c0c13400010010144c4c3030001300000304c0cc3000534000c4000440c004433c074011100000d00000c000c00d00013043000000104c005001740c0c0c0d0f0fdc04000003c070004000403007400c0cf04030000030040c00000003c01040c450003cf310730c0000fc0c00103344007d0000fc10c0303001310fc1300cc0104c100000441013300040cc100041047cf010f1c040000450130c100007300140400fc3030010007500300147431450001003745c100000000c0c01105c003030400d10f011005f000f3003044;
rom_uints[159] = 8192'h1100010014410040000c4040ff01c000040440c30740530304403dc30300000000f0c3c0030f0000c37000c001c0130303c411f0c103c1340110c003030300c0000300c001000040000004430340000000004043f30001000c0050000c030001c33001410000c0401301030c0cc00c1000c0c040c300300f130c40400c4107c00703000000c0000d0403000003000c030000000000004400004c040043c13400004301400000310001030c0004070000000343410000001303010014c00000314333030300005113c00c0000004fc001c40107000000034003c1030ccc14004000000c4104070000cf030051434d00003313f40c000c00f0c0004140030000c10010404f130001000c00d40015000300071c0441000f0301c100c303010001c0c0110000330400000040110c01403040430001000137f0405033d001cc01cf010103030004040100130001cd0000c0044043010d00c03041c3c1f10100c340c000c10103c0340007d0414411001343c343f0004403c100000000040c00c300c0030301c304cc0000400700430404010f330003044001540105000d000c40740314c00740400000304041c003d40513030000400003030003004000007003fc43c043c0000c000031000f0001010000c14340c303000c014000000300300000c00f000041100f000c04700000f1030103cd40044100010030000303010303004c00400011c300004300430000cf0df40f0c010003430003050013000300000040c000430041c10c0000d4410400000f30100c100001c000004cd30100c30000c14c0100c300c10700000033c00c01c000404317004f03f1c10c51014fc143401f00045400f00003034000000f01030000f403433301c7430300000000c14c44c4074c0300050100cc00c04103010cd5c00011c5070005100140c10c010d33310c44c0000130010c00f10405000dc04710000fc00100000001340c044d0cc3c001330043c0c00000c0010100000303003403c0c0c4000c000c0140c303000703430300030004c30f0043c101f0404f0f03000c03c70001040000030c0100030d0000100c004c3300010300030003c3c04c43030000c0410000100100cc43c0000330d1000fc501004000414000034cc0030c03313f03f007c0030d4f010143c10103304301c4cc000040003c010100f00301c0010100c1010140c103000c03000444000041c045004003030300040000410340c040000cc30403400004c0000000cc00030001000d3000000043000000c50000344001c0000011101000c000043300004000c401c00300000c4cc700c00300c4000310000733000000000541030303c017f000c4030c0300000000000040000003030041004c05c1d140010100c0c0000300017300304040100c41d0030044c0c00010010054440c000507c10000;
rom_uints[160] = 8192'h71005000003301c0030303c31040c4d0003d47114fc37300004000004400047000c0cf30c03c000000c03000c00d0001c37c4141300040d000004c030500010300c00347100300704000000300c0c000104300000343fd30303011000001cc0300104300330043000100f03003503300c000304000c03300000001337000c040f3c00104300000c0c0300000d1103000c0d0000000000d0001c100303014130010c00130f000d30030304100c100c000031010300010134400000031cc303303d00c000000304c00c0750003cc3034c100100c000c0430c000d100d141110000500c00401030c000000c0071417340103301c0c00300000000c00000000000003011301000c040440000010141cc00000041f074130000001033304040c7c00003741c0000113330000301f000cc300000c0004000c000314003304000030001d0000030c0c034007703c11c000033004000400040300030fc4031300303405000400d00d13cf03044c00031700101100040000000403030c3c7c0f0c7c3011000000700c0134000340030000143400103000033c000010011001030f00340c0503f3000100000400000000000013041740040131000c0c003000c3000053303c04444c0400c300000330001c3003400d1c1004000d074c330d000040000c010c300400d3dc000471333c44000c0010440404034c40000fcd0c000ccf00000373f00cc40400400d0331344d1003c0310000f00000343c4c000f0037cc100101040003d03300040cc001000000101003305014100003c1030c003f33041001100c70000001000f0100301000c010050fcf0003000003c03000070010110300001cc700110033000c003003000007103001313000400c04300c0001110c300cc0000453030c7c00000030c0c10333005cc34d1d0030030470040300c0033730000403300f303c00c0000330c4300f30374c00000f0000000c0003000730033c3000300f04000003000d000000000010003000000003000c0003700400f034303305c00071004000310000070104000030043c0000300403000000400000c0440004001000c0f0300c04000c04100010000c0d30fc05300c0334003c034c0003103ff3400507000000000400050005040104000000000cd0000004c104c1000d1011d00100c30133700304040007d0000c30c00f300704040c4fc140000c041f00030c05010300300c07c00000100004c0000015100001000000001004c3403300043c0c074000000000c3307c401030f30d000011c00100030010101004000000001001030043030c0470300000004000000370001750013c001c003000037000040df01c330cf0301003001c300503000c0001000400c001f00c00030c000333000000300300000f34130010000410f030000000370c003740000330000001000;
rom_uints[161] = 8192'hc0000c4000000000044010000300030000000001c074000c434003c1c000044013100000400000000000c000014100030107400c104f0003c00400000c0000c00c10000000c0400004ccc1c00001000c0300f0000000014300d0c000c100c1030c4c4140000000000000000003000c4c0c0040c0c503cc0d0001004741000cc4440530000000c0c30000c0000310000000c00004000000c34000030140400000004000470400c01cc04000000001400000000000c03f00045000400004000d0300000400011100cd014d400c40cdc0001040015403400100c300004140000400000c31f04040c0c31041cc014003c10003c00103100000000100c004400701030441c10300005c0004000040c00300fc0d0d30004c030dc0000cc0007300040d440000300001c30010440504010000000c41300c3400000001c01300010041403000000c400000c00000000304c00c40c40d0f4043fc0d0050c4000010c00005400400c0000000010440cc0c43c3000000c00000cf10000307100c0040c0c0300003c0030000c131c04c0000007030300300000003d300000003ccc00033c300cdc030000d0440000041044040710140cc0c000001040c400cf04100c10cd300030cc3000000014003000333030040c003000300c00433c00d0400004340f3c00c030104c300700100000040c300cf0031300c03300004007030010000000000340404000000040300d33334044000404c0040000041000c00010313130d04400d00d0c4c4c00000740c430000c300040c1100041031c001c000cc4040c340cc0c00c0c00030010c4000c0000300000c000000c10cf4000dc00c00000003c11070007f010000f0000043100d4000113300cd33400c00010cc0400c030040c0000035c1000303000000400470c7400f0100010000c00c30c10000000034000030c00fc44000c00c0c03403c040100140c340d005030070c000c034000040040000000cc000000f0c001400003c00000004c000c010c344c33000c400000cd000000c001c000c00d000000000c00407c0001c0f0004000c3130103437000c00000c00100000304004c43000001000000370c70000400c00041400140d0040c45700000014c000c00044103400000c0c0030300c0c4c000c00c0c00104000d000f500c300000c0001c004400000c74000500000100370000d0000c0030cc3f30100000c4003000c03400010007007400c0044400003c04004c0000305003c000110c00c00000c0000000000c003c0030300034000300c400303d0000c0c00c0030000030c00004c0000000000400004300004c3130043003000040000400cc00000c700c013004000c0c0410100100344500040430dc004c3410010f00d4104c00000400001000000407040c01040c00104000000c1c43c01d0000c000040c40;
rom_uints[162] = 8192'h445000000014100000000c0c7000044001010100330c03000d0414007cc004100003000005700000030000c000c30c00010c1434000100000000000f0704000000040003c10c0140000300030f03070004030c0130f1c70c01430300347cf030473c0404131d00000040fc0040440004001004f07000043c00453cf10033000113c50c0013c0c7000000371000300130003404c00f001c0ff70f00304400000303f1000700004005000100400f04003000074c000c01300005000310100001040103010c0c010130cc3000000003c3d40331c00004000c0303c0370d0403000474000cccc0c1cc00c0100fc00001c00000045313c0400c000c0c03400000004c030c13c0003140133c01400c1cf00c00c1300000013400001d13004cdc40c4040c110000013c04c003040007c00cc010400004030444000000030440c7001c04c40431000c3c004c0c0003734040100ccc44c434011c0107d1010cccfc0d050c050401031c000000041d00070500000101c004410305030f0f0000100003c044040000330c00c34c17c00007dc0300304000400f000000004c000300500c04f007df0c03c3040d00040100011001dd0d013313c000cc0000c300000cc00110300011c3333f300cc4ff100003304c00040000000c3330c30003030004c0ccf00c001c40331c04500403f00100000c0c0303c0c0ff01000300c00000400c30d347000c0dc01cf00001074c074c1cc4c070000c4003c4cf03030404303f0c00cf05107d0f1c00400440050c300f130c30000c00000010340000040430010010010c3fcc70000000040c001037dd00f0c000400f3003000c30034fc00c004000cc53c10000c03000004000030000cd0004f11d003d000330000030333004003100000000cc13040c0000000054440001c743c004c03c033105cf00043300400130fcc3d40c0003f3330fc004510404c30c051401440c0300000c030d4c10000300cd00000000100c0003300004000000000c0c3003f0c300cd0c0044030fcc30300140003000c300f00c00333403330100100c00071c4000c0000000c00d5000100040400000fc00001d4000c00003c0c0030000303003c0c1040403010f750001101c00c000d03c03000d10300c3035c00000c7033033010000100004cc400773000f4340040003c00c03010440030100000303073005300c3034c00c00000c040c1f000c00cc00cdcd370c030000010c0400110c00004c00030010030000001c3037031400f000340c10040f34cc04c0130c11000400300004dfd10c04100c0c0013c3000c70c0040000403030000000100c04030c0000100c0030c0000013030007001700c0c4403000f1c00005000c00140d010000c000400c30d0c0c00c03f400000c00cd0cc0410c00070d01130003f000400000050c001110003440c0030;
rom_uints[163] = 8192'h1034400c0401c0c43700040c40004004300040f0300040400133104040c140c00033c04cf440101040c00c07c0ccdc3070f00035d0730fc0d0430030033300700000701041c0000c400000031004f3c0043340703c1c301fdc3070d00070f10040fc51343130000033d37103c0c70404140011c004000010300c05c0c0100000003cfc000000071011c00000c031c4f00010c000000000000000305030c040003030d0303c04000010405005040001d00000400004501440000000c0000004040cd0300000310000304013f3f00330d000030003f04003f0c31000fd15700004300400030c00004cc07034c000d3d440f0000010340000000040000030001004c0001034c005c5d0407cf04c400f000f401cc0430030301004100cc050474000c011000003c100c03000c003003000d000f0047110c0c0004040000300010010000100003cd0100170c04011003033d05cf010133000000c0001c3104000033003c400ccf000001005fc0133000000330340304000104c103070010000000c0300007000030c543404c00000c0050f03c003300c0043043400400c10340010407c3330004000d150401c1c0000dfc0015300017034c0003000001010103c1000c10000cd50005000000070c70004000100f030001007000010003030000c004001433003334000433045000c1000533c10001300100017f0000370000004050100301014744104300030400001007041c3fc1001300510cc0000c1c7304c04cc30c300001031000000d43003d300013007c030000cf410d331f00000101030c0704000f0401000133740c771040000d00030f0003000300001c0c304d0000030f0d00004dc040030004cc33000004000001f7333000040043013400030dc01330c500000000000040003100d00f0300c0400c0104cd0004000103030c000c0300050030100d050f0c130c00300103c40c0c1f0d010000400040400503c0033104c00011010001000c0001010c0400c400c40000000000cc0440450c400307c003000000000c5101400d1c0c00000ccd0000070dc01101030000c15301c40100003000003013003c03000010330004033d0004100c34410100040c1d30000c034c0300000105c0030000010c030000130000300103c000010037030c0043c13730c033010300d000000010c033000d00030300010304054c0c00c00000033c3c00d40400cf0c00010c400d03c1000000c00c0c4101030f030c310000000c1005103c0700000c100034c4310411330c0000033d04003010003010cf00000d100000470000000c0c00040f031d04000c0700c3d007110007000301000000c14003cc33070fc0040337c0000000001c00000f00000004333f4001014100000100030001030170d30103100003001c0c1100040300cc0701030c070c0ccc0c070c00;
rom_uints[164] = 8192'h1c010000c010d00cc0004333000d11d10c4400c40f04043004401303174311140c3000030c00000430c0003c340401300c000000050410001c0501df0000000c000c30104003000c00000d0000010403c0030000000c0404004d0c0000034c00030410054c00041001dd000100353035000405343004100000c00c30c3c1000d500500110d0000410c140000c0000007100c0000000c03071400700c000001700004030000330d100004100c40000c100703040001043c0d0000000c7104000c0013000000054f030301100d0000cf0c0037403400c003000f040c101f30c0010c300031005100003cc0034007310000000cc70404000103000344033401030c0c00110c0000040c004400040c0003100000c0000001001c703c0100040430041c0010000000000000000c04000400040000000c30003000000305f031000c3c0c0301000f0c0000000003cc031001044f0401070130330d000ff507000000300401001c4000040c0c0c1100044300040103c0000100c0000c01000300000300330410000c000c0000004000000500c1000cc3000000004d0c4000cc0001000c44c003000f00171f00c000035c0703074001c430000377033c00040010000000700c0cc0040031100300040010000000dc37c4000c3104000000cc01340003300f041000003fc000cf0c003041000f0cc000410f1d40013c00070130070d0400100034041100030c00001c00300d1c701000040101004c00010400000005000000040004307f01c00001000c7c000f0300300400030003004c0d0407000001c30000100c00c0040c0f000070011400100cc011003410001c05400d0304030d01040c0c00c0000c0c0c00010c0300000400040c00101431000030000015341d10040500c00100007d00c31f00c1310d030c0d00010c0401000041000c030c03071c400c00000d340d1c07744004001f34030401011030ccc000c0005040003000000300400000000c0000403100010000330403033f30044400000430040004f030000100000005000000030030030704000303c30404100001030d003c011cc43300000401100c4300050700000103000010330c040d04005000011f003c04140c400000040000100004041c10070000010c00300c03031000c00d01100c0c0400300000170c0010043c1f000c00000c40104f41c00300013001000001400cc40fc0cfc0000400043001000404040000003000003d01010004d00433100d070301c1340500030404010f0c3d030003303004d100030c30130300c0004d00000f0103040c00004c00030001140c00470000d40c0f100010100030000100110300003c0000c47004000c040c050d000c04000410000c0001c107c00c1c3010c00c0d040000000100c407040f0003140003c00401100104001cc010101c0070300;
rom_uints[165] = 8192'hf10000001c03003400c007414001c0c0c1c0100004f000000000c00040007000000000404030000004000300c005c00004000cc0034c1740c0cc0004400000004000130000000c004000c0c5000030004c3000044000c00000d0c03041c0100015c000c003c5301d00c3c000c4030cc70c000040040700c504010000c4c030cc040c31100040c5ccc000c004040044004000030000000040034c0000700100033c0c110040000c0000314c01000000000400400000c0c403000000d03c0000c400400000000050c30000c40000030000000010f300f370043000010000000000c0000cc403c04003c041071043c0c0303000fd30c100000101000030000000004000430030c3300041010c0dc04003cf3cd0c0000000c0c7c01000c4004dc44004c000000003c0000c0c14c3d000000100c00f00040303000c30040330c0000400c4c3c000001000c3451143c0ccc0001101c00000000cc30000c0c000c0c40303c0c037fc000033100f0cc100c30300010000c1005f001040cf03053000c000c000c100f0100110100000400c0c1100f00d01c0000000000c004000c30c00400f0c4340000000f003000000c0fcc10000c300700c0400400001011c1103d0c0cc1010004010c00004c0c00000040000c330000cc4004c00000300c0c0c00040000c0dc4f04100400d04010337004000400000c4000c0404011030040050031c03104030004300c00000100c0cc30d00c7cc400f0c0340cf03c001c1510f413f1c0010044030c00000cd0003c10000010300000000050000040003c0000033000041c30000010100c1103050001003010c00000003cc040d04d300000d04400c73c000c4c4000c0cf00c0000c0000f00340100c0c00f0c0000c10000000000003d0cc40003c044003040c00c0c00c404005004c107c0014000f030c10f0cc0dc0070c00fc0c00d13003cc00010000c4c004d10c000000040d0010340c000000000000dc0000010f400c000000f440c0000431300400c07740441c0040d41c000000014010c030c000300c41000d00c01000000c00f4000003000f00fc440140dd0c000c003cd010c00030c0f3000c400000000c0304400000c100cc000c0c0c0c0100404c0000000c1c0c00100000000c00f0000c1400000c40003000300d1104041c400c04fc0001cc0c000c03000c00c00c0004054043cc000f100000c0c01c00001d00fcc00c04000003c0001000013cc30000000c01330c01100c0c0f040003ccd00c00c10004004070000c034004c40f00c10c40000c104010000c03000c0000c000400d000400000005030c0c0033c0004d01100001405c00034c300430c313f07c10c0c403c00c000000c0000c040000004010500c0000110000001340400004141040400cd03000000d304cc00c0c0c000040f01000700c4c0000c3;
rom_uints[166] = 8192'h5000440c03310c04000310c030504d001c0000f40c10003134107013c0000fc0131330000c0c00030f000000cc003c0100101100300030044701500010100f3c440010c005300003c471100c00f0301004f4043c40c0003d10110050f0103040c0c010000003100f7000005100370cc0141c10110000c00470c0444c000dcc40000001400000043000c0000410c00040001001001d03d100000000170c50c0c03000004000c00330000000004dc00303c500000c4010400010514000035001c00300000c01000030010010333010501004400cc130000d40c011cc00500010000000000030400030001000c03011f40300105c000041404073004c000d01fc003c0101340cc0031000005c00411037dc3101410d0400303004001033043c10c150001040f0311300000350000013c351303000001030100d10c0430130404030d04000f04000f3c04c0000c0333000c01040c07130f030dc010005550000000004c01c0000c01044000400310013001414400410f0f03051040c000134530314105340010030c000003c1101003030000040cc0f11013144730000f0400dc01000301000043004440001f3cc0000c00c0cc441c00c30000f3c01d00030d33404000000434031017400000001f0403d000004101413c00d0000501c50334c0007000c000331301140c300700000105000017010370340103d0044000c1033f000304c00010c0001d0f340cc00500cd0c000300050f31010000731140341403343f0004014434c0c0010004f10000003d000040300030001105000000010000c1034005000000300000350031150000740f10000f4400000c0c0301c310c1453f000003c40000000400050003000100100401030c0c000043c0000c304340c0000c050f00030505130001c3403034c014350374040014030010000f300400041430304003040d1340d10040c70c3100131c04000100cf03000d0010100033c000c0010000003045000014000000400330d0c3c00cc03f00333503007c330000004003410100300000c300001c000f03030534040f300c04300c300431530040011000751000c4110c1010010040f0010c0c00110000300334cc13d1c400c0c3010000030400cc00000c013c00400000dc040c3005c014f400c310033c040000040000300000d10100401040001f30050c0004400314c33c00000000010350cf00310c40030303c0010000030000c0c004011c310401000cfc400dd0c103034000403134000300301310ff44040400010030000010c1407510c10f15310c131340001003010c14101c0000000c0010007300041c00c1300000f000144000004035c014d0d400340070004030300040301c300030300035c1d340003c57100005100004c00100030cc3050500001440000000000130303f7013000031003300;
rom_uints[167] = 8192'h40000001f13000130c001c03100c00c000410300030c001004014003c0c1003004304cd000000303040000030000c45c0330c3433003010301300011c00c00010000c1c000c00003400330c01000040300c00fcff01000c000034100c003000003d000015000c000000f70c0001013000430c0d0c0c1130100c300030fc3700c000c41033000003000410030700100c0000003000017401d0003000000c310030f30c000004d400000c3000c01c300014141100000130103030000300c00000000400000000110c00070000000c143f0030100c0004c00000031f000017000005c0000c30fc000000100000cccc10c0040034000133000c000c00000010030c00c00c0c10000f401d13010c001040000c403c00000c300c1c41030400140070001030000400000c04001c000040300704003310100001001c30500000040c003cc31004c3001000010100fc05000400554007c004013d037310c5dc000c0f000114c0003f3004cc10003c0000d0000c00300c0c005c1f0044f4c0100000740004703034f4340c040000000003011cf07000003000005400300030cd1000340c0c1f7700300003300003000004130404103007000c0435130030000000cc010c030f003c0040f03030cc340003000c00c0040c000c0003c4043c0030000cdf30000000300004333400301c04000d00001000100400100000000400c00c100cdf10000000041000000000000004f00035000000000d00c0341c003c370c00f0000c03001c11c0000c0000003cc000340c14c3034030303c0f30d03000510030c00c00300d00c000140ccc3c0cc007000000044400040c0c3030000000074c0c00030f0000003c00000004001044001030740c040cdc3300c4000cf00c100c00f00000c00000000c001c0303030730dc300d33044000f500300000f000310cc40c3c3c000c003f331034f004000001001cc00300340c000000000c04c1000000c000cd0000030030040000003000030d040000040000303c3010031030400300000300cc00000400000004010c004000300000103500000000c0003030cf1d0c0c4010003033300730c0000000000c0000300000300c0d1c10000500c010300000151c000c000300140000000030100c0000f0030000c003000310003300000c030cfc300c000c00001130300c703f0c0000000c0c00f00c1333103000cc10f4300300000030d00030c1100c001c000034000004470010100354130c3410c0040c0c0c040000003d040000300f0cc0010c10000010133000000014040004000030100c1034cc140400100000ccc400c01400cc1001cd00000c0000400000400300fc0001c404000000000c700c0010300c000000000c4c0001f0000c0003030c003010300c537000f004000c00001030000001100cc3100d10740c0cf00c000030;
rom_uints[168] = 8192'h33c440c44010c00cc000c003000050d0005c031000c0c0c100c300c00cc000044c00040ccc30400004040040104c00c4c004334103040041c04fccc40400010c00034c0c0c00c0c000000051004c10000cc4c1ccd1c500040500400007000001c3041300400cc004000440300004000300004740004101005df01040c000c0cc000c000000000070c1400000500f7dc000c00040010cc0100c00c00c00c0df00c30c4000c110004000100004410003010500c04000010004c040010010c000fc0fc4050c50c0100000c10c0f03c3000cc000000c40434ccc034010cc00444040f35001004013100043300d04313140ccc00340007c4000c00000404000000000c3300044400f0000404040051040000c01c0403c000cd00c71c04c0030c003000000c00c554c0c0000c00c40404c000c000c00c470003000100000030140040053c30040d0040ccc0000044000fdc0c500005007d001011f4040c073c010c0404140cc00400c0fc0dc030344004c034c00001000040c40430cc04000ccc4400c004cd0104403400c3000000c401d4000c0000000c00440005010c00000c0000000c000004000c000030300000c51c0c1c0030003077040c1c0c0c0c004c15400000c0040c0400c40c0040000c0c0400040000041c0c1300c0004c0000d1000c340cc040400c003d000c00001010033c7000c0010340c0c0040c0000c4000030c41000000010c00c04cc00c070f1010c00c0530000040cc04004ccc00c40450d01f000013444000000075400404c00cc03445004c0003300cc07001114004000c440d14000001c00000f0000fc000c040df00c040c054440cc4403000010040030100100dc300c0c04000004000000c70000300000cc4c0c00000000c0040030000000001c000c00000c100100c040c440ccc10100010c4d0004000000c0f040c00500c0c0050004c404cc00c004c04044300cc101000040000c0453000c00043c400c0c00000c0400001040c030040000c054c00103cc54000c3cdc0000cf300000000030c4c0f00c050000c400c0cc40040000401000c40000404000710400040300c0c00001000c00040400040000d000c4c000040410400fd0cd003000001140100c1c400c0000100105000c0004000cf4ccc0040000c500003c00000440001c000000370010000cf014c4c04000000cc0000003001cc0300100c0040000100000100070000d400004010c400cc00c40014d00000000000700f40400c000fc00c03000c04000f0000cc50440030031c10c044d0f041004474c00000400000c4401cc0c050c3403003400400c0000cc004000130000000000010000c0050000c3300501cc0543040000c10400430000c0540c4004001c4100000cfc00c0c10cc00040040c00cc041c0000044c00000100001c00c40c00d000c04004400004;
rom_uints[169] = 8192'hc00d0000055100000000c3000400004c003d00000000110000073400400c40000013c700000000000101300000000030c00041000c1005300c0000000341030000110013000000000300030070000f030040030c3001441100340003000d03010070004030330044005c040314030300100011100010003010030033300003004030c01011000011104000c00f000c030010000000071030000c0001c0f4010300310d30c0041000000300000c00000c003001c0000143074100000414700041cf0000000000000000000000110cc40300000400030000001311cf4004c000000d00000c0304010100070100c0040704c300350007cc00010001000400000003c0700000403f400000cf1404c4003000c1fd0dc0044f0c0044000005303101007114c00000500400040000133030d0100030c33103003000034000c10141f4000c433c1030401040040001100f00004d0007701c4d07000304000d40040000000300010304413000040307000073c0000c00410034c5000c0030500000c100000c00004104031d00c00c0000030017c00000030000000044000400041c40000003c0000300300004004000000700300c414010303010030000401500000c100130c0003003400300011000c030000f4140003001030030f10d0c100113000000000c0030040710c030331030300c000034cc004040334000df000000c40310c5000000470c0000033300000000003c03100071000f0000c0450000000f4110300010000004430010000730c04c4c30004404000101c00050000011034300334d0311130001000000050004310000015000c0070000c00700d05003011100003701050000413100030000030400cc0300301030330100001c01003d000303000100d001000001000010101310011c003443440c00300100010001400013100c00c11f0d00c00f000c13cc0003004000f07010c30c000010010040100100431070040300d3030031000101010000010d00013700400100300001030d00330301000000001c0d0010000301c0c10111000f0010f0d00003040c30000010000010001000000010f00c300c034000003010c00303400303000010010000c030700130030000d0000000000300014000010d004010ccc00004010404010c1c00c00100003103130030104c0010c40341cd100041c00003c00000100731c00003cfc04c1c01010d400000000c00000c0100100031070141d000c03403140003003103400030040150000300c1000c0340000040c0130040003103004500450003c00000043c0c3000001c0000000011c004100300100003330000c01000030000c041000003cf04000310310000030041c4001c00c005c000510050000100000010340000130000100301340131004c100403004d703000000000d00004010f00010040;
rom_uints[170] = 8192'hc0000130104040303340400000d331c00103000040000000d103000000c0004300cc0440004000c000000c000303030300000c30ccf3500000004000000c000000c0003000c00000c4041c00f70400310501cc00003110c0cd11300000010000400c000000030000030001000000000400c0403000050051c300c10047001d000304c1000040000000000c004031030000c00000303100010001000c14330003d00000040c0150c40000004100400000000000010000c00300c0c3d0000c30450c30c0004c005040c071000041030014c3c003d54000c3c70000000c00c40003000110c44001004c000101f0c01001110c4340030001000000400300000040c000000010014f000cc043c5000000c1004c110000cc00000030330005c00310400000053c110004001040000000c03300000143030000014003c030001000070130c000014000000000c0000043c0c10011404103000170433300c007030300003003000f0310000010034f03040c0303000000000100000400014300d40001000c01105700403001000000001013400003400000030003000000004110ccc0ff03430301041000c00d000005000001030005d005040104010001100401010301000000c00000000503013000110003040000c0040f730000030000c100010c0040010304001dd01000010c0c0040c04101c140000330440000c015000140050000140fc000000300000003100000000001000c10010300000343f0030440f30000c0410303000100300141010400040400000000000703030d00010000c0010000030cc003003000300c00c1c0010c000000400107400030400103410300001000004c0040000003010303000410405000100014c0030300000000c001000001c04300c03001010000c03000f300310003c0000000c300c0000043fc0000c1000c0400001f00007030c1000c00c1000300000540c0000000c03000000300c003014000000001c000f003000c0004c000c00000031c03050dc1c000031100030000000000000000000000010000010000c34400f0000000c403000f0000004000003000030000004011001010c003300040004c00d1051c0300000003000035010307c105304110300100000100000040c0cd0001c1400301430000030300000c000000d000030001c1040003300033000001410f4c4000000040c0f030c14000000c000000010c0101100100f0030100c0c00003000010030000030310c10c0004d1300003414c110044d30000c03c0c00c11c130000cf00000003004030c0c000c04500000110000001c0000000013700003c00140c0001440000000143c000070c3030000000c00c07c1cc000000400c3c0000c0000000c00033170000430000010103014cc001c50001c05030c00300000040c0315000000000004100;
rom_uints[171] = 8192'hf000004c00c34c0040400c43d0c0c100c0c030c000c03000040c11100003c0c0000003030c30000c70000f000100f10c01c01000c1033400001040cc10000000d031115000400033300f0003000010000010c0334c3c0100414c1050001003000310ccccc000000000001300c40010300d1003cc0000030000000c13004000004031c0000400c04041000c0cc10400c00030000000000c01000000000100413000103000300543011f000044c0c3001000130000000103c3700101c74043031404000cc0d001030304004000000310c40033007003044434000000054100000000f0000c30c10c0300c001d3f3c133cc00030c0001c0004000000c01c00001011cc00007c40051c05100c50110d000c0f3c000d04740c043c010c0000000007000c00000c01300c10001cc10f0000000c4000c000000c00f00041d3dc0000c00c40ddc0043c3300ff03c0f000000c0003010c000c5000400c101000030d400004d3000030c10d0110000000104c01010c00c340c7110000037c35c000033004000c440c015000000000000310401c000300000000000f000f04c0c00d4000004cc03004cc001c0400400000100c00100100000c00000c00303034104c0003400f4440000100000014c140304d000c00303100300000cc3000d0300c00cc047d000003000000c0c0c0501000c104400c0c00100c11cc00c014c404c4f40101f7000300000400010c0c000030cc00c0cc0f043041f40040030130003c10003400030003004000c0070011d0000100000141330c0000000c4d001d140c500000fc40c070c40c000000000c0003034c00000000040101000000301c000dc003300c100300501f000303003001150000000443001000c00c00000404c30cc0f0340034150700030030150c140004300301c00f0100300d340c3300c300000041403c400100000100f0034f041c4103000010c0510300010000000300c0340400c034003000110400f0000400000000003400000400f01000300c44010004103c00c00100010710cc30400f040040f00010000030cd43400034000400c3cc010c01004000003c411000105c0c000000040131000100c05d00000100c0101000000030100c00004031004cc040000000030d000c0d70f00c3400000c000004000030f00d0c03000400005003f3f000573000000000d00403430010c1cc1400705007370c30cc0f0000000013c00340c40000300c0c0c01000d0c4000c0001000000c00700c000411000000c30431300150110c034c004400110c00c0000c001c04cc0031001011d11cdc10100040010500100000fd1000430000c0000300000010330030cc300000c3010034004c0c0f10340000c00000000c03100c07f0041f1400c104000000033004c400000001000003001010cc0041000014c000040003100000;
rom_uints[172] = 8192'h47000000000107004101004013300100000d0c000040c0410041000043c410000003c04003000c047030cf300100d354c300013f00d13dcc01030013c7010000cc70101c000fc000430017c0c000f0cc001c1d317010ccc031000c1c3c3000004300c0343030c530007050000c0001003000f75c0040c1300044000010410403000147300c000047033000c04350100c0000000000001011cc00c00003000003dc033301041000c0100f0104c0c073000100000100030010000010313440007040c3003c00c000004110c00143010fc07043f100000303000ccccc001d13c000003000c00017d710000030cc001cc10cd0010400c4300000010100300d000040c00001043041031543c13c10100000313f1007400040c1c040c1404f140cf3c43015c10003f103f40000f01000000330071000f304300400c00040d300031000040000130000d000500000001007c40001c00034c1130040c4cc33100df1c0000030d0070c01000314000043c045d10c030c0040344d00c403400c00c00411f0050d0c00c700f0003500000001d0300cc0000300cf004c010000030340c1d010000c4300c4400000c000c3d030100c010d3c4c0340400c0301404310c1331c70003cc0041d000303011f0503000030cc400f0c00c010f003c00c000044c0003000c000f3001300c0300110c3011400d310c0011d400000c040000130c00104d41370003c1100100030c0104700340c0107f40100040014030000c7030c405000c000000003300040c0003c13050100010033c10000430100304115cd0000d3c070c00000300005dc00d0000000cc5c400043100100303c000fc3c4000031404100040000140714440004001070c01140001101c10100c00037c000c00300000000000c74040c304d00c1000070430003c0c1030401434500c0040003540007303d01c00cc3c300cc1c40000c1030100301d00043d30033c041333001c00033301fc00300000010c4000c01c0c00c030000500d4f000400001d3c1047010043070c00000c4c30c003c01d0005000000c000400d44000c0000400003003c10110034300040401100703100403340501000304004c0c00000010000300000430c1040c100c0c471c4d11001100c0040f00000005730104d10c41031010000c0c30f0030103c0340401100c00c0040303330000000000737051413000fc00c000300c031d0c0000c00f0c01f03410d0dcc10d000000040cc0101f0c0000c4033070100f00303c0003403004000130c00047c0030030c005300000c3c0040001010001d3c03411000300410004370c003310000030040530011000000000040004701000047dd3c013005334031300040004000d01000003031c0c34450c030000040000cc401003030170c03fd01100c54005310d0405044fcc01411043c4000070f;
rom_uints[173] = 8192'h400000100000c30000c000000000000040c003fc100c007d0400000400400030003100c0000cc3c0000040000400c000000c4c04700000c00c00c00c000004c0cd00004300100000c4044400c040000cc0040c41c0000c70000000c3000cc0c00d00400401000c0cf0040004500400000014c300004000c000073040c00040700400100000000400000c000000c0c0d0004000c0000000400000c4304c05cc0040000440c0c0000c0000c300000c40000c0000400000000400c3003000400c00000000040c000001000000c00c4c43040043400c00cc1000c40c4c14400404c4004c00cc000000c04040004000040000004040100000000000c000040000000000c000c0445000000030c30000c0045130040010400030400440000c0000400c400000cc000434004c030c00034cc000000c0000000000000000030304000c040030030000000c000034c0004000450040000040003c0f10c05430034004005c004000000000f0000003000ccc0c44040000c040040cc3c404c0c1000000c03050c00cc30000000c00000c444000400410000000000010000c010000c0c004c000cc0c00404000000c4300040000400000c000104000f400000000c04000174400c00000300000c0c0400f00050cccc0c0000cd005c0000c00c0000cc004c0000004030500040000c04004c004c00100043cc04000400cc30c04c3c0cc040c0700300c104000000c400c10000004c0400300004005004000450400004c00441f00000010004c00c0040000c00cc440c40c00000c0001000c00000000c404f00004040000304c3ccc3c0000c1300004c000000043000c000000000000000040000000100000040000000000444000c40040c0000000000000000034000000004dc400000004000cf000c05000c0004c7300000400c040000000404004c00c300c0cc00000000410134004000c000000000044000000c000004c00000000c004c00000000000c00040400000c0040000fc0000010030c04000000cc4c001003000000000300000001340404011c003000cc44c0044c10000c00000c0c001c4c100c00003c000c0000034000c0040c000c000000c00040040003040c03000fc0300000c00c001000c430c4000000c0000c400c00c0040003c00005c0000000c000000c10c000000400700000c00000000c030000040001000000004001414430000400f13c40043000000000500040000c003300010c00000000003000030004000004000c00400000000cc00cd0400d010441040004c00403304000040c00000000c04d10000c0c000000040000000004400000500f3c00c0000000004040044c404000000000c0cc004044c0300000000400000c40003c00000000000c03034040cc00d03000040410c0000000c00c0000000300033400c0000c0c0000004;
rom_uints[174] = 8192'hcc0f10000010000000034100c40003004413011310330cc40077c700010100010133030d0034030001110c1c0c00011070c7300d31471014cc300c14f000f000000003c0010d00117d00404000003cd0000d330d00301f00c0030fcc000c130c0cc0044000c0c000043013003f10c00c00f300030041c1134c01100c10003d011f1330034110003c70000540400c0c7c3403010c00c3101411101440010004c303347f010d1f104cf04104000000c0040c101400000003d340c000ccd030040030c41007c0004001010050000300dc30100001300030100c00000c0405130d3000000300407d5700000c001c00c50701c005100000110007010000000000004f030d010405004c33000d33040c1010c000104510030c400030cf0000110001c0000017000510000d004c00001014000300430001fc43110040400c3c300cc000300f3100530cc030750113c00c404c1c00c0100c10d3334cc0c1c300010070030c00334053434c3dcc031403cf0304d00010004c040c713030014cc00cc4100341500d031000300040010030f3113c0400000001000000034d10003c0333000003c050000000005400000050003d310d05c3000d00cc130c300d0430000c333d0f000303fd100c0300030400c0000f0440000c0030107430000001005100f00c0100010d100010c300010cc30014003f1c000c430410000300101000c10c33037c0000cc043f07400c337110c0d0c03d40400300043c0300500330300f0104333f540100000c3d0404c00f001301100040cc3300000000001034c3d0d00010c47010330310c00101050030000c0c00400040030003400c00c0001000dc010c10f040100037100001004000c03000100400007000430000cf40001000010c400300710c0d710013403c1c7400714cd317c1101300504c33000030c000fd00030c013f400100331f30041000f1313004100347104040c00c1311301001c0700004004003fc000000041010000f03c400510001470f0cfc00100040003d0c4071051000d0700dc50000000000330000c0003dc451f405005000140004000010c030cdc303003c17000331300000000003000300303cf0c1000003100030000c001001cf00001d0003005054300003010c41040f403c000140000700140cc30704100001403c03000cf4010101f07d0dc400c00303030153030303cc4001000000704100c0010040057c00010f00c10070c00114d000010013000404004d0001c0ccf0003300000003c00c010140000ccc0f0300070100c03100040c1404f0300100170c4c0110033001c0003d0c14013004007d4001c3030dd500c7400003401340000d100050c031c4000c0043030d0040000017030003d1000343d73c0004100c3010041370110050000005d0000304000c001c00000001714c43040000000000;
rom_uints[175] = 8192'hc40dc00000440300400c4040741000040cf00100000010001000000000c00f1400003fcc00440000040c40f00004500000300301050000401000d0c0c34000c000300000000000040100c3141700000430300030cc0000ccc040c04c00c30000c04071707010000000c300113f407cc00010c03000c00c004014c000c000c0c0cc00500c14000004004100030000007100c400000043d0c4cd3c40033040010010d000300000401000f0cc00c0004040000000000000000000040000d0c3c1f0c0010000410044307000000cc0000003c000000000040fc3c0300033c13500500044000000f3010000c001c0000000c0410fc0003070001030c04000000040440c0340c00700100000300040c0c0000000c0df01c3c0cc00000300c0003c00000300c10001300400c000c00030044000100000010000000000001341304344407400c301004110c0c040400040000110000000403001447000cd0437c40c104403310301c04000d30c0445100000030000300004c00105010044030010c003300c1cc1334400004300c00000c304007040000001030000c33400c34f40d35000c3d30300400000010010c014010114c10100000044000400003c03011413010710000000000400000100000000000001c007010000433000411004c07c1003c004000450d340000110410000070000103c0404003003c030003c00400003dc54c0000030300c3000410041c40444011c000c00c04c40c04400130cc0c3104c000100cc0073301004000000000c03001030404440000040c0d0cfc00000000345000c0c4300c01c00000030c000c0c0c0000117000c000000001704c0401070d0c40100c01c0000034044000000010130c000010c00c0c4c300001100303c4045000100c010c0004c0000c01714100040403707004073000000000c0043400010c03cccf051444030004c04000040d300000000000000c040dcc0410000f04000004304000000004c3f0001400000c3150030340c3000d330f10000c00000c0000000000004cc1c00100110004c400c11701003034047104003000400401000c00303300440001000c0010300000300334040000015000300004100cd13c0000c01c000400040000130410c0000c00c004340004000300c000c000010404007c0c3f01330000440040310c14140030000c01340400c3000f0040031100000001000c000dd1310000045034cc30c00c000000440c1c0400010410300c0000000c31c14c0c00000030040c00030300f00000cf7400000c00000c007110040000c00c3c000ccc004d4c0400010d00100014000c04100000000c0004000004051d3400040043044c07dcc10000000001110440040c000000340004700cc1040f0000000c300330f410303c000c3c000cd4000110010070000f0c000c00110c0c00000;
rom_uints[176] = 8192'hc000c3c0d0001000c000000000c4400c000cc00030103001004003c000040000004300c0000031c100001001044100ccc000c0f000100cc044030340c00003001000107d00c311c0000401000c000c030c151fd5f0c0001143030000f1d030fcfc3cc040000000f0440010010000c440410051034001410c0400d00010c0c0703f3c000000c000c700004c00300000041c0000000410040c0000cc3431004c0300400001004400500c00c1c0000d0000040400014000c000d0047000000c000c0014c000c041f010014000000051700001000003ff00cdcf00700000c040c00010000d0700303c141004c0c0f4000c0043030404710000c0000c00000000cc43030041040330004cf00000c05040000430c00c00c0c04cd44044003004cc0000400000001000030c00004cd1000000300043001400000000cdc00cc3007000000d03c00000c00000441c40c4c0000430c004400010304310cd0010040000015000000044f303070030c3000cf340004c00c0d034000000cfdc10cc0004d000c30400c000c400010c00c0c071c440c51000704c000000c4001000301c3100011014c01000d00c00000000301000040100c04300c3410c010000c00040041000140040400400045c0000004f000110c040c03000f040c004c00000004500c00c0005000011004450f33440030040000040040d000000c00004d50000300010c1c00c0cfd4410013050300000001070404141000044f01c0c004300fc50000004000100417fc305c0000c04001100030005c00040c0004000cc400070000c1000c0000000000400000003000010000000c0000c40003100404110100000c000100140100300400000f000c0000043003c0000c0c00000c3d0cc10000f3000c00000000040000c003041c4003c3500d003000040400c7cc4000c0740070001c000c070c0000c00300000cc1430007140003000cc0000000100300040c000c0cc40c0c03000000c000300f0017000c000300000c0c000330001d0c4030c4000030f30000000c45040c0c400033000430070c14cc0000c00004c0001c00340c44404d000000c0cf00c04000400003440013170c000044001410004004300c0040401c01040051040c000440d40000100400d000f00c0cd00c0c34100c4d0300001045010c0400000c00004c00c01000cd00030f130f003300cd0d00100000440c00000d700c00f00050cc031104040c0000004d301001341007c000000c0c030000404743004000033c00134c0504c00001c040d4043c0c3400c0c1500074040000c5000044cd000005403000700000043f0041c30d7000400540011300007c00000cf0000c01d3cc01003300000f0c0304003014000c04005c041c300f00010300300000110003140304fccc040540c4100c000c000000004100d100c001030000;
rom_uints[177] = 8192'hc00c34f0704c04301000100030040040430010d01100000000040f04301c00c1403400c00c0000000000c00f4c04f300441411cc030d50000014c01001000400c0000000004010040000000c001000c4c000dc1f0c04030030103c00053003340c10400004704071c000340040003000100cd4c3040011403c03340c003001400000000000c0c000d0017000c0003000000000000030404000c1c030c0000c000000000cfcc13040300f0010000cf00000000300000330400c0000000000000000000c0044c0c00000000004c0000f43000340407cdc437c303d4470000004c0000c0010700000c00c140c7000001c1fcc104c00000000300000000000011c0130001c001031004c00c0343001000f0300cc00007404c0d00f53030030000010700017000410010040134c0d0c00d000041cf70014003c0410040c3000d13000001c000430700c0c30300030c31534004d040d51040c330c440004dc007000143000c310340cc5300cc40341c33000cf053300c47c50d1f4c0040c00700c03c0000d01d00010d000043c1011110f000030c00000414000c00010c053c330cc30311d00c0004000040c03741c1004100004003c401000c0c0c000c0000000300000000300300140d400000000330f01d0031000d4f10000f010c0000000013000700004143fc041030041c03000341000f500001c00030400000c00c0004c1c001c0003300050c0004400f13c40004c0010344dc3110440030c503c4d301c1cc0c030400000000c4000c4000040000010400001c030c000300013000c0034c00c00000003000014300030400003000001d00010100c0000100040f0c030301000004f4000000030040c000c4c10430000000440007030000010000030c001040c3cc0104300000c0c30003010000cc0300c00d010000000000001010c1000cc300400c000f34d00d050cc0440c4004c00431004130c0310d00400000000300000c130000433d3d00300000c03000001d4f3f0c100000444c7010c00c0041330010400100000400f00003400000004000130d0013010030000c433f430c00003000c00000000dc0000300114403030d1000001010330303c00000c000000c01730004010c40000031450400c00500000f0303000d00430343030001d0304034400003010c300000c00000cd0003003c040770cd0000711c04c1000003cd01c50c40000ccc000c010070004101000010000000ccc3cc000d0700c500010d0cc0c40d301000c0004300004c3300cc430fd335404014040004c0f40010000040070f00004140c0005000cc00341500000000c14f0100040d00000000000130400000000330334010000c33433000c000000c3003403100c50300c31c300f000c430000004c013014044040ccc00000000004000000f3400f000001cc00070000;
rom_uints[178] = 8192'hf114000000301001000040304040d003050000c4c040d000004100000004041000500130c00000c0c1cc0000c04cc1c0040000500340f03300cc10fc310c30010050f00c4050c00c100000d3fc00c3c000007000c3ccc030c3f10300000c414d10f00c004000300cc300c000f0310f3c00001040d040c0c1404dc04cc0301330c3ff074040c0034c1cd0000040034001c00000c00003c0fc00004301413013f000c04400c00c0104403030c000100054000ff40000d0000dc0f340c0010f00035045c0c0c000000000001110000c03030301c03c000300000c444c04344c03c0040100500fc4c0000000c04000f03f400c0150134f3501c00000000cc00000c150c30c0000c30004404005d371400044c315c4c00001040000dc3c10c4d30041c310c000100cd010340303003000000304070c0300d4000000c00cf0707c000043000000003100000000c03cc0c110c01d0000c104c33c411050f43c000000314030c3030c00047030400401c3c3c7014031300cc00d0c1030300c03c400f000f000100054cc000c00c00100c4004dc7c00000000c00700035d0003c5003100d0100010000c0001500c010c004500000c0f0030113300000401000400c34c000c700c0c040c00000000f03010104c10003c00440075350f000d0c000400cf05c400401d0004004c010c330030c0c050400c0004c0400c000c050c030107003005c00c004f10c30c000004004333300304100003100c03000030014040400c307c1500000054500c100040c00ffc00007c030fc0004003040000013cfc10000c04000c00040400404c431c3444000310c00000c304c04cc00343c15d3f4c0410043c03000f000030000d31c0c03301003c00310430004430c003cc000000004c3c40401400c0300cc3000344c5c5c0000c0c1430cc043c0c00c00c0003c0cd3c0400c070000f3cd4d3c0003410c000041c0040300c404ccc300004c0c00ccc000c003000000003400c0c000000004c110c04000f5304f00043f01000c0c40000004000000533000000000c3f400c44040430000c3000010000f10007001fcc3c00d3000c000c400400040cc0100004c71410440300000cc0f000c004000c30000544c0cc0c003070001c0c0c4cc000000c00000c0c001c004f4fc001000d4440044400c3110400c00c10404301dc104c0030000000400000010c05c0040d0c0104400000300cc0010300cd004330000004334d3f441c0000000c7c000f0000c30c3d1c04100003003c100004000000cfc3001c40d404c70c03034c004fc43000104003001740f13c070004c003c04100400d00000c100130000c057000010dc0430000403100400c00000d401000100000004340c00cc000000503303c0400050c0f000301140004004c0040000041301530003cc3000f0011c001003053000c0;
rom_uints[179] = 8192'h40300c0070000c7c0c0300000c00c00cc00044300000000004c0000000c1000040000c3d00c4000004044c30c000400000c044f400000c100000043070000000000c0cc10030000400000c41f000c0340d041000c3c40c30c0c04c0003004000d300f004040000000000000d0034040300030334c0000400030000403c444000cc00303c300000430040003c300400043c0d0000000030003004c001010014000c00440000c0f0040cc4000c400000f000d0040000c00c000c0000100c00cc0c0c0400000000f010011000003000c00030000f40040000c00470001004040010000000000c30c0c0000000301007f000310100c3000300000104d40cc10000000340000034010040000c300407000000004700c0dc400040500f0c003004c00c00440c00c0d0c000400c0030f0c0c70000100004400c7000000000c4733300004c00c434c000c100f0000100000000000300000035f00014c3014074c4000c040004c0c00c1cc5000031c10d1c000c0404003000000d07001c3c010000c0403c0000001c7c41000cc40030440100f00c000040000000400440c4fc044000cc01033030000c00000000c10000000405c007300c040d40c0000c000c04c00cf0144c00400000c00c340000c0000104dc004dc40000000cf3c00c000000040050000000000c00404c033f0cc000070134000303c0d1cd000004400004000c00004000c03070c03030c00101000c3cc1c004000c1c04cc0c0c0c000014c30c0c300000430400c04c000000404300400000c0000c0404c000103040c00c10030000c3004054000cc000003500cc0c0000c0000034100300c4001c4f00030000100d0c000005000010c07c400c040000340003000c0000c00044430000001c3400cd0c0004400030000013313c00104c4030033300d00cc04c00cc00cc040030c07c430ccc0004350c0c00003034c43404c0f00100c300c0c10430c40dc04000004c001001c000000010c03000141300000c4000010c01c0c30c5344000104c0000004c400c01cc00430040001405003340004d73010cd00040000000004000d0300000100030cc1c0004014001300000c00ccc000c0c00c331d000003040400041000040000003410003003070404400403000001c014c03c000cc4430c000cc00c0fcd175c10000f400000500004340030c000c0001000000044300000000030c040000ccc070000000c0710000000000000007c4403000cc00000300074f03c0c00400c00010400ccc4005003c0ccc007007c0040040004c4c0000c040004c0000001000f13070004410000040c7400003100c0040041000cc00000c400000000c500003c10c0cc04000c0c400003400000c0000040000c00cc0c00700000c000c00c00000c043c401c040400000001cc00000000c0000cc00700f100cc0000000c;
rom_uints[180] = 8192'hc30001c04c00030000000040c0c00f10c040c0030103cc0011c03000000d0d040c000400c003cf30c0000000070070c00000c40c030137010c30000000430400044000003000400000404f01000c310000104103010c00c0015330c000400101000040710fc1000d0d00410003300d3100c00003c003004c13000c03100c0c00c3000100c0c000c000030f0c0003d000000000000003040374c0030d05c003004c0005000c00010043010444c0003004c0f04003000c0031000100c0c00000000300c00400400000000000030c044100003403300c03000500000301000003fcc005030004c300cd010400044c0000004c0c000000000014000000000000044c4040c0030c00000c400c0110000c140040c3000c000004000001c0040301410c5000000f0444000004404030c44040c030430100c0c00400450000c0400405400c000000040000404003010001010c070c0f0c0d0000010003c300000040010003c30000c4000151001071100f10030040000cc1c100010c000103c301c00cc1c00001c300000010404404030f470300cc030040000001030d00000000c0000dc10041010000030cf00c00010300c00000130303000305074cc000030000400100c405030007c103400000300300000f0d0000000c41c00430003040f40000000c41f1c0c00000040403c40f000400c040000c0030c031c0000000010001550000030010000300c3004c0000000040000001030000010330040000070013011d0401004d30030000450c0fc3033003101f0000000f0000f10007c30103f1c00300c00403c0c3010300003304c3c33f0304400007300004004000010003000c4100000f000f0000000300043301d00030040350c400400000030004000cc0c0011700c0007403430fc000100300d03701000f040104000040c700044300c0c0004030010104000040003c4c0035005003c001000043000000043000000001f4c003014000030000000301000040010001c10cc0034305040c0004c3c0030400c00000c00003400000030000cc0000400040c303c44cc000c000004f004f03000000c0050004c7c410000c0030000f03c0c000000103000035040c100cc40cc3c3c00003c407000cc00000000f4140000030f10c0c001d0dc01001430433013cc4f004c03001000c007c4000300000000030001000000f1d0540c3000045033000040d0540000003c04000c3100cc00c0000410c3c0cd4c331000000004103c051cc010010010c33c00000400300c7c033403c400c03400031000000500004101f0440c011050370100d00c300005cc30514440cc0c04c0343004000c0030000000c4d00000c34400000f000cd0000033100000000000400d0c304003c00000000040f0003330f000043c740030f0c0004004101110030c1c3100c010000000;
rom_uints[181] = 8192'hf300003400c405040000c005401074000400317f1cdff00000f1c0000100043004df1504130030cc1070300400cc0043000303c4001d3d400c0000f1503030001c1003100ddd03001000f400010100000c00400141331d70c03441000370d010113c004110053c1003c0c00c0170077000000310001c4000140033d00df13c7c300cc1010100c00c0311000004001131c000000001f403cd0311c04c503dc0f0003fc00004cc7030000034037010401c040f00300001c340300040353100030313c000dd310000c4d310c7130030505f0433370003c75010c40343430330040c00000310f1c13004035443030cf1000100175c1500003000441004c140c00030d04004301037f4d01701300300010001c300d500f01300044d0c40017c73051147000005c4c31000004004014030c004071f130350004c0300340330000040301c0343703030000411100034c001d00f04100c370cc1c4d414110c0cc34cccc000cc00051107111030dcf030000744300033f33400cff10314c0cc0345001c0f444f140dd000001d1000000430c0dd3430304001000c1001c00c01340000cc3f7c470fd0c14001000340000113300001c03c03510f14dcc000504000014d3044130040307c003c0400003003100014330010711030401040c140f003510000003000c00100d77000740304400170341070d030c0001070000310300100001c30130004d0fd300c400043144c30c10030000033c1d034c01050c1303c00703000f000f30003140000007c01447040000c0c033100001070000000001c50300010104331c00000700c300000530310300013303330001c000c4c04100070cdf00001f3c000c010057010431400003007014030103001000c0003c03000100000c110c00110f0c000000c300404041004d37000100004c40000000300040317030cc0c01c10c1c0001303d000173d000331c03c30c0ccd00470300000c00300c100400f00000000000c0000c0f000c004c04dc0cc7000d00110c00000fc70003c00000040000400033000f300431054c010101c74000c00c000400c330cf03100400070000401f40d073000c3004130cc0c4113f0c341300cc0300413004000040c13100003411470010d400c330c0c0c0003c0004001c304000f3000d03304400001040000100c0000003c0001c04dc103300cc4c40c303001d00000030f03000d0004c300cf3000cc33c4000c000c3003710400005070000c53000000cc035c0f703c0300400ff001000343d0047400c100c10140100040c4c0433c0070100003004000ccc01314330300400c30000c000c1000403000504f00011000f0c010f000703100c0100cf01000100300f03001c001300050107033d00070f010c0dd1000411430c100000070f040440c00d0000000030030400fd4d40c00100004000;
rom_uints[182] = 8192'h3111030d000cc4300304f1470040000c030101700cc00000f000000001000c000010c0100000040c000701ccc31007440034443040000510133044c003400d110c331c1101111030000c0d10001c0000001010fd0c001c30000050c473030001103000d015001000013c50c4114c00c014040043c003cc04cc0c7c04f00003330040000000000410000070000030d4c03000000310010f300c0404000070144000f0000c05030000000003013c00c00d0330000011d35333001c0003f0c0301f4d00001000f4c00040c00370010dd300111000007030010c14000f431c10000010000c0c0000031031013c1c0f030c0043d05300500030300000c33000010cc3100001410114300040004c4c1f00400d000c00473d031c001044f01c1000100330000004c001cd110000401010c004303c03000030100000014100004040005d1011100d1100003c000dd00004f10000f054070c11114fd730000000100000001700431000f03c4f00000000004000005001333003c00003341031000c5004700300034450131ccf000130010f131100001000000c4c00130c00011c0100d0c00000307000500000c0333007100c30000044c0004050001007303c00307013041100c04ff430d40111430300040300d000001c0113c00000100001000404d01033fcc0403010507c7c300000c0000d401d0144340000c0d0f00cc3003c73307030007414000d0057100410750000000011143400001700d0c007130c3410040434cc0cc03c5400000dc0001040440000404003070110300000c00140004014334104000c050300043000333000000034004101000004011d031c011000030770c100003000030440f0c00cf010000d000d0013c03073040313400001f40103003000300cc0cc0010031003033f04010c51000310310c000000001734033000c0000400400400c0500d00001f0040c03d0004f001311c15c000c0000030030000000cc0000dc403dc0001c003040f3c034034d43140cc40300030301430333100000400303c1300000000000c1000103c01000000d01c00c0040400133c00003000003d0010110c3000001000000000104c000d00000000c001030011303130c10c0100010000050000010003000000c110400304000003000400c41044d40004c00710f000014cf30f4000f0100000050100370100043000100014c0473f0dc3c0403c310001c5533501000000000040017040300040c510300c4000000c0033f340c000000000300007c4d400010fc0041f13004c000ccc10340c54c001000c1c10040c3c07000000040001400040030d000cc0014cdc10cc70010034103001d303000070100c0501040d0301c1001400010000d1001d003c0000c0100004001000ccc030c4f0103c0c400c00000c3300010000140300c03000403c35000;
rom_uints[183] = 8192'hc00000000004000c00cc0041101430130000150c3404003030c00c000c4400000c10cc0000000030000003c400037c1300000c0c10000c147c00503f001c3c000c010000030cc33000cd0c7400004c0c00c5030dc004000070f440c00c0c030470c030300cf044030000003030003c0000041033f000c00000300fc4d00030030c1c0034040400100c100c500044d100000000000310400300c0c40c0444004010c400c01c3c35000c0000501c3047003000000000004cc04c0004f4000c00df0c30101c00050c00c1005010340c3c1c1c3fcc0c4000c000001010d3140cd003000000c0c400030c700014313f10000f00040003050000004030003c0c0000100c0330340000413050701300100c04000034031010300c30440cc03400000140340000140000001d00f00c0c330c30c0000004fc0530000cc0303400100c033c04131c04c01300040000fc30c0dc0040000030530000005c000400040c0cc000000040c040044c1050000cc03cc000000004c01000300400cc030004100000c0044c001c100010d300040c4c304c040100300c00000c30004333440c001430007f0004400000000c3010030000003c03c400107f100010c1000430030c14340cc005044c30001400c043000f300cc40740301c14c4004f0000300c0004003000700c10300c1c10003c4000000f0400300000d0700f340000030c00131c103000000013f00cd03400c00cd44c1003cc10c0c40c0010044f50000514f0300414f00fd00d4f0c003c003c04c40c00000c000400043710350c003c004c00000073340c040fcc00c030cc40000c30150c1431c31400c0001f0c0030300000014c0051140000d000003c033010000000400001141c0cc000000330cc00300000001c0c15170c0000c00003c4c0300430041030c001001301cc500c0400007c300300c0000440400c130fd00c7c30dc70000f400c00001400340000030cc001003c0ccc30000c0000c41004303000000404003050df00310004c0c3300010401f00000c0000004313007000c30030000114500c103c100000140c0043300c030c040030030c040c0c00f5fcc000c000030c0010403000700c00c4040000000004fcc1d41c00003410000000c004041c003c0000140c040033f500c00030340400c00004f000f000000f0000000000f4003f03000c10000034000440301400cc04030cf41c4000000c0004301400c03010f004040013040c0c133c0c301000101c0334f03004000c340c0430000c3000ccc50c0034007045c00c101037f0004c1000000c033cc0c00030000c00000400001c04000c103cc4040000000f0c001300040c401031000c4cc0c4000304dc1010300c3004c00030340c0000000040c3d40100400070300000c0150000fc0000000c00d00c300430001c1405d4011001000004;
rom_uints[184] = 8192'hc000004000f004d3430010cc0051000c003c3c003350440c00300000003003000040105000703000000000500000000030c3c011c0301040c4110000c3c0000000300340000000c0000010c000007000004000c05404003300cc111300500400304050c10000c300000011010400103040f00050303cc00000500030000f0001100c01130004007500010000010000133400401c00000003f3001000140c4c410050100000007134000340c0ccd0c0000000f0300000400c030000c000c300c04101c00000001010013050000000000031010ccc00c0f000141040053dc0400d000000c0c00300000141c0030c0000c0c300413000000000304000c0c0c000f003c13000000345304000f04001400001303c3410300403c0f00001500000103003c00000140000004000c301c000f440f101440370000000c0f000033000010000404035330dd000f31000530000501000001040301000434030d100000c300054c000c1110003f03054010103cc5530000000c0c040440001cd4c0000f00400c0000011040443013370010000004000c00054041000000000c4004340001000003c103400f0304000000030fc1000cf00003030c07030000400fc0c3cd01370c003500000c01040c00301007f30003011000030445003f1000c001100d0d04000c0031c00004c40c0f003c0304300f30000030000c000000cc00300f37c3000c100000050530000403c00d0d0c00040401303f0100030c0c3005305410c3000073c3000003d0000000000333d00c1000100015400703000300000c03000c1d0300044000100c0103000f03cf00030c0c0000400000004c340c101000100305d30000100331100001110c040004000c0f00430300014c00000c030101050c00000001000030000000030540010c4dc10c040401000d0f0c00040c300ff0cf030f0f0000031c0010001013040411005031001f030033040033000c0cc0000000000000070c00000001100c00040041014300153000000130100f0c03000003000400000003000000000000030f04040043c010c040c005440000040105cf30300f000000130040000c400131000c30000010000100c001040000000300000c04050d3040000c00000c0c1400300004c005040c1100000f00430104004047010dc30c0c0500c3000001000013000000050c000c01010000003040000001c00f5c03300fccc00000000500010000000300040f000c0307c0011000000c0c1003100f00000c01000c00030003000500000004004107000100040c14100c070c3003300103010030003000000000c000000c0004000c00c00c0004000c00030c010300000cfd400f04003301040000000100000c0033030540440cc03000050c73303500c030000c100c30034fc31010011543110f01000403c7044300301f0000040;
rom_uints[185] = 8192'hf0000000303df4f45100cdcc5343c151cc3030140331c37300f44300303000000004cc0f754430c00410c04c3c0033d03004043030033c4c10000030110000000100704c000400cc04003d01cc0c101040300ddd0cfc7014fc40500c00c0047d001400f00c0cfc0000c07c00c0d04f0c4051301704300c30000c01cf30010400f173300430c0000400340c001040c01c000000300000003c3c033c0c114015401000310c007043044400040c440d0004cd417c0000fcc00103704040c0fc3030d3040000000030304c0000000003cc057004003000c110000303445444411c0010000031c03140004000100cc0303d000cf0030040030000000d3000000c00530030cc111c0c50400000007c341000dc0104c4700cc0f03001fc0c04f030f010403c77000c01300173cd740370003400000000744305000041040000c50310003300030000400d003c0d000004000000cdc100403c4300405777140c00140300c010000c40000104733004003c000c4c00400c0c3000c30000301000003c40000c004000ff3c04010c100c0040c0dc35c000d03c000003405030c30000c0c100cd0f040c73cc400400f000003700300030c0cfc10ddc300c7ccc00000c01fc50043c1c11070c33c3030070405007c000c51040c000cd331ff01100400034c010c030c001c0fc54030040003040c00001111040000340c0c004307030314c0c3c3c0c00ff000c77110c100041c0c170c000040000010c0000430110131c033cdc00d004c0d3f740f0000744005c01003010f00c0000731000445040000c10ccc00330cc300030000740313440375c0000c4df0c030d40000300cc04004000f3070c0010130c4000dd0c01c000f000530010c0000030cc0ccc0141000011c04d000044f003cc74c00050c7304131c033001c401cc00000c0c000003300cc00330030400000740d00c303015400000c000003000000c003c0c0c0c00c3c30cc3000fcc0004400000031c03444400033f00c010c000430000d730c0c004001000c30540030000f4000030c4300104011340030d00cf1f03f0010f0010000403034c01fd003000f0714000000300430cc33c00c3010005044f17004700100d000100031410030c0fdc0000c4c00cf00c134004030013c001d00040ccc0030003f4505000000000410303c40c300000cd0040004c0000cc0400cc00000cc0100410c3004003445300104f103400dd0c03044cc503c3c0040045c50dc040040000001cc00004c030000403c0c0044c114104f0050c030d0401710004444300104f3c00010000c1f3410340c40300310400400700070400c00001c5400c001000cf00d000010f47c300030743c00140c1300300d1000001030445040fcf4040c5400fc30000c0c0c0030003c0000340000040000104304cc3c40400ff03c3030330010c0;
rom_uints[186] = 8192'h4000000c000000c0f140000ccc0010404004400340400011000c40040c000003c0c000c303300000000cc0010000040c0f0c4c03c0004c003c0c0343033004030030000c0000000000011005003cc000000ccc054400c0c3344c0d005c0100040c0330001003c40d0df0000000000431f000430403010000404c040c3000010100cc040f010030000100000130c0033334010c0000111003410000310300f04c0345000000f140001c000010130043001000030040000400c100050f000000740c010400000050007015003300000000c3000100550c1040fdc00c000000000050000451030000000003504310f44c000100f4c00000000700011003c034014300301040053000c10003f0430014004017000c4f4c500c0304c0001c4000030007010000000040030003010011040000000000c0400c00031c00133cc3304ccc01000043000c300400137407c033040400000103f03033c1000c300004000000030d110c0c00000701000c03043cc3000004000037140001c7001050033c0003c0000ccd030030041000003c00040c000000030000001c0f000c004040400000c300000000000d00010003031040c440000c4f40f0103000140100040c430000014000f00101f000000000c0c0100c00010300003dc0304030030001000300000004100c00107310c303c0c001404c0c010103040001010d00000040cc43100f000c0030440f50c0300400c05000070c0103001000430c0f000c3c3c03c1300000c3334dfc0c00000003010040000030cc000000c0f0000003005301000003430030300000c4003c03000000d0000044300c00404fc04000100010c0143010000010000f0030c0030000340101043001400030001f00f0500d000030000100000000c400000c010000f0010100000c4033dd11145c4440004c3f00040041c0d0cc000400c00d04f31d0040f00003100f3c000110004040c400040c30400000000000030000c0003010000000c0401000000400003011331000003000034c00f00000040330300000000403030000440300100000000c0030000040f1003700c0000000c030c00100003010401c0100301000000400000007340000004300034510000043f00013044140004004100000c30003000d0400f3000c0d00000c0007000c001c300000100c4d073c0000000000010100004000f1434c0000111c0c0400044411c000000c00000001000000030c0c0f03f0c00f0d010000000c00000410f0004300c400c343040030c0c0004c0141f00034f700100c10003300000430f000004000c03304034004f000f0f00001000000030310c0000000f0140cc0000001c31100413f0c3000004c04000000000043003003000040c00011300031000300000000005c01030c0000040c41c0010005000000371503000003cc0001;
rom_uints[187] = 8192'hc40d00000cc000c00d000f010004030304110cc00435000cc0040000300000003c1c0101000004000d00010000c40d40010430001000440000000c57c000000c00141c00000c31000000000001000000030d01cdc30f00050c4000004c0c000300c407000000000004000000100010000cc010000c04031cf4104c100000c000c00c00300c0440000c00000000040000000c00000000401c044c0d001000c0000043000f04003410100000000c7f04000c0001000000d0043000004c040c000c00000000000400040000000100010c0300401000c3040400434cf3001400000040000000c0300000000011c11dc000001d400031000000003400700c000cc310c0030000c0070000100000070c0c405c1133d000c4000400304c0c0044130300040000440d440000050300cc01cc00014000044c010000030c41001000004400300c3c00000400c400000c00c03c000301000cc4c400403c00370504000c000001000d100000000300040c310000100c101000004f00304001010434c0000c00cf0c0100000000130c00000f000c050000c0000000040404040c0004000500001c00c000fc00040000000140040301000000040c0304000003cc04100434000400033c000d00340000000333000000f10000000100010c003331000f0004000070010001500004cc000f00030c0004040040c0031c04000400000cc04c34cc010c0001050000040030dcc44d440000c0c040100100000000000d004d00c104030c0003001330c1000350003033c0300050000000c570100c4cc40c10001c0c4040030000000c000407c00cc0001c00c43030000c000c0c005c010000000300c4040000c300000c000c001f0c00000c00050004c00d4c0c0c0300000c01003000070300000000030f0c4c003000030003300f0d4c11000001040000c00cc400030c00040305000001000c070100001f33000c00040c000c04c10c410000000c0c010000000000000003003003c40030004100c0000c0344110400330c0d000000000c001d400f000075040004c00000010100050000050c000c010000000304011c03000c007340440000030000000d0500340043010000030c00c03c104c0007570000c04000000000040004c0140c000c01000100000007000c30040030031d4031000030004c00040000050c0c000c0c0c0301030447c00c01000c0000c10c0000d00c0d0005001005004cc0340000dd74000c00300040c0003c0400000050c00400100000040000c00300cd40043c040000000403340f44c000330400340f000000001000050cc00000300007cc001c1300c7043001000000000c0c05c1000cc0710c0c00350004304c00130c0c043c04040004010c0114cf017c00100f0010300d000c00c0004004030c03000130000000cc000c03c000c0010003000c;
rom_uints[188] = 8192'h5f000000001000c00000f00000c033000000001c000014004030000130cc13405130300d30c303300010000044030301000057cd50c001310300dd0031c001000100310110000044c00007044000fd40000330c04c03700c4040003d03cc040030cc000f00003350cc00313101000407401000c0c030403f00004003c033041044300001100000dc00400011000003c0040000030030c00000031001310401c10014c3000000c01000d10c1030040040000d00c400003030d04000000c400140c0c000000100000300c3100000c0004c0f0031030000040510f1ff10003501000d000000300031000001010005c4330300130c71440000000000c4400000003f0400000450000c100004040300010030c1d00000d000f703030300cccc3000c140100c00c0400000c401310c010074111031301dcc00010001000000c000c004740001dd3001030007010c01f310c000f430410c0074030005c03c74c7c0c30304410cc0000000033030c00c0430f400c0000353400003c1370341010003c000030003d044c30300040000040d0301070000010f300001000305003c0c00000000010400440010cc001d0004400c34c000000000f001430003004013700c701047d30000041003c000303000040034105c74100000fc070100304c1d0000030c010103c00033cdc41077011300c0030430300cc70c30133f300010003003c014010000001f0100010d30040c0404400c0150c3100400c04144c0cc3cf1500000d304003c3401100000c031030c0d0000107003000030303001dcd00001000d45000103000c430100d000000d00000d1c03c03700d0f00000305040070d133001000f03001341d40300000100cccd40030c0300f107000430cd00130005000040000c0c43004000330100437003037014454011c0f0500070030c000004011fc0d00c000001370000300001f00c5100c341010050040050010000400300d00300f030003000000013cd4300400000c3040000030c0005c000c3000c0000001dc00c0001040c00010d04c34c0dc001303030403411000410f00c01000001f7400010400c101dc40c4d0000000001000333310000000744300310450100010d000000310033000430000000133300000000c000d130003f0001f010c010000000000010c40f010000031013d1301c010001400c30331c5000434405c30000c041000700751040f000c00c3100343c00d00300040cc00000c0353010000c03000c040000c110000044000cc000030c00c031c100cc3100c031004040100331030400c000001334404001430303013d000100003030001c0010c1000000000004c000003c13c00000f00030c01000400300040001c00000fc0030470c00c100000000c10c040000130004cc03f40c0050040007003043030010004703c0031d000000;
rom_uints[189] = 8192'h3001300300c0c0100000f0d1001100000000001010004001c0040300001000100000000000000000000c30000001033070730001f033004011f030003000031011d000300040000000f15000c0100030070310c01000400000010130c0c0100030003000c030000100013000001110000c40030000300c000f10c00010413000c0c040300033000000010000f00040000300004000303000030111f0000133c00000000c003000100003030003303100300001003001300001000000000000c000f000040010d40010300000300000300c030000000c7000004003000000030000100000f00300000004000cc00000000040333000d0000010310c000000003030034c0030000f00040000c10003070cc0300051303000300040c43010000001000130700f00001000c0003303000100c00041c0c0000103013100313013000f30000000300cc0000000000000300000301030c0003cd33030401001c030100c713133000010c104d3003c0030300130c03030311000c3004001000010030000013010c00003007033030000c0c0f00140301007103034000003d007300c0000f400c3403000001300000330031000033301f01010000000100030403300000000300040c1c0c0103000f131003340100300310430300003000003100000003000d0100000000000033031303000300000000031000010070040c000010300f0f30000300010001000043000c000000030103000c0c0310030f010000031f307c00030070300000001000040000004000000001003000f400300001030f315000030300000043030000003c000410030000300c3c0000340010100d3010001c34000c1110304300040005000000c003100c03100105000403131003000000000300001c003003010004000000004177c1070c04c003000103000d00030d0000000f1c0010c00310030d00000000000004004c000000030000030000010110004100300003001003000010031001000100000000c00000000301040c0001130000303000000c010301030001400c403300030300000c030f1100030304000c0010000d130030030000000033000311000c0000001000000c000c0101000f0c030403043000031000040300030c0005000c010003c0041cc003043f03c103000400031100030c300053000c00001000030003300130001c430300001f0331f10000010103000c00030330000310000001034130100f010f05003403100030d0c10031000003000300010cc3003015000400004144000000040400030300c01000000000000104010000010c030000001d000000000f1000000c000c0c030000033003000104000000013004c000000010000000100000000000001d00030113000100000300100300030700001310300300c003000001c000010000000000;
rom_uints[190] = 8192'h300c000034430cc0000000004c00001000c000cc43c000000dc444000cc00404071004701130c030000c04314040004000c0100040d000044c00100cc00000c00c3c041000000300500cd1d03000f000cc000044c0000400c1750030300c0300c04cc4000000000cc0000440000004441c00041ccc0000000ccc0001300c301df0c30000000c044000100700300000004000000000000c0000c00000305c00034ccd0c307df04c141400c0c4c00000304003cc000c300d0cc0c0004ff0fc0cc04c400000000cd0c0f010003cfc0004000c0c70400c00c1c30ff00000c140004c00000040400c0c0000414c70000d3c4cc0004410cc3004004040000000000400000004c0f4004c00dc4430c0000c00407d03300c0cccc41301000010300070103d00000c0c00000040310014c00703300040c0004000400d040c0130033c4044000034000400c0c4010004043010100d0030105000ccc0001007c1000c0c10000003c00040c000c14000135004f0400c0004000cf000f0001334000030ff00d14cf410c0c00000005c400000030d03dc300000c000040c0c3c00c3c700000001c70000c0004400dc4040100034cd313cf4301c711c40c0000c440c014c013040000d0000c000000040c0cc04000100c7c43000000400c7000000004c01000000c00c301400040030c0000d00fcd0ccc00001700101300040c0c00000100007100004c000c0c0cc00343310040000c00cccc40400d440f700c0c0004000000070034c40cc43471cd0000c4c000000000040000040000005c00044c00c340f00c0404040d0000100d30100cfc0dd40cc00000fc4000c3000030700cc340c30fc4400300000c0c0007040400d40004410000c004d00cc0c00c074cc4000700047d0c04c004000c0700044403300f401c0c0043c00d14704f030000000000450dc004400c4c75403000337540d00000001c0303057001c00000d40c10f1c00c007c0440c0014c000000000000400000cc0340410c40c0440c030c000130170c3000040070000400300100cc0c0c000404c000c000000f0c04000c0000100400cc00044ccf0434310437df00001540000dc0400000004031c000c44c30c0030c0007c0d00000040000000c1c001400c0c0f000c074070000000dcf0300c100c04000000301410103c033c4cc0100c0340000c03c40400040010f700c0c0040057100000300d4014c0c000030cc040400010004000000040414c7c004007000cc0000110c000010000000c0040c03430c3c4000c00000000cc3030045c303070004100d000c3011000cc000004040000010c0007100c0450000cc000003000044c00c41040040030f00cc0000c000010c0c000f0000d4000000000f0004010404003cc0cc0c0007c000ccc0cc0c00000100000400000004000cc00000cc7000040400;
rom_uints[191] = 8192'h1400d100c0011000130c0070170050130c41000404040700c0410400c40000c4c00003300043c040c0d0030300000c1f3070110000000070010100045d0d1003f1c03f0f000c0001000014001400c1cc00010c000400c0430430370c00030c4007040c71300100c0c1100440c0000004000070c17f3cc4c00010d10304030001040300000401000fc000000f100353044400000000000003400300001001d00fcc0c004c001000700013030503d10014400033000040c1d04100001035c4000010403cc4000003000100c415440003000500f40c431404431453d3100013000ccc0400001450400040000701c00c00c001c40010034300004f00000c0c1001cf00030103c5c0f0400c13c4cc170000740c0c050405150c00034400c070300c40070000000300440c04000140c7033cd00000cfc040004010c0010c7000d0030310040074c00c100017000c0c010405c03d0c103c0cc000054173d30c00400133040001400303c4000710c03503c4100340400705443d004c4110d074030404030040000014107000cc01310d43000cd001004000dc00c30000c0c4030d001100c4c10431cc0513000cc1300c044c040c00030c030c10ccc00400043000dc753c5c00340c0c0003c10403c0007c300c4015040000004f170c00030c31000400c1004501d00700004004c000c3c00d00cf4f01cdc0030c10030c0000c0040c00c540c10c040700f30c01d00c000f0103cd503074000d054010010133104f010000040d4f004f033dc00044cc430500d0000440c000044040000030000f010043f0400cc53300507410000300300cc3cc01004414c01041c1001c30531330044d105344f100014f4004c0c101003033000701440110c01300d1033c030040c304c004cc1000c13000303d3317000000c300cc1400c3034401c10c311c004dfc00003d010133c0c10cc0134c3f3c1331d40f440005350330c40c43100040040500000001030000000c030330000c1300000000030000300000030000c0f54cc0c4000f000000cc00f10cc473cd014c014004300ccc000c0d04030000cc1073000d00000070040c0401441400c0cf0000c0000f030c30cccf00ccc003300500c1010000d000c04000104000000100000000400043c50f0c0d000004000d1001c0030000015c4300000000cc0044010543010300c1f00c05400001017f040000010010340003c000fc00000cc000053f00c100000400050ccc53050cc700cf0400470300430f03c1001c007c44fc13100fcfc033504400cd003c0004450c05cc4c401d00d001c3000ccc00030cd000300010300343c3031011c00000000400c1040d0d00030335f000310300011300c5d700cd104333040c3004dfc0c441030f40000f40430100000c30013704001c00c00d04c00f4fd0010133c403c047054403cc00;
rom_uints[192] = 8192'h110404043000300000003000000103100011000000fc0000010350000003300014000750001000300000000101101040113c0f04003c00d00000110ccc0c110c0300300000103004000000070c0400003d030cc40400fc03d010010cc00300000030040c400000c000030000c00c0cdc00000000000030003070003c044f000030000000300003040000000404000c000000030000000c330c3040d000000030000c3004040000440400000000000000cc040c005400003c000030041010140001370004100004050110000c0f0000001d30f0c5c304001033100c010000104030070000c03053405c0000741c3d33001000500001c014700030000000413000303004300114400040301000c0040c00041c001ccc00000000100500cc300010000c010007003400000c10003107303c030000c03050300c110000000c0004000014004c00000cf044c4111c04c0c0100000f40c00070004500003000c000c1004143c31f00300051014000000030df00c0000000003010000000cf100314000150000000c0c4010001c0340003440140004004030100003040340100055100700c00700f0000c04030c00010000f00d0400040000fc0103101c03314c000001001000000334003000003ff404000cc0d41430cc00300000f0044c0401445c50570401107d001000400cc010407014000c0005000000004c441404005014010450340c0000000fc07140c0013000040400110440144000050c1004003c0c04c41c0003001c000f03101040001050000000001c0030353000003d1cc100530010c40cc0341000000c00050c0430140c00c0500410010410505400f00003c5303300341000c003c00c00c0000030f0010030000300003700303000c0030c00500030011c0030c100050004001f143c3044301033000734003110301c4c401000f04440000001070033c00400d03c000c000d10000000300100f400f0100413300000010c0f0000000c0014000cc401c00014440001043c3100110c003000001041010f0c4440003000c30c100c1010f31003000000010c040430300001130004fc0430000c0001c40000004307cc303c0000003010001c0003300003031000001100013400300004440c0000144000000c00000034000000400047100f301433301c0c0000000d00330003000c000c0c0d100c00c00c00003003000004100c0000000040070300000c00003401000414c40c000c10000030100cf000000400010c000cc0000100170c003007c4000000cc000c000400c00000400000040040005003004100000330000000300040003c040000401001c50000c040000000040014c1003100401700035000040030000300000000041070303c000000400000000000103300040c0c00004010c0340000010031500033cc000004000f;
rom_uints[193] = 8192'h40000004401c00f301000040044310001000070c03340000007013004001000103c300c30000000c103000f3c00f00040045000f0c04c0144000000000000d100704000400000000043c0030c00000011000d10f00c0000c0033d0c11c000000400c040404030c4c0000400c0010c300133100001004d00001c00000c00010c700700041000000000000014000003013000000000000f0c410c00c0c00003c01100000c010001000c000000400103c070000000c3000c0005000003331dc00c0100100000c04400d00000007f4300430010000415010cf034cc011503000000030000c001c0000014000000010000004470cc003400104000000001400c000004000cf400313ffc0c303040000c003f110000000074c0500f0401100c1000040c0000303000004000000004000c040130c00c3c001000000000330711000000c004003c404000000000fc004004000000c5c0440313100d01c315000010c00004000054340331003300307077003030cc30300001033000500c00000c40033c001100000c04c0000c00000000d0d000010300400004000c00c0000010d0004400130400103004003100c005000000300000041030c00000303d00c4c400000011010000000001000c0100001000010440000c01000400000cc000103c11c0dc40000140030c3000410c001000000000003003071c300010000000000041305010000400110000040c01d03414000000003c403c001000f000f3c10000c0d0000c01400043043000f00c3c0300c0dc0004040000c040c0c0340110034040c00000100c04000c013100c00014d440c000c0c003100113301017310f0010031400400003c000000000000030f03030000d0040000000c0c003000430003c00340000100300c0000c013330ccd00030000000c0000c0004cc00c00000d400c100110c04000510c3010c145000cc00001400c040c0c00003000000c03c100000300c00400100000030001000000000000000340040300010c04c000c0c30000001030000c31330003110cc000300000010300000c0c00300000000c0140301410100040c0010c000030000003c0c300000fc01f040000000000000000100007c00510000cc0000000003404000000c310c000750033000000040cc1c000000dc43cc0c00f00000c0300103040300404000701c004c000300030f000000cc10c03000000010001d0000030000174000340c4004051430007c4000340c400111040c10c015300000c030004000c0300400400000440c0403c000044401003c3c0000440001001000170000300001cf00004c00cc0c00000000000000000000000073c04c5470c300050000d00004000fc010143004000030000dc003014001f04001400300fc000000c000034030000000010000000c00013c003000700400004000;
rom_uints[194] = 8192'h140000000000c0c403c0000004000010044000004c401d0000cd4000c04c004000cc0c5c044c30000004c00c0100000c0f4c440c0030c004000340400d040000c0000c0c03010005010000c033c0c0330500004c7c000440c0fc01c0c00c0c003c034010000c00c000c00cc0c0043c404000331403374c7300d0004400c4000040400c000c430000000c000000c0700000f400000000400c0400104c10000000000001050010004070030040c04c004dc003300000c00043c0cc044c704000c04310000030000140000c00100c000c030014ff10004001c41007d50cc004c000000c000c000030000040004404c04c104c00400004c0000000000000000400c004000400007010040cc4010c1c000000007000c00040400034400000c4407104f3045000c0cc004400000300000000000c0c004c4000c000000044f0041003000f00000c1000c100400000c34100401c00c00400401000400300c330c001cc0c00000000030cc0401041c004c0c0000440430741c0000000044ccc030c40000040400c0043c43000004040400c05c0c00c0400400000c400040c110000d04000344441004004001000000c00c440400004001040c0000c4041404300c0dd000000d101040000c007000c040074000040c010cc40c000f40043c0000040001d40c01000cc103034030300400fc0c04001c00040000000c0030c040003400c40c040c1ccc0c00010030c000000c0000000c3d0000000c100040cd000c000c30000104040010333104004c310000000000030c0d0004440000c0c004c00c30010d0000700c030034000000c0043001c00c4400000000044cc0100d0003c030c4101000000c003400000040c03100c004c0c300000f0301004c001d033c0400040c100c0c1000000034c004cc7d44001014ccf0c50000000003000300c0370c0d000044dc00401cc3c04d4045f000c030171c00f004c004cc0c300000100404141f3c3010000c0003003040000c003c00500000c00400cc044c30430403300000003c0003c04440300000040cc00000c0004c4c0004c00000000300040040041000000c00400ddc500c0000c000000000000f00300000c00c000c010000000400031d0c0c00040000040030040000000000000013000000000000c40045c04340000c000c00740c0440010001000c00c0c004000000040000c45000c0000700000000000040010010000c00504000f00004000d4000c0400cc0c00000040c0001c000f000040400001740000000304c000c001c0130004000000fcc11305004004300000c400c0005cc00c0040ccc0000040000cc0407100000530c000000044000011000cdc00030c000001073c004000000304000500040003100030fc40c4007000c0c0043007c0010050000000010c04000000000c0040c44000400c00c000c0;
rom_uints[195] = 8192'h43130c00c0000100007000001700130003030d000001030000040300030004000000000100000000000c000000000133330c03c305400c030000400c10004300100d00030100cc000000004403000000000307010301000100030405000301000103030000001000c30c03000000013301000010c00d000d0300000c0000010003000500030300000013000000000400013000000000000300010000030c01030330300401010004010003000000000410033c000000000000c00001010000003d400400000004c40374004003004341001000004001000003000400033f0000130300000300c000030000400000010c0100c710f0410000000300300100000000000100000037030c000400040000030d0303010303000000000000003d313000001c000400010100000040010031000443000c0c041000010030030c0d0311c100034700000100000003cd1500100040000000000001700c0713cd03034000001000001d000001000004c000030003000040c00300f0000000030c030004030c4000c001404030000d000010004101c000000000000303c000000400000300004033000001011400000c03003314003300000d340001f00401310300143000034f03010101030c000107003c030400c0001300000100d100cc01c00000351c0410300104000040000c00000103000003000074000000030000000031370401000004001300c30c000001030404001c01000303301001c1043307000300310040030000041c043000041003100c0c0000003300000c0300000300000300000c300c0700040011010000310040104c00030000000001031040400003000130c000070001000000000404c0031c0300001000030030c10000004f000000000003004c000400000001000c000370441303100400300000055100c00c0111300c000000130100000000300310313030c430030f001000100c0003000300000400000004010000000100000f00c0030303040007010c0f01030100000c00010003300000000400010030300c00430f1d00050c04030100f40000010001040000010004000000010300155000300d10000040cc00030040000330f001004013030000000000000000000000433004000c1c300000100000430f00003000033303000004110001000030000000400f0701000d10330000040f000101300300314000400100000000c3001413000000030000010104040400100304000400330000040043300000100001000100033103000f010033000f00010c00d0000334400c00000300301f0000010001030000c3001000000000110000050400000100004430000c011430040100000301010103000300100103030001007100c30c00c130c001000fc000070003000000000c00000c0000001000030001300400c30000100000;
rom_uints[196] = 8192'hc0030040c000403000403000000300c00000000004000000053000000000000004fc3000d0000004000003f000400cc000c0c000d0000400000000040000000004401000d40000040044033000000400000c000cc0040000cc4c01001004c4007003000000c0000c044cc00000004c4441c040c4c000000000c000c0000300c0000c0000030040000000000c00000000c3000000400c00c30c0cc00c04c1000001400c00400004004c00c00000000701000c0c00c00000040c4000000405000400cc000000c0c03010000c00c003400000f00ccc01400cc00c40c0000c00c0000300000c0000000040000f1350000403004440030d000100004004000000000000c0c0c3f00c0c004d00004d4000c0000000050f00c000c0c7401000304000001c0000410000004000c03040000c00000000000004010000001300000000004100000000000400000040304400c400000000c400c0004041c03fc0004c000000f0c030d00040400000000000c0000c00000cc000404000000000c00004110004c00010c410000000c00000cc0001ccc000c0000000000000010050c040c0000c53d000000c400000c00000000c400000000031004400c0140000000c07c000c40c10c000c0000000000000000100000401400001415430c00100c000f30c04000000000000400005c4400400040440d00000030000000000040004c04c4040000400003fc43000000000000001c00041c0c000000040040400c4c0400000000004c00c00c0cc00004070000400c000001c130007f40400000300004c0000310000c0010000000000004400400000000000040000c1c000010c3000000104c4000000003004040f00c00040c040100000c0040000004000004fc00000000000c00040000000000000000c007000030030c0000004005003000000000501c00000010040000dc4000000000133014040000c04000000004000000030c0c0033010000004000000303c000000000000000044c004f04cc000000004004053c00c030000c00300304000cc4040030000c0000113c10000c40000000000fc000000cc44040ccc00c4cc0c000005000000004d05c0000040c0000000400000000000fd00000403000cc4000c00110000000000300c4c0040c0004c30c103c000c0c000301000c44400cc000040000c010c04003000000010007044000400c00cc00040000001000000000040000c0000004000110c10c0c000040000000000400000cf30cc4000000000c000004003000c000c0c010000004000030400c000c000c00000000c1cc000000000000030000c40000000000000c000000001000050000000400100c04000cc000000c00310000000040c00000400440c0000004400000004000c00000000040001030040470400010030000c40041010c00400000c0000;
rom_uints[197] = 8192'h30110000001000030f034001c1040c00100031f0010335030004cc00000001000104037d03040000000f000d0d0000cf400c10400007c000300404004d30000000000004300400010000000c040000040000000cc00c000101000c000000c700010000c0010c01000000c0400000310c0300c0000403410007340034f3000300c1000040000001030000000c430c001c300000010000000001000030000403003100c00c33cf0001000000000f0100400107c00000c00d003301330c000000010f4303000c0004000d400c00000004010d040c0fc00010f337c000c300cc000000c001000ccfcc0c000000d100d4000470051d0130000000000c0000000000030004000004cc310000cc04f45c00c3000015cc41c003000000f543c0d4001c0001040000030c0403c001000c000303300cc300003c0300000100330c0100c0000f00070c000f01003700000004000d000407000111c4030007010040300300000400000c00000000000700000c0500c0000030003100031300030000030400c0000304000403000f400c0400310044000c000300000043000000000300000000000103000000000101010c0700000000430c3001333307000000f0100001000d030c110310070101010f00000000100344300000000c440d000c400c300131100004000d0000c3c004004104003c001037001147030001000c0000043373000c00000c400d00300001c040c00045c1c0030cc300f001000c050c1313300000000f030c0d003011c700030c004100c003500004000000004103f0c00404004104030010000c0000000350c03000040301000405300001c3000004030f400043400000000000000100000103c30c0c070000011c0000004100100003c003003000000013000c00cf01000c000c03c00000010414330c40050d400c0000134000c0401c010300030d00300003130f000003c4031000000001000100130c0000000c00040011400000000d00000c000c00030104c30c00000c30cf00050c100001030f00030304000000000c001000d003000034330c030400000040400000434100c0000100100310f00c000003014030030f40100040000c030004100c000000c00101000000001c0c004f03004000c1c3000dc0000cc000000c0003c1030010c004030030000003c0000000cc0500400000034ccdc0010c4104100000030000c0000001c3000f000000010c001100000c00300040001c000040000043004c0030100700070100c0000000100001000d0c03070403000c0c0005000703c300000000010301130d500d00030d400c000c30001300004300300f004c0000000400000000070c0c000000000000003100000c0000c000000303330000405c00330c0004000f00c00000340d00000c45010c0031030000000004400030c30c01010000;
rom_uints[198] = 8192'h10300c000030004c400000003000003004004443c0c0f000c040400000744c000c0544d1cfdc000c1000100300c141d00c030c00c0014440000000ccc00110c0c0000dc000300000c00000f100000d33d000c103100f300c0f00501000c034000104400000c00001000410cc04004010ccc00000300004400dd00444445300c7c0004c000c0000300c10010dd00300d010000000000c0000001000c0100030010000070000cc401000010004d030c0c00031000000c00074000031303c101001d000c00000000c001000100cc00c0000034c410101341110c070110c07d0040cc0d400fc00c3c00010400330c070400001043d40010c00c003c00000c000000c01010041c003c010c0000000030cc007003c000003dc005030400c00040000513430400030100fc0000030044103410c0f0000000030000000003030013d0cc43c0133dc1403c00003f5034030c0000c0d4000d44010f01000000010003cc0000010150031000003c400d0044000504cc007c40c0070000343c00000c0c0010004f4340030000043c0041101100d0140100000c000000000400c0000d04704040d0c000330000100101000004401003070504000f00cf013c040300000c040c70c0000400000000c000400144000c07d01d0000cc013f0000300000cc0c017c0dc0000c0004c400000f11140000003fc0304c0f0c000010400c1003300c00c704c1000700000000000d000500cc30300d700011050003c0034044001c0303000c4040300c34001100d00c047f0010c00037d00000d1030fc00300531000cfcc0c01740330cc00000000cc0cc00f11700c0100c10000c00310000010d400700000331100440000000400144003300000000140cc103000d1c1d000003134300c0500c0300000000c0c0c440100003000030013330040003f003d300000000003013003071d0f334040430d040000000c1d0004004040000404c100373c0c00040303000c00000040700000000000c00c0100c40103c03304004d433c00000dc01400c130000000440077100004c00cc100110c00001404000010c30c0c3f3040000000000010c000cf00010100070007151c0c0d0f003d0300300001d000c000fc0f0000c03f34000013c4004000000101300300cd0c0030014000030515c503050000441007440400041c0c0104c0c00311000000704000c0400000000c0c10001c00004310033c000c7000440000000c0033cc0007c000c4040047000c0f000310100130004000110c030f000f400000100501000000000000ff040144000050c00000c3000c0d0f0000010000007400cf007000000000c00d0000010031c00000c011001400000100010c100100c11000044500030040013004fc0744000000cc004000cc0000010110dc000040cc030003c030000301ff000c0040003100;
rom_uints[199] = 8192'hc300000030040000f03000340000c010043000000000103000c000000000000000000000001000000030000c0c00000c0000501040c4004000c4000040000000004070000010000c00000030400c500000000000c3300c10101001000030c4000c0cc00c0000c00000001000030004700c000000c0c00000040300c0000400f037c0143000100000400000c0c4c00040d0c0000000000c40000434c00f00004c0000404c0000c0cc003001003000c3000000000000400040c013f00c00300030000000003c00000030500cd00000400c00c0103000c40003d4c10031104c00c400000000003004003c404004404cd40000000d0004d00010c004000000000000c30000c000001c000000400015400000c00000400014c0000c4c00c3000040d3044d30000d30100000c0c0c0c00000c01c0000000000c000000044c0000001000070030c00004000044000000000010040040300004130d03010400400400010000000c00000403430405c000033300c000000c0004c30c0100033000000040030400030c030000040300030c01000710000c0001010c0000011000030c00000540c10004000f001000040c000ccd0300010c03000c470001100c3000040013cc030400c00300000000000003000040004010000000c40f000000000c0f0103003000000d0003000d100400040c0c0400000004004300c003000043000141000101000100000003000400070100470010400100030404400c0001040c0f030011cc301100000401000000c0040000000704010004000c03030c430000000c00000401000400000c01c44fcc00c4104334000000000c0000001000c000c0000c000500000c0c000031040f0304c0030000c0010704000003c000000000000040000000400000300c000c0c070000c4000c0150030000004044000c0000040300c30c0000000000040d40410c0cc00103000c000cc000000000c0040400010303040c000000000000030003000000000000c00004c0000304c7000f3000000440450003000030c000000000000404c40100010f4c03040000030000c00001400001000000000510cd10400004c000000000010400040300000000000003c400c5051440000004040cc000c00d0000c00000010c10c000c00100c00c000d0d04d000040000c00000000300001000000d03003c4004000400040103000c00000c0c000000000000000404c3000d04004004c00140011c00011d0001000000040000300005d000000030c10004040007000000000013000007000000000100030000c05c00000400000000000000000004000004000400000110000000000000000003000d0000cc0300000004c300014000000000140004010c000c03c1000000004d0300000000d00c0001044300000004000000040000000004000003000000000;
rom_uints[200] = 8192'h103140000030030003000000000040004400001000304300304030001400c004000500034400000000010030000010000000000dc040544004000000004000003000c030003000000000000000000010003030700c000c303004f03000004000000000000000040c000001003000c00000110000013000000053000010000000330c1500004000000000004040000c0003000000000000c040cf0000000000300000000004000000300014000000007000000000003000004010030c30000000000000000000000000400004400001000000004000010c4300101041000c000300000000300000000030000000d03050c0003000000000000030000c0000000000c00000040000300404000001000070300c30c04000330000c100c00040000310000400000000000040404010001000000000000c0044000000003000d040000000003c0000c00000013014000000c00010000040010040101000000000000000140050000000c000000010000000000000003040c03010003303400000400c0030104005047000000000000c000014000000000000000c00001000301030400000c00100000015003000001000010000000000000000000c000000001000000010001000000c300000000000000000300000100000c0000000004000000c140000000000010040000000001000000104c03000c0400040000000000000010000000031440400003000c0101000000400144000000000000000000000501000000001c000000003000100c0003000000011000000000000000050000000005000000400000000000000c0000000704000400000c000000000d400300000c030040100001000000300000310c0c0013000000000000000c000000000c00000400400c40004040000040000d004301001000c0000004cc033000000000000000000000000001030004000050003c0001000000000000c300440000003003000001030c000100000000c0000c000003000000000003000000073000300300000000000003000300404000010000004003000001000001000000000cc0000c030000310400000400000000003440000000000000030450000000000c0300c00c030d0000000000000000010000100c0c0000030300000700000000f04c0000010004300003400000000000010000003040c000000000000300015400000000000000040c110000010c040000030011c0000001001110030000004c000001300000000000503000003000300100003004010104001070044010010003d00c1000040440000401400000000000000100000000000100000000040000001000000300000000140000000403000000000000000003014000030000c000304f00000000000000000031100000000000c00100000c04000000f0000000c04010003000000;
rom_uints[201] = 8192'h30000000000c000430000000000000040f000004c03030000c130030000400000010000c041300000004000000103030003c00c005001000c000040034000000010c041000000000000001004000c010000c0071001c000400003410003c10100003100034c000000000c00c0c40041c000100001c0134000c50003c4c00000c7cf0150c00c0000000303cd00d300001040c000000043c140c04001000403c1300310030000c0400040010004c0c0000141f000000000000000000000000000c301c10000000040000140000000105350c0c003c00003000000000100c00010430000010000c00004000305130040000300430000010000113003034000004141c0000300030c03000000000010000100301040400000000104000000530007430000000c400300000001010c0100400340010000c0003000000410313501000040cf03400000000000000d4030000004c3000000cc11001c400000010000010044c0000010c3c00000013003004c00000030c000c3000000c0c30001010000c00000100111000000c3000000030110430000000040000000031000030300000410400000030000000000c0c3c0c01313c0010300c1c1104040000014010403f00407000300004c0000000000d0000003cc0000013c0300c00030000cc0000010001040001000f1cc030003401000c001c30000c3c40c3103c000000000035300c0000300401400c103400140c1c000c0c140c000000003015000703cc0000044f0003300c10030400003f004010141000110100000c00101000000c0c00c000000010100010000030001000000110000030000000001110010d000010410c0c0130000303000004001003003000101435333cc0000c3000040037000c00301c000000040000401400040c0050007030000004040c30314c0000000440040c001000300c100400001c3004130300000c00103030300104000010001001300000000001303c00003000100300001000040000100400710000400000000030000dc70000005d1c0004003014400000000000001f0000070401450c04001030000000001030000000dc4d00001300341c1310c01000010000003004000000311c00cd0000004000000c001031003004000400030000030c000430300300000000000400cc000c14000300000c00000000100030000401500030000c300000300c00000c304c0d300001170c300004000c0000c10000100003001403000000003010400004000c003c0404000000000000000c00000c30c030007c0000000034000c0c0c3c04003300300000001430000c3000030c711004cc040c00f0000130303440300dd000000030000d000c0004000001000030000000100c00003000000c00000f00100010000400000c0c003c00000f000040000000003400010000000000;
rom_uints[202] = 8192'h140c00301c040000003c135003000000cc000014300c000c0010031030003000000030000c0c000030001000303030c4cc303100001c000430300000000000000c30001c0000000040000c30013000003c000c30000000003030151000003c0030040c1000000400100c04000c10300000000000000c0430000c00300400003c0c1c03000030000030340000003014140030000000000400300010000010000000001000100400300c0010000104100030000c3000000410001400411010301000000c0000000c3010000010c00010040054300000100c0cf014000000c00000001010000010301000c0000500c1000000010300300000000c0000003000007c3c0d000031003000000110000410001c3c04000c10000c003004003400300010301d0400033000000000000010004c1000000c000c03040034c01dcc1000040030001d13000f30300c001000303034000000343000043010001000301c0000f00030041030001c301c0403000031101004041c001004dc000010011c3c10001000107000000030300c3000001003000003001c0000101540700400100c30000001d0c01400000004300c000c003000040c0000000030300c00000c00cc01c40030010400043000340000141030300000300000003c33103030000000003010101014000000000040143400340030000c103030f003000c00003c0000f40c000c000c0c300004000004003c1000100004000c30003000003c003003300300000010000030300014c000100000750400001c003100100004000001073000000410cc1000000000040000100c0c0044300c0c040410300014140031000c00003c301004000034000000000000000000000034303000300000100010300010000000010100000400000000000010100004044100043403c00030003c0000340c00000c300c000030000030400c401003100010103034003400003000500030001000cc000030000030001300000010000003000000300c000033300c00000010000000000000100000000c3440000030000000001033100c000010003c0430007000000100003c103070050c000c0030100003040c10700000000d5030000004000043010000100410000001300000303000001004d00c10303c001c000400dc04000000003000000000000017100400000c101c000400000000003c040000343030301c1000000000001c0030110000000010100410100400440c0c000c0c00040c000040000000100030040c10040c1030000004000000000011050d000104040010300014000030304400003000001400003000003c003300003000000004330c0004100000100c000000000400010000000000000c003000000cdc30300c001c04003000dc00300014301000000434007004000c0030001c0000100030340030;
rom_uints[203] = 8192'h3300400300ffc00000000300c0000000030100c010000000000c000000000300000300330010000000310003003000400000010000c300100000000000000004030171070000000300004000030010000700000033711000010000000033140000010103300300030000100300f00cc000110100c00000010103730001310030130300000000000000400000000000000001000000030000030003001f003000431003000000010003030000f50000c00000000100030010110000500010000000110000030001c0030100001300400310010003000400001001030003c100000300000000030000001000030040000000000003300100000300003000000007000003010700000144c0030010000003001100000000000003000000003033c000013000010000030000001000000000010103011000001000000001000000030100030c00000300030301000003100040030000000000131000f000030000c1030000003133c330431100000030000030000303000000001c0703000100014000010001300000110300000000005300c00000000000000001000040000000000107000000030000000031010001103000000000001103030000000000c300300133000070000000004000000010000010000100000040030103000400000000003000030010c01000000c0000000000000040c000000143310400000000100000030001f0400000030000300103700c10000000010010030000010000f000031301001043100010001003010000030000010000030000c00004300311000003030010000000000000430003003003000003000000030000001500000103001000100303c170000301330000000000000300004001000000003001001001000000c00300300000000301010000000001300401010000300300300000704300000043000003040100c0000000010000400003303001000000010003000000000003300003000000010000300000010003000003003d43f000000001000117300c010000000313000100310010001000130010000d30030000300004000001000103000000330000c0030000000000000040000000400013000040031000000f10030300000000000010000100000000000003000000333100100001001103c0000000000140000103030003300c400000010700c003c1010057010103031c0340c00300000300000331100000310000000000c013131100001010000103401000010040000000010003000000033031070401010030300000c01010000001003310030303c00100030300000000001301003300000000000000001300030010013001c10000000c330000c00300000300000001000000000303130003010101000300000003030100c0000003100301000031004000004043003001c000000000;
rom_uints[204] = 8192'hc00004003000000040000c0000000c30000c0000c0c030000450030003340c0400404011000004c0300c00c000c000000000dc030014040000044c0000c04000cc33c004c00cc0c0000330000100c0000000100d00c000c411040c0cc00010001400043000f0000410100000c00300310000043700303001dc0400c7530004003000000000044103300000c0010000004400400000000c000f00401400300000f000401c00c0400c0004033ccc00c003400000000000c300000c00040400000050000000110000100c0010c00c1030c440303000c0000000c0c30040c00040001000000000300000c00c0001f030040400100c30300400c704000c0000000c0c30000c300c000c00001c0c1000c010433f00700400c00c4100000ccc30c4100c3330004c70000010c0d404430f40c534040043010000000000c40030c01c000010c444000040000c134f10300030010c0000003c301450000cc0000cc40c00045004000c0004000030435044f300c0c13c0c00d004000c00d33003000000c0300c0400cc000000310000c03000004010001000000fc0044010cc000010004050c010c00c1c00013301440044000c003004410004dc01110004c0000c010c0330cc04030c3000000c04000440000000c000000ccf3d3c040c4000000005dfd010c0000000031411c0000c00430c000c0050400c430d00377000000430c40034040c0c00000000001000400174d03010001000140101300c00010000330031000400110000cc04c00c0c0000300004000d10c100c4c030c000c03074000cc00000000000040000303034f0c0c0000001000d00010001c000000400307d00c310000004503000000000001f4f500c0000d0300cc0003004000000000414040334000400000400c010000c0300f000000c30003000005034000100000103001c033c00c03000040310004700c10c010f403010040000000000c0c040443030044cd000c001400c0071140000300700c0000d31c300010010703000000c3010103000011010c000000c0070001400c0001d000404500000000000003c000c07000c0000000f010010000004000000440c000c00000c0c0000000c30045c00f040c000c0043035001434c075f000000000003004010004c43001000450c440f003300c5004440004014c001030000000000304c00f3404005034c1441000004040c00010000000100c000000300300300000010c000050010110c4c03700f0100c00000c43100000003004100c000010001010000000001c4003f00cc01c047000c310c0001cc730500040003000301010300f001fdc0005001004000004003401300000c04000cd04000c000000000300030000000300000c000010047c0041d331000000400030010004c000003c040000f0000000300f0d0cc0c000300004101;
rom_uints[205] = 8192'h1101000000300100c0c40340110001000001001001cc3000004304110000ccc00000100503c0c000400f0000714003000c30005d4014401f103c000000000000004c00f0d030005100000c01d00040400000007cc440010ff1403c00000c0c3000411000000543000000000104040070000100000300033300d04c0013404000ccc0433001000004003c00005000000400c400300013c1001cc0070000f30005031330000010030330000000d30130c05110f000000c114000c100300c00030c40410000010340000103c0d000407000001104c0033cc400d0d1d0000013000010000000f00d100000fc010100fc100000333d40100000030000001d43000051d00000c400011104000100104f0d400000030c0f03003100c3013000000300c003000000003c030300051c010000000030013103050350004100cc410011400000c0030001010000c0000c5c130c1001030010010050404050100400000c3303000040001013f30000ccc4c1c000140c00c0017c000033000331c0000000010040001301500300000033000010005313001004000004450005004153000300000c70cc0c010300000031340000050340ff00000f40041c333031010030000cf3100010005000005c00030030004110000f3040003d403370010000000333c30c4010010c00440500031003000000003c13000d0037003100040000010cc00001d0cc00031053000001c000300041c350530d3100140d0f00003000405500cc00cf0c00c030010000000010001c304300300004000c4d4d0030000003070040030c30c010010000000033000000004000000c00030c000c40100c1133c10300001013503010000010004dc450313403000100000000000000f007040c0034010c00ccd300000001c40000001114000101430000000104000000003000504c403c0000010300d0000110f11101c5c0000330040100104100100000400c1103c004cfc00001c0000000110000c000100001301000000701c1003c03004101cf4c10050000300d404000c014d010c3500000030344400030000000003000011000004d30300033030d0111c003c300c003000500000000001c30000c010434013c0c001d1000f30000cc113000010040000f03003d33000130011030100dc0000030033000013c4100c030303041703003014033d000000444000c000500f0c0343000110cc00010000007d00000030040000000000f01000030003c00d5000c0c3330c047400cc000000000c0f3c011077155040000000000000400011c50004000430d015003000c0100000c0004014015007c100000001fc0c000c00000300000004450030c07000c0000003000c300001c0003c0c0dd0000100004001d0c0000000040033040101033033330400300400040000d010000000d00300101100100;
rom_uints[206] = 8192'hc00000c000000000000100000000000c104000c00000003cd00004101000400030d0c0f00cc03000001000004001c004000401f04040000c300400400000c00000c0c0000000000000c43004443040c0000c00300000c0c000c04430301001000000001000100000c000c00000c00c000000000000000000000000000004c000000000000c0000000c0c00003010003000000434304340c00050000010c000000000000100c00000001000400430000c0000000c44000000c010c000000000000100c00000c01030003000354c144030100000c0c00030000070c4000000700010c000100000000000000004c000c00010400000000033003000000000047000000000c000503f0000c0341000000430c4c030cc001010300c00400000404400400110100000000c40c000004cc00c000000c40c00001010c000c0100000c00030c00010c00100000000000c40043000300c100000c0004044000044300000004000003000001000c010c04c00300300000c004c0c000c1000c0000000300000004000c0000440001000000030001000000000000400c0000430300000040550c000000c000000040c004f0c003000000000f0003c10001000000004c00030300c400000001040c000030004cc1000cc000000c0fc100000f000fcccc00001c044d000f0400c400000400000043030000430300001400000c000000000c0d0007cc0c0f000001000c000cc100030300c00000004000040d400000c0000000c0040000f0c0140000430040000000015d04000000000000c0000010000c1000000cc0400c0d0000400701470000004c000000000103000373010c0000403d040000000000004000000004000014c00d00c30000c00000303300000cc00c0000c403030003000000000dc0000040c0c30c040303c4040c000000000001000040040c100c0030c50000000cc040013310cc000040010c00000003000d0300015f030000c00000010000030000000000404000f10041040c0c00c00c0c4004000000005307000000000000000040010c030000c000400c0000000000000c0c00000040000010c0c000c000030cc100000010000c0c004c000044310c030c00001c0000000c0000c0000300010001000000400c0000c3c000000000000000c40040c003010000030000c0dc0030000000030000c100430000407400000c00c10000010d040000000400010d0c40000040001000001000040043410000010104100003010000400000000c0000004c0301040cc000000401010500c00001040000000300004300000000000000400c040d00030400000007000000000040030c000004dc0300c44d040000030c0540000000c00040004004000c00000c0400000f00300000000000c00c04400c00000501300004000d00010c0000c04005000000;
rom_uints[207] = 8192'h5c004000304404003030340000000c103000c00400040c030000300c00044314000004f030040000100c0003300400140000040303300c3c0c001001140070f000000004144404000000301004100c1400000000340d170040003c0c00041c0c000c0000000001100f00cc0000c11030d4000c001c0c041c000c0410000d0010000444c00010000c040000010000003000030000003010c4011c003400c0000400400000001030cf44000000000000000010300000c000000c0c10000004403c1000300000000030f03c040000014414000cd70d00001300500000054d00000f00000c0000000c0c30110074003000000471030410000000c10000000d0000040400000000141000001000453000c00c0110500c304010300c00001c14c70500000000001c30033000000c0c301004000c000004cc000c00100c000330003c0407000100c00000000c070004c300001c000000440031075c143c0000c0000c0d0044044001f0f4000400040cf000003c0001010cc000001c000c5c0c000000000430003c140c413000100004000001003c0c0300170000000000000c000410000410c00c10070400040000000c0f3410000040001c410300000000000004cc00c30c0000c010300000340c0c1000000f1100003c1010003000001400100000000c000c4f0c00143d0cdf3403c40000f401004037040c000c300700000003400c1330340040304c5007000000001c0400000000005c0c44000000000c00013000f00030040000000400c000000000000c3130400000c0c004c034000c4c0000100c1034003c040010100414030400400c0400040004300c000c4000000000035014004000141400040000030df4030400040c0c003041c004340c000c00501310400c0c04001000c300000c0c1c00000004040410003c300400c00004d0004c3401c44c045004000c4c3c140c00101c1c030100100c0c3004000044000400f0000417c4100c0000000c0000003c0c0c1c00070dc70000c0003c0c0004c400c01c140000300400000004cfc40000140000004003c00030000c0100171c0003000000003400003100cc0d000c35005030040400000c0414000400c010000014fc000c0000c00004000c00f1004c00000400000000f0000d3c00003c00d00c00c0004134340000003c001c070c304c0000103030400c0cc000c410000c0c04000000000c00041004000004100c0030000c1400000c341c0001000c0000100d03000c3017001400001c50000030040c3c0004000c4c00113100000000140c0010000d3c000010301cd40c0440044c300c30100c340c0404000c00000010000c000c0000cc503c041000000000c40000000000000c0c040010001000f01400104c00000c001000140000400c0d3010400c1c000400000000100431c40141030c00003c;
rom_uints[208] = 8192'h4100000004000c0504030000040f35010f000113040f44000100040011330003001c030f00000005000100f10001003300040034000f01030403004c0401000f0c00150f0003434c00000c054400c00f040c44044f40000405c50f0c0130dc0400c4150004000005000fcc0c0c00054000c00404000c07c40c010d470550440100041c00000f00040400001000040003010100000010400533051f000c0c0100304f000507141005000d00444000000f00043004000c01c30104010f00030c4f30cf03c0c00004043fc7000f0c00cc000301f140000fc0410c0c01000c4003c50cc1000005003500000c0c070cd304410004000c05050c0001010105000c00000f000c0503c505441c0d00100f0c014f0f0300104c00000003000030c4040003004c0300000000030c4431030000000c0d000c0000000000010043c50f000c00c10007040501f0044000041c030dff00cf000000000014000c0007040c0c030500003300c0400c4d0f00010101070f00000400000d000f100f0d0c000c400c0004030304400001040c37004f004ccc1000010c0400000c30050d115000010404404c0f173000c0c50000000141f50f0003c0000f010fdf0c00000500000c47340541c00c050d350c04040000c00400010d0c000001001431040c000130040001400004c1301c010300050f04140107cf000004f30fc00d000400000c040000cd00000f04114c3c010000c000000100010c01000c05001f01c00400040000c30f00400cf1c011000f000c001c030000004c141304030c0504044f0504130c0c0f7c0c00000c010305300f000c03130030414c33070ff0000300030104d500043c0004000c140000010030030000c40f101501050c0400000f0f4001011c04000c0cc10f000000001501033c0140034005c3040405003400c300050304150c00030c00010c0c0110000c070c00050f3c00c00f0404010403000d0d0fc10300030c00000f0104003004703000030f110c0103cc030c040c01000c410000030f0d0105000c0f03cc0c110005001c07df0000041f0f00004f0500430cc301cd050c0101031305000c00114100000f00470f00c40f000100010d04041c000303043c0005310135030304050007070503c40104040403c30030040100300fcf040c05350c0f3c050001000c040033c004cf1f03003f00040f4c04470c00040403070104100cc0cf034004041700040f03003003041005cf3c0100301c0c0104000100000c000105000005040100001f010c01c40513040300030c0000030000000730303c01014c10040f01c003000c040000040c0f0100c3000000c00031000c030400001041000001c0010c0f10f04c1300c001004100050c0535010f0c01c0000c00400c0103000c001300000f000f4301050f0005000000040f00000c0004040000;
rom_uints[209] = 8192'h33030000000c000710030300c000000f001004000d300000000431000411000003330d01030c0000300000f0cc04440c300140000301070001010000070000c00300143c040c00c4000030034c0400003010100d0d0300010c3070c3034c00000014103730300c004c34013000001000100f11343d0000000004030400140c34f300f000000f000001010000040000100005000000000c17000700113410c100000c00003003000c000f0400403000cf04d00c0000000304110000400000000000d73300000011400101c0040400c00700c0c400000000fc004300000010000000c0000300001c0000c0000007430c00017d000300c0000000000003030000000c4330147c0000100c40070001003000000d0c0000033f00030d3100043f371100500000330d0404030000f031000d40000c04000000030000004c0000140000040440000004000030000007100000000000330c00cc04c0140c00400003001c033041003f010c0103011004010c00100000000000000300c1f0010000100c0c000fcc0d301000013c01300400000001f000040c04000500140030030000110341f330010330030000000c00000301003c01043000513f34001101343440001000040004000c3000001030040400040110300c0004040137010300000ccc5000070000f40004040f04c0100000100c0c0003000c0c0000010c040000314440000130c11c001301330005000000030c0000040100110003040400c400c0000f30010c0433040100000010001040004000030043333300040c0000cc0f10000403300401110000000c3000000030c00700303040000403cf00000c000c00000c30074c0003130300370503141003000000041c3c00010044070cc41000150005c071050001003004d0340d003434c0301100310000c30000c000000103c00430003000330c300000000c000f0405040000300004001000301700040f4000000c000000100000000031000300000001030f000c010d0c3304340c300104000133300000c0040000000400110010001f030400040ccd03001100010c000300d0010430400330330000fc010000010000000434c400030004030000c0031040003c00c044370c3c0f000c000d00000145000300043c0000f10c000c00150c05000430003300140c040100000100000330010001cc000df040040fc01c110300f00100300403000000000300000000410000cc00c0003304013f30070100150004040331000f010000000c3401000c0f0010000403010c300100000c00410400100300400330000d1d0000c00000040000040d000010000010c1030c103000f00c001c001007f130040f30300300000010000030000401003300000404340103011d0c030004100000001401000c00100010030d1000000000110c0f04010101000007;
rom_uints[210] = 8192'hd000c000000000c0400000c1100000c470c0005000c00c04c001304000104000410003f00000000000c04000c0c3000030000000c000005c000c000400000000300001c00c11041cc00000004030105000000000c0c003003070300040005000cc4000300000003010f44000000c04c00000300000c05c300000c0c07030c4340dc0040054d000cc0010030410c010003400000000000100c03030003c00010004040000004000c0303300f00440301000c43cc0000000400040000000f03030c1500100000cc0f4f01000500010500004400000034001c0414011500410000000c00c0004000000300000100f100000303f4100f040000030c0c014000000c01000300430fcf00041007000000010c13344330135c430cc0010c043100000400740000c030040c11540000000030000c0000d00c010000040c0c000c05040cc34d04c00370cc0c0000030404000004000500034005c0030500010000010003010f0f000304c03f0c000400003400040000400003040c0000000000cd101d500300000000000f00000c00000c0000450400000004100d000c130005400000004300010003000107000300034300030000000000110c010cc100cc00010504000c010103030c00700c000c0000004400431c00000c00010000030d001c4414350001070110c40003000c04c100300100050000000000c307010c0c0400c000000103c00f00444000000c040c0500100000030c400400010c0100f03145030000004f03000c00030000340c040000000041c0010000030000011cf000000010001c00000000cc00030001c00f04011c030c30040d30030100400000000400430310030c000510003134000044cf0004c00d0010010700000000000c0000cc000400300000001c0f000300300001110004140010c010030010300c100003000c00330f00100304c3040000100300300300100c000c40c00f04030c00cf0c0300000101030000000c0c340700340000070c00100304000004c00c433c0cc000000000001d5c01030030000f34c1000100000040010f0041c0030c000004000c00000c0000000003c0c0000000010c000f01030000431f00040c0305074c001c30000000000c31c000000f40000c000c004000000c04000f00004c0404c00f03040031ccc0004001000f0c0003000c005400c403030004010301050430000c300310000404050001010500000000000000100300c400030000c001000000000f0c000c0111cc0300000043000041000400100401057110400000000c053010c0045007434314040c04430000000004100013003004000c000001000003004f000000000010370003401c0001010100f00c0000000700000000110000000004004000400000030f0c000d0340410d0005000c01000400030000400100030000000000;
rom_uints[211] = 8192'h30f000000030101350000054c000f040303010040c70000000000000c03030101010300000f04000001000000000503000f4300003300c3000300003700000000000004040f30004100140043011013000c00040f07000000300d000300030003010001040000000c000030cc04c101041130d103330003000003000c01000043001400000040000000000000041000000c0c000003000003000000c4050c03001004030d040130010000001d04004c04333c0000000000cf0000014303000303cc03000000003001130001000000050000000c000301000301010c3c5c0304050f000500013301001d0004000107000000000130500003400001050000000413d000c10f000140c50100030001000000110010040f0300f00700030710050030100300310f00110d0045f0c000133c01000100011ff000010c00330c00000401000c01000013030f07000405030300074043370c031300100c1013000000030000030307000105011033310c0f00c100000c1000050100400f30004f30000f4f014f0310000003040c0c103100040000000000100001000c000000000140003301400f0100040000040f330c0df000030c01000f04170000050c0100130f30033000000303001704c401003010000c4f043000000350010300010301000c0c000003000010000f0303114304070000030000000f000c3000070f03030110010130c40005040c0300010030100c000400000f00000010050000310c01300f0000313500071f0403000515000700003300130c0001000304033003000000000c00103300c00000000017030000050300000c0104003303000007010300010f4f1d300300033400050003000000000701401f0f0003003d010000400310000d030c00c1030400010000100001110c0000300300030000130100030003c3010f050000003000000300030303013d04010fc3010030004003013041030453000501030003000000030404000000000c300c000003040310000003133300000000000000000313030031000d0004014000031000310001000100011c0401000c030330001700000001073000030005300003c100300c47010000000144000403000001400403540000000003001c130445070f04300100300f00000c00030c00000010050030040000310134300001000d0303303400c00330101003000030000c001000000504010041010003000130001400104010310f0103040c000d7304400000000300010001004300004331000103c100330001100400030f0000003300000c0100c1040004303000c004000c0030000c01303700cf000000000000100f0c00010c1cc30007003404001f3c000001000cc003000000330101310004000003df3000004000030000001300000030000c0c0000000340004001030000000000;
rom_uints[212] = 8192'h10001000cc000400040004c040400c0000000000000013000043030030004404003c35340c0000004004000000004100130000f000100c0400130030340000140030f0000000300000000300003c3c01000010c4031000c03300033500000c0ccc0040c3003c0400140c000f3004c4000430000000000405001001001000310010f003001000003c000000000034000000400000000000f0000000000000c000000000000001400c000010000c050004003010c00000040cc000001404000000c03c001000000000000000000c000000344c000100d0f03c053031003f3c000c30000000310c0404000000010c0300410410303400000400003000350c00040005cc0404000000030030f0001030000c0c000000101c0c003c140c3010040010000040003100001030c410000001f004000c0030000c0c000030100000100034300c00334000040010000c3004000000100010000004c003001cf010cc305000000c00001c043c04000034000c0c043c14040cc40040100000000c0000000c003cc00c04000c000034000000c0041030000000300000000030030004000c00001fc00410c40004310033000c0031171100000c00f00300000001300003001300c05c10300001000430f030100000000d003000000c0034ff040cf400c134d010c00000000f00300cc040000400010003c00c0010001c0c10103000140c001030000000f004000000000c0000330000300401000004000440000030000000100050033000000000100000300400c000040fcc140000000000300005c01000043d0c3000053000040c0000000040000c0c00041404004030000430000c30100c4c0004003cf0040004000000010c00040004003c00103000c0400c0c0010000000000c0400000000c000130c30c03d1030340c000400ccd0040000f00014000c0c100010000c0000300000044000000410df040300c0000000000010340c00040000000000000004030c1000040c0000300030100000c00100c00c00300000001034000040000c00300000000c0c4400100c0000000000040000c00000000000000c03c000ff0044c0100000400000000030003000003000c000340c00f00400007431000010001c3d0300140000000c0000000000001000000000000040100c004d040040000c000000340300000000000000003004100034430c04300400000c040cc04cc000040070f00000000043040c00f10300000c005040000400cc00001c35f1000400300050040000040c303001100040100c0400100005403440000013000c070400c000300030003030101300ff3104040000000000000010043c003035c40c0000000000040000000000310000cc000c00000100430000001000041000000030310030031c100013000500300c00000000004c0004c00000004000;
rom_uints[213] = 8192'h4000000000410340c0000003004100c1144300cc000010000d000000030000000100c7000d00c0010300c40d000405c00030100c01c00030000000000000c10000c101040000000000070cc0c00c010040404440f1000c4ccc0400c00c01000004c0400f0000c0000044000301c00c0003c0000101030000051c00c100000000440003000140050044000001000000004040000003c000000000c0440c00d10301c0030004c300000004404010c00000000c400000c000000c0004c0000000c000c10140ccc00000c00000010004040304030000000c4c0000c1000c00400040c00000040c0000000734041000c0004000133100430000000000030000000c0003000000100c04c1c00c01c0c001000cc4040041cc004ccc00001300400004c0c000000cf00000d0000404c000400000000000c000000000004010000000c1c4004000c003014001000400c10c010300044401c0400d0701c0c0c30d003100000300050755003040000004000cd100000000cd4100030707000010c0f1000500404000400000000000404004c00105044304000000c0130040c004c00300004055040000004400c0000000400304d0000c00044c0011004f430003000014004c0403c0000c0003c000000001000010004100000cc30c50000cc000000100007001d00d00000001cc0043c00d04000001cc04000000000500004000000c00c030000c0000c01010000000004c0d040000040000004000c3004303030040000000010033c0c000000000c00001d00400034c401000050f000140c041c00000c0c0000001c30cc00000000d00040400100c00044000000d000001004001000c400003c10001c100000005400500400000033000010c40000004050000030000010cc00000000003c00101400000cc0010000144cc0000001d000c3cc00c7100c00000000c00c0000041000100000c044403000003000000040001050000c004c00c0040000000000003c1000c00000000c001c10040000c00c3034000c0cc00000000010040010ccc00030034c0c0c0300c010d03f00140c00000000001cc41c0004000040041030000130001c00000cc00000000000000100c00c301040000c43f001000040c4047000d0000000004000000000000050000040c4005c3440033030000c0400000000000cdc000040d0100c00000000c400040cc00000c40000100000000c003400300c0030000c00d4000000cc001c3010004000000000cc00c01c0403040000d000c4100c44000000c03400c10f004000000c0c0c004c44001000c00000000000000c0004c00c00000030000c400400c00700003000040034000004001000c00000100000c00000000000000000004c0013400000004000001000cc0010000c00103010140000d000c000000010400000c03004100004000000;
rom_uints[214] = 8192'h501000c4003000100000010000011300c000000000003004030000300040000043310101401000010041401001130000300330c0000040007000003000400000001030100000c000005050001c003000400033100000001000010000000303c300000030030000000070001003f010000000f0030000f03040c00001100100103000000000004001000100400000c0000000500030000000c0000001101000113000f0c03010004030010010000300c00000000011301033000001100010000001004000007040000000f000300000503300f0c04000c3400000330c100101f1100000103010000010000000c00000010310101000004000000000c00003003031301040004000530000000100c413003040000070700050410030c300000440100000003301040001c10001000040401000c0000010300000030010040313000000300003000303d040d0f0004040300001003033037030030340f01000c0100000414041300410c05140307000000030000011000003130000301010c030300000310001003033c03031010001004000403300034000c000010147100000413070404001303000000040000000331000310300403013000000100040f30010000141c000100001313000700103c0000040000c003030001040c033430110000000004300000000c01000004000100000003000c30000c000000033304003300030004101030000014003c0404030030300400100f301c0000310000c400001001f003300000000c0c00000300000001170c00100001000500030c000c0000040000010100030001000c001c0001000007100700000c0313010004030f04004007053f00000d0100030000000000000000013000001000000101300030001400003003003dc003003001000001000003450030310004003100000f0000000013050c04051030300017000030030730010100000030000d004001310000300c00000000000000000030300103000000000304000000000004003001000c030000110000000c00000c0100130f00000000031f1000010010003000040003000000030000001000000100010000000c033001004000003c000100030c000c330f0c000c0000000401003403030c00000300140c000100000730001000040000101c0000100c000004003c00040300000001000103000003003c4c00000700100031000000000000300003000000000030031f3014030000050500300401110c000f130c1400000000000c00000100043c03033f0431000004003400030000040700050000010000103000010100010700000f110000330000000100033f0300001c17700500c703040c000400300000070c000000000f3000000104040000070000340033000000000001000004000030000c0400050c03031d0400000c1010;
rom_uints[215] = 8192'h70cc004040c00070300000000000004c000000400000000000004c000000300000c0c04c00040000c0700400030000cc3010c050c00041010040000000304000000000d00000000000001000400010004004000400c0f040000300004000c4000c4000404100000c3000c0000040004c00000c0100000400000d0000000c0040f000d3000000000000c000004000c000000000430000c040c000000000701c1000000c0c0c00001c00c0400040c400f004c000000070000040000c000c004000400000c0000000000cc400000000c470300000c04040030004c00400004c004cc040000000040c004c0c00c40fc4c40007d44c00400000000000c00000000004f400c000c00c0c1000c000c0504000c000040c0000400000000010c000300000000001000000300000000003004cc4000000000c0c0000c00040000c00f000c04040007c0040f400c0004c13c000000000000cc00011001cc41000450000c4004010000011c4c000000000001c10003000000000000040000040000cc0000c000c0004010030c000c0f400c000c000c0000004c0000000400003400000300040500cc00000300000c00c0040004c17c0010000430014c04000000f4040c405c00000004004c000000c04c00c00000400050000d40400c04c000cc0000410440400c040000000400040c01000044000c00100ccc010000031040004c0000040c0030004400c0400400040c4000404000040000c0000000500000000c040000400000c00000c00c000000c00c000003400000000000c0000004000c0c30000c0400040d0c00030070000000040c004000c0040c000c40cc5c000c4000c04000000000c0000f00c00c0400000040c00c4004c00000004000300c0004000500040c40000f40000000c001000040030c0000004040c00c00004000010d000c400003030400000030400000440dc0c0343001000c040034c000030c000c00c00000000c4001010000000000cc0c01430000100c000c410030000c000000000000000010f000000c0c0000000000000c000000c000004030100000000000001400cc0004c000000c00000cc0040000400004000c0000c000040400000000c0000cc000000c0000000c000400c10c040c400cc0c05400000300c0000034c00c0000f4000000000403c4c000030030c000cc004000030400000110000000cf00000100300c040433000c000100f040c00040000000c0000004004cd00400c00030033cc0004c0010c0000c000430000000000c050000c0040000040000400000003000000100001c0c5001040000040000030000000c4c0000000000000000000c0c0000000c343c00040000100040004434000001c00400c0000003c00014003004cc404004040040c00040c5004403004100000c4c000000000c00cc0000c000c000040;
rom_uints[216] = 8192'hc0cc00000003c0000f000000c30c0c4cc00043000000000004c000000c0301010f53030000400c0000004300cc00070000000cc1040040004f000000050004400c000f0000030700000000c0c000400c0c00cc03c00004040c070000c40040c00c00c0000100000000000c00030d0000c30004000000014300cd0c0000010000cfc4410000c0030000c0010303000000000c000000000000010300000001400400c0030c0000010000070c0c074007c1000500000000000400000005001400000c00000c0000010003440000c403cc00c1014004c100040000030c000f00000004000c040cc500040f0003400040010c00400340000000000004004000000100c40000000c040304000004400000000007c00147400c000c04100c074100000c000fc0000000c40c00000c0000004104ccc004c0c00c0f0d0d0403000c00040c00c7000c0f0000000c000300c00000044d00000c000c40031000c10000000000000007cc0f000000000d00400000040504030100000000034d0c0c000401030000c00003004000030000000404000c40000f00000003010c41000000000f0c000054010c0000000004c0c4004c440000000001cd0f000504410c000c0100c30f07040c00010700000004030c000101030000044401cc000c0f0005000000040400c10104000c00050d03410000000303c000000f00c00f0c00050c004000004c0403010f00000c000cc000cc01000c03004c05c0000000030044030001400040c0c400030cc404000007c0000c000100014400030003c0000300000000000d000c4000010000000003004504000c030004044003c00000000300000c054400c30c000c00000001000000000004000000440003000f04000003400003004040000dc3040000c000000003000000c0c0030000014003040000000c000d0c0000044000cf0000000c000c0c0000c00403450c0000030c0303040003000c04000040400d000000000004c0000700c300050007070c0000000c00000001000045110c00000703030004040c4003030c0c00000700000004040c030c0100cc410c000100000004074c0d05cc0043000d0300030d00000000000cc4440000040000000d000003000000c0000000c00001400007000c040403400040000043000004cd0300034c00030100000c0c0c0c0c000000c40d00000000c403000c0004c00100004004010c0100000c0c0c0000000000040001004400c00407cc000c430100010704000100c005000000000004cc000d00030503c0c300c0000000004c0004000fc0c0000cc10140c04c000c00000c0c000f000c0fc00040000c00000003004100000dc040044d000400000c000000000c0f04000003040c00070c0c0c030c0d000f010407000001c0040001070c010101cc00c0000000c40314040d010000000;
rom_uints[217] = 8192'h5010c000300000030000000cc0c00000300004000c10c00000c00010000000404110333030000000000070301000043000c41400c4703000304000c030000000000000c070100100100110140004cc00000030c470d004040c30f00c040cc000300c004070030030003000307700c40110003400000040100f3000c10cc0dc0014340c0000000d04001000000030c01000c000300044103c3000f04030c0000000c4c0000cc0cc00dc000000001000100010f0000000c0d0000000100403c000104030c0000cc0100404000400c04004540070014044000cc040f00014f04000700000031000000004440010043400c01410300cc00000300000000c0000004300400000131030cc0000000000000004f0004c000c00503c700040c040c000014000300004400000c0010c440034c04000c00030c01070c1000000004030c00110101000c000000000047000100c000000001c0000303c05c00440400440c0c00000340d104400c100c00c0030503c0000107cd0f00000100c014304c00400c300c0070c0cc010340000000c30cc30f0c00c30110004400c40f0003c00000031500110dc0c00c0c000030000105000d01000c040004c4004d014c000003c001c0015400c00000000303000000000101c1000340000000370030000001c000000000c0000701010c300d034003040003fc00000d3000430c400000000003003f0400470403d003c400000d0040c1000005000000400c000070000ccc030340030143000000050000000000003300c1c0000101000cc0000000000000410005040001030c003341000000000045040003000103000103400dc0d4030c000d01f0000f000500000004000f00000c700130430c0c01034cc7d00000cdc0000c000000c10140040000000dc3070300014400010c40310c000515003300000d0f0404010000010304000c100403000004000004c07c4301010303440f4033000000030001000c00000000000c0000030001cc4000000400cc000030000003440303400c000c000100300c100c0f474700000000030c5003004c0073010000c301c00000440005400cc13000000c000001000c430103f000c000000f000000070f00000c1d000c000044c1044c000300000500000031030000000c533c000100c0070033000003004001c0c0370004c4400000040fc30000400000130071003c000000010301000503000c43cd000430000004000040c4c300030c00000043047f00004400d00c04005c000400000000c0c01401004407000000004001c1c3d0000101000000c04c41c7000000040000000043000100040000300005000000004100030000000f003707c344000000040c000c04000f5040c1000c0000400300300c010100000f03c100fc001101c0040001000501400000404c03c0c03007400000c0;
rom_uints[218] = 8192'h4d000100cc1c010100004c4000001c01c0c1011403c01d00004040030300404003c30c0c00f1000303100c0004030cc03003000117c1003100400c01cc010100c000330004000041000001c100000003cc00111035110000c00f00000010c3000330030100000000c107000300330000c0300040000340000054c13c41000c00410c000041004000000104000400000c001000000000004340004000340003f001100000030c00cc0040000c100c000000004100000c00400000000000c00040000100010000404301000001010071c0010043010100030103300000011100030100000f0000c3010c00004d0c01010000343300030000000300010300000000400410000000310c330000c100330000004100030003000003400000000d700040004c0000c00000011d000000000305000003030c003500000000c301044003030004c0c30300004540c030000050034003c100004c0700c101000700c00003013400011f010000c1ccc000c00000010c00000c00000000011000000000c101000101c303c0000000c40000011000030001c4301000010c0340010100403700100d0000cc0504400000000103cf7c000000000000c30003c1c0f00003044c00001501c30000f00d331001000300030104000040030dc30300c300000000003000011003c10c004c0400010400000001010000000300c50d01000300cc0300400304407000010007300003ccc004010141030010c000100000c401010c003100010c0000040001110000310c1c00100003130700000101cf030411430000010300401011c3004c000000007000000000000110000400000144000003c3400047010d000034010c00030c03c0c70f000c00010c0003d0400033c1c400070c030000004000300000f107400001400041c334c701c01c3000300003000040000000030c040030c4c3cc010301030003001000000f000000010c00000000004000030010040000000000010403c001030100003404303003000311130033c3130104c00000c001003100000003310130c003000011310040300000010700034103000c30000000003c004000000301000000100333000100010c033fc03000010c044401000d1000110000400001134301000400c0000071000001df030001010000133000c301000300000c00c0000000030041030c41000001c0c30303000133c110004000c000000f000000c10c4000cc001d000401311300c000000374014100410c40030300c3000300300300c0010f00110c30010030000007c0030cc00001100011001000330000c0300f030140000003000000000000000003001c01c000010100030007400d050107130100000000005c0000c000c00100000c031000c0110003000044043000411df11000030004010030c1c50c000000033c0c000330;
rom_uints[219] = 8192'h1034000001000000c1000000400000000000000100f000000100100000c00030004100c03030000000000000100001000000004c30c01000100000000000c00300c100300040000000001004c100003000300300410030101000c0c00000001f0041003010000000000000000000c30503001000000f000000cc000010310000d000000000100040000003000000000100000000003000100003000001003000000000c30010000300000000000001000000c30000000100000c0030000000000000003301000000000010300000440d00000040000f00d003c0003c030000000000000000100000010000f0300303400000104000030000000000000000000d0000033000105300c0000000100000c0300000000000c00003000040000001410000500040d00030000000110c004003030000000000110000003003010f1030c001000030014300c000c004d30000000300000000000c03000001000001001000001050f000300030c0000100c0c0000000000010030000300c100000031400000440000000000030300000000000c00000000000004c030000000000000000c00000000000004300000400000000000000010104cc003143000010c0010000c0404000c00000d000000000100000000100000300c00300000130403300104100033000c000004000000100001003001000003300000300110000001300c000c0000c00100000c004c0304000000000c010030000000000000010440040030001000000030041000000300001000000000333000000100100110300c1000300000100000400000300000003400000010050000000034000c00000c000000300011000101000000100010000004000c010030031000000003040300000010000000000000000c000030010f101004100fccf30030000000000000000c0005000033030004004000c1340300000c01000000040000000c03010000000031000100000c000000030100003004000000300000000000030c0c0103013d0000011003000000070001003000330501300000000c300c00000000000003c000100000000010000010000c0000040010000000000c000000000000000010000000010000000001030000000010100000000000000001010003001000000000100030000500000000150000000c040010001300003030000003100400000000000100000300000000000000000001300000000000010004000c000107100000000d3100000303000c00000000000040100001100000340003001f00040407000000000000100001c413000000000000170000100003000007100f0000000d000000010304001c01000c0c1103000304000f00030c0010000000000300300300100103030001000000040000c5101000000000000000000000300000300001030c3000000;
rom_uints[220] = 8192'hc14310c0003301000401000000003341f000000404cf01001c1000100100000030c3003c0013000000040030100047c1000000cc40330cd371030010c300d000030003d30310003110000c14c0003300310001001040330400d0101103df00000004040c300000001000c00300000040030400430f430f1000c10100c04100100cc073010014004040100043c130c000003000000033000030000c404013010010c00130031100c1000000000100000000401000003030c40030c0001700003c0004001000004010f0400000c000000000000310000340010105c104c10100003001000010000100f003003000433300304030100130000000000000003000c0007f0c0100001101100100033033004c10103000c3c013400000000300400300004373000130030000000003401041d100030100000003000000100300c3c3033010000101300000000370f30000033003001014730c3000330001300003130100f3300100000001c001311030c30010001110033010000000f0f0000000000030c3000000fc10004000100011400000000000300300010004000140000001c30003100000010010001030130034000000300033f0c0034300000000c0000310001110001003000300100000c4000001410000000d00313000000000c3d1300000cc00c13700110330103330f0c0000004000000c100010040ccc0300004300000007040c0000000c330101030c010303000010000103301030070000500c031c10000000034000000c0000074000004003300000000330300130c03f003c0000c003100c40000003000000010c000014000c0101300c0001130010004011003413000c033030030000c01000c0013030100030030400110001000c001400c1000c0003000100010000301d10010010003c10300400003d000013000cf000d031dc00000010000000100400301f000110f100010010300030001400000000000f3100300000000005003000003c4000100d00c03431000303000010003031100050011304033004300010000003003010030105f001011000000030101c01f000003031000d000300001300010140003403000c0100000300003400030c000c300c1003003c0404010100030003310300030130000d0000030c100133100043000f00305100040000100c13011030040700300000040010303330000010000d00000d0000300400130c0000003001000300141130000001050030104000000005f00100140000400c1000033c100c0f005d1010c00000000410030f1000000004f13031003013330004010000111f130000300004101f0430304300000110000100711f0000300c111c000c300001010c030004140004031000001c0040010000001c001000003c00c0000d170010000030000d1004040000030000000010010;
rom_uints[221] = 8192'h3000000000000030000000c704300d3003003000300c00000000000000000000051c00010c0000000c00400c000130000c100000310000000000007000000000010130000000c0000001000000000001030000001000c00c03000f0000040001340300004400000c004004300010000000000000300000c00000100311000000c0000000040004000400000000300c000000000000040000000000000000004000700000000000300000000030000000c000000030c070100300000003c0000004000000040000004000003000440000000000000c000100c00000003c00000c0000000c4c000030c0040d00400000001000010000004000000000000000100000000c300c0000000000000000000000c000000000400050000000340000000001030010c0000000000000c0c040000001000000000000400001c030000001100300000000300000c000cf000044000300000040030004c4fc00400000000000d000c41001001000030000000c0003000000000c00000000300040000000001000001c0c300000300400004000c01400000100000010001300001000000000110100000000000300000c00000c0300004400000400000000000000000100001007040c00d0000300000000c1000000040c0d0000000000c0cd000000000004000440400c0000c00c00cc000000000030000000000c0000000000000c0000000000000c014f00000000004c00000010c0130001100000400000004300304003000c0000003000000000000001000000000000000030000000000000c000030000001300000000000000000000000000000000000000000000000000000010040000040110000000000001101000000c00000000000000000400100000000000000000004000000000c003000c00401000401ccc070cc000000c1c00000000010000000000100400000004c000000030c00400030000000c003000000000000000000000000001c0000000000000000000c03000000100003f00100cc3000300000000000100000000000c0400c000040c0001100000100000000000001000000000000000000000c000000000000000001000000000000000000300400000003f70000000001000004000000000000003000000003400000340000000300040100c00130c004000000100000c0000000040000c00001000001000000000000d000000311040000cd00000000f000000000c00300000005034000000000c0000030000004000000000000000000001410000000300000c000004000003100000140030000000400c3000000c000000000074004004000000000000000000000004110c004000013c0300f00040040004000000000000000c000000000443300000000100000000000000100004010c031000030300c41000733c0c0013000000;
rom_uints[222] = 8192'hc7c3000044000301000c53c300000c040dcc04011044100300433300c41fc01440003337401c0000104501c0c00301c1500f03c31d1000dd337410000404000304103c03440300d310000115100001dc0145c0010010c003004730140013400c00030034040003c110000040303034d4c00000050030040300000c0407001030f110c00104030333ccc3303000000c03000000050000004034000030c000400c00c10130403043400c05030000c04013001041140000000000000000100c77303000000030007010744001000400d0c0c3c001034044041031c000000301000000104000d0f10100004030c01111c00003000fd3030000c0004004c0730300c0100740000100c00140c00001303005004071c140030100004003000300417733000030000d31000430c0033300cc0004040000431001440040010340110703003041030c007d000041430170d0030400400cc00000d000001010000005314500f1034c0031c0400070100007301c0300d0040104340041c00c0031400000c00cc0001300c330040000000000000c043c04004c100000f300dc4700003404004cf1141c0300000433300000100c534701413003440df40003000003000004c01140c0c0300c400001df30000040000000770014007000ddf0007340c0053404040000110104dc000c001070d30301d030c100c0000101c000c0014500030300470304300000013001300044c70003010040300cc001001000c30100040034c000000700c0c0c00400000f100c34010054000dc001c010ff000c0330004000c3111341010f01001000340000300000007000110403c00411030040000d0c00c13713300c00cfc000000000033133001c00d0c04c044000c00303030c30700304c004340410c0000003401035041417c3c03430cc0c343004c030010000c004c30144d4040c0000000004cdcc43c3450031c1400fd0011f007030000c0500000004c114100030000000003000c0000c000000d107cd03d03c000041c3d0030110010c001310dc3034c000cc00c00000400000111037c01c004000111000000074003700110300c043403300417300cc0300c050004100000140000cc05000cc440040f00000d0000070000100cc004034010100000003770000300145170004f700040c070c10cc01303500340014000013004400d000c10010c030030410000c1400000c700000000100c001000300c3d000d0f300073c00d05030003037173741300041000000000000003000100c0030000d104400300c413303303040cc0030c0007430f000000413cc07030c04301000f00304c30003004000300010d0d100c0df1034f0000004c0140000c0c000010040000c0001c000000f04000c40000001000130010400130007d000040410010303034040010c010144000030030005;
rom_uints[223] = 8192'h1003000000104040000000000003000301c00000c007000000400d010400400000c10c0300050000004000c000c10000043c11c0c300003000d4c3050300000000000cc1000300000000c30501001f004c043330c710000301050100000300000ccc05400dc0cc4c00000300c00030c401c1c000c0030100c00044000000040004000303000000c000000400000003030000c0c0000140000c0000030f0440000c034040000003400100000c01c300400004440000c00307040c0400c101000003cf0040000040050cc040000403c300c00c070100c0400f000c030004c40c0003000000040044300dc300c34000c3000010000c0000000000000000000000c3c0000030110300000000010d11030000c04c404000040000000100c00300c70c01cc0c000cc00007c00000cc0030004047004c00c007c0000100040cc000c000000403000000400004c000c0400000000001010000c13000c00c3d040000100001c00f03010100000001000000d13f07040000040001040cc3000100030000c10f03c303000f0000040000000040144300030300004000000104c0000401030010070301004003000000000400000007000cc100430003004300000000c3c0040015010f00000cc0413000000100040403000000400f404000004000000005c340030054010330d030c10c010003c003000c0000430541000400030100c004430040030c000400c0000f04004fc00000c30101010001004000010300c305040300f0000100c3000300000303c0000000045c14000003c3c400c4c00001000300030001404300004000130003c0c10000004340000300c1004f00000c01040707010d40000c040003404301c0c0030000000001000103000343c4000003004400400043030000000004c00000034000c1c140c00700cd1001000100c00400cf0044c50500000033030c00c400400040100130c40100cc0000000000400f40000c00440000000004000000000dc003014c000004c3c040004c0040c3c304070400c0000403c4c003010004000c01c30000c0000033000100000003000000030000430103430c0003004000c000000001034c030000c143040041000c00cf01030043c0000cc0c10c000000010000c3c0000000310f03000000004000c344430c0000000000010000404143c0c0430fc000c00401030304010000c0c000400f4c0343400300c00100010c000000c0040403000c300043c00041030340000003000cc0404000010001004c0100030003c0010003000305010000d1c00040000000000103000101010003110000030c010000031043c300004003c0c00f00040107000003440d0043000000030000010f0040c10c0040400c004043000303000104c700c000004143c4010000c0000c01000003c00004c0000c5001400cc40000c000;
rom_uints[224] = 8192'h40000000000000c10000000010400000410040c1c000000000400300c000c0000000004300300000c0c00000c300000003034100f1404000100000004100004040c000004000000000000100d0000100c10000c033000000007040400001000300d3f00000000001000030000000000000000301000c0400011001000300c000c3004100000000000000000000000104c0000000004000c000010000c0401003c000c0003000100000004000c10000000003000000c000000000004043c0000000400000004001000040000100000001c0000300000400c0400300c001c00000411000010000000000000031007001000001c3c000000000000000c001000000000000c0010043c0430000000000000003400000000000003003000041300000003400000000404003c000c000003300000000c303000000000300004c430040c0010100c00000004000c10000000333410040000000000000000300030040d00000400051400003430000334001c00000000000100000c000030000d00300000000040003404000030300c04000040040000000000050400000003000001300014c0000400103000040c0000000000000000003c100000000c0c000004000000040000000000001000700403000000300000000100000000000004005c300430000000041f0c00003000100400100000000000000400300c000400000c000000300c000000100c0000303c00000030001030003c00000c040000300c040000000c04003000f00c0004001c0000100000000410000000000000003304000500000c0100000c000000301000004004000c001004040000000004100000030000c00030000c30000000000000000400000c000c00000c00300000000000000010000004140c0c00030400043c0004041030400c0c00103010300000100474001000c300000000000c000000000c0400040050000300040000000003043400000000000c000030003c0c000000000000100000040000000c34003c3c0c0c0000300c0000000000000030000000000100000030040330000000000c04000cf00000050010000400300004400000000c04000f0130000000000000043c0000000000300010000000000c0c00000c0c00000c0000041000003000003c000001300c3001040c003000000000003030000000000400400c100014000c000c0000001000000c000000000000000c00000c0031000000000030000c0000000000000034000000003000000c330400300c000034300c00001000000000040010000000000c100000100010000c040000000c00000000000010000000000000100000000000000c001000013030000000000c0010000400010c0000000030000000000000700100300000040000300000040000001000000000300000000c040001000000000;
rom_uints[225] = 8192'h10000010000000001c000000400000c030000000000cc40c004400000c0000100000000c3030000c4c300c0000101000303000404004040000140c30003004003000100000000c0000001c0000100c0c0030000cf000000c30040c3c000c3000304000d0c00c0000c03000000c00000000000c00000000000000001014c0f000001004000000001c000000000400000030300010000000001c0000303c0430000cd00000001c0000300c1400140004100000300000000010000100000c003000d010000000000000000000103c100c1c0030040c1010000c10d0103c040000100c0000001c3cf4300000003c00f4000010000040000000000c3000300000001000100400300014000cc0000005003000000c0040003000000010000c000c000454001000000c000000001c004000100000300000000000000000c00000000000101c10000030d0000004001c00004400c00c00000014000410301000000000f4004400040c000030c00030c00001000c0400003030000400003c003000303c000c00103c101000000000000000c040000000000010001030004000001c0000000510000400000c000000f000000044000c00000000001000000c00f05010040000c00000f0001030000004000f00000050400000003c100c00000030103000400000c000041c00033400000000c000000c0000003000000400000000f0d0040010000000c00cc0004000400c00100c1004f030000c000000000c041000001400140007c0000000300c141c0000300c00303c04001000100000d40000303000001c10003c0000300000000000500000c0003000000c000c000c10000c0000304010040000100030c030000c301004000c14340c00040cd00000100c00000c0000000c10003010000c00003000d040040040000010703031000cf0f000040400000000003c000c0c001000040000400040040004c000000010303034003000000010400c00000000000c3000000000000c0040001000400000fc300c304010000404000c003000000000cc0cd01c100414000000000000000000000c000010300000400c101030004004000000000000043c400c0000000000001000043c040000700000000000c0001004000400001cc01000001c0c30000000c0001000143c0000000c0000000c0c0010300c000004003030000c300400100c3000000c100c0000c0100010000000c40c0c0000040400300014040000000010003000003014000000000010000c10003000000000cc54001004c00400c000140c0000c400103c301000300c10103000001000f00c0400000c0c00000000000000100000300c3c000004fc10300000001014303000000001000400001c0000000000001030303c3000000000400000d400043c0054f0000c300000c010400c3c00000000000000;
rom_uints[226] = 8192'h44000000300030000400001000074000000000000c000000010100c000c001000000300c0000c004c10000040000040003c003000000000c0000400c004000000050000c000005000040000000000000003c004000c40c000104040000c000044070504040000003c44c00340041070000040c00c000c00001010000000000404001c0040c000f0400004c4000c00c0c00000000cd0000c04c00c004100c0d040c0000000004000040000000c500000104400000040c100300001114000c014000004c0000000040c00c00400c404c03000c300c0c40040c030040c000000001000cc0000000000300037d0cc11c000c000405fc0c0c00300000c000000000f534c00c040001300000004c100300c4000301c00043410004110004c100001040000000c0f00051000040000000000030040000000040000040c04001000001030033300400f300cc11430100000c00d0c04c004311c1404c00c0f03cc000c0004100000000c0405040c0304c4403030050000103000010c44070000440000043400cf301000c0034000001440101cc170004003c000740c404000040300040104c0f1000c1400d00040000034310000010004cc4c00d000c010400c0f01100c40010c0f0c0c00c00314000000400000001001000000c0404000c004c403000c00004c00000004c00100000003001c003000100c044c40000000304100000c04003c0c0000d4c0000400330c0000c410030c0104440cc0003330dc730000f001c4400400004000700c000c0c100000100c50000000400c000334d10d00030c0040c00c003000000000c0000c40040f000003c003050c00000300000001003040010000c0c500005040000400000000000000f00f0040000c4300004400000c1404003c00100000c0c000007000001443d0c0000000000400000000111000000004c40cc0400c000ff4741047f030d10100c000000000000c00004c0d10c0000c0c0cc40430000300000000c000300000000f000404c00c0c0034001c10f0c00000000c000040000c0c00000000010100c0030400c00004000c03100c0400d0000300c0040c004c10400000000303000c11c040001000000300000003000044000000000c14c004004000004030000cc00004030400037004000000003400700f3c4f44c440700000000005000400c0000300000001300010003030000000000010003c000300001c1000000030000000000c00c4004c04004c4000003000cc004000c10000000400fc000cc00303c00400010005c00000c00c003c05c00000000400031f00001440c0000400043000c00cc0000cc000c0000000100000033000000010fc0004130430c000000c00000414003c00000000000c400000cccc40c50340cc0c000300000000004c0003000300004000000000cf00d100040003400;
rom_uints[227] = 8192'h1c0304c004040300000c000744000070330000c0000400000000410c010c011c040c0c77007000000000000130400c0c04010043c0c400300c000004000700030000040c001f00030300c00d01000f00000000000c3d0000f10c0001010f0300040c0c07350000400c01f30001000044004101000000010c0001444000003000317000000447040c0d1000000c000000000000000000404041040001030400004000100000530440000000030d4030400100c0400030030341000010400100000f1f00c00000000c341000c30300030d0100c00f0000000003010f0f10000400033300010000440000000001100101030f01400d00000000040000000700000c44c0040c0d30100c041300000f00000000400c0407000f4001410c0f0405031430c500000075000700c0000f010cc4000003300704000c0040cc000000000010cc00004300030400000404040c000c00050000400400401004000c0d030010000503004d00000001004f000cc0c1fc03000000040040000c03100100300040000300170000c00400000000c3403f41c0300ff30000001d40000005000301004000000f000007000000400100000f00000400400400410310000301400000014d0c015100010100f544044000030000010f3f00000300003300030c044040c0000010c304000010d4744014410001000004000c030000310000050000000c00340f03c401000c3000000000010000440c103c00000c00003c0540c3030301050c000000cc33d0000000004300000c000000dc0c0500030100c34d3400010000000714000f04000000cc000037101100010007c040030c00c30c414cc01c0007030f0c0c10fd00000433000c13300001003d000000300001cc0f000000030c300400100c04c10000400304310f17031000c1544c0103310001003000010d000d00c70501000300470f104f0c030c303c0c04130f0d000005040030003507003001040304000100000004030000000000040000c00000003c0004007000000f010100004f00400000000070000d0400000c010d030001000004040004004f0c01003011040000c00c100000000000004400c00c40004000300300000000000000c3134f0000010cc00040dc01000cc000000103103103070c00c00700030c000d000400000c0000000c0000000c00000c04030000000000011000040c00004000030c0314000c3c01000010000000000004c4100ccc00040f0c130d000c000000c0c00c030040000000070504c540003401cc4c0c04000100000c000d0c0c00000d03000440c0010f001403000c05000c03000303401c004004c0003000030c000400c00f4f040405040100c30c0101000c0000c30004000001003330000331000003000000070301000010000010004104010f00010000440103040c010d000c00;
rom_uints[228] = 8192'h1100d00000040000c004c000fc00c1c0c10d414041307c40004103004401004100c30007004c00004c0c00000cd04010701040013040000100c10001330000040410c330000030000c0000c0cc000400300100c140010f004f1007c40030144c0030014004c44043014cc0f0030f000040c70000433000000003c001110400000c03040000030004001101400d030041014c0000000410c30400c000c04000c03001000000c700100000004030000c0c03000c40000c003c010010700001000000000000c400033030c000000c000c3400c0041040013c000000000031c30404000c00000000d00000000031300c50104400c03440000000000000c000000000c470000040000000030443c0f3070c3003000034400d000043100010400140410000000003000040c000c0c044000700500d000000000400c30000004000c003000070c00030000000c300f300000010c0f0100040c0c03114413c000000c4c04011000dc7004000c3c100c4044000431c04000043040000c0c0000000000c0c40000000100044000401010034c000c70000004000000cc001004c00c00cccc0cc7c010030f0401000031050000f310000030400cc0000400c00100d300051f1c0c10100c050401d00f01000c100c00001d0000040030c030007c0c000000c00000c01c03000110000c0044d000c40305c000051fcc04040000000034140c0000000704010c00f00c040071000c0c0d000d0cc40000000c040c34000c040433000415cc3c344c0100000070c0030c00000c470030000c0400030d000000000400100c000c30000000001400341040000000101040030cc01c0c410cc03300d0501000000400c00000003c3d000404104100dc0c30004400000000000010000100000404300000030000000c0d010310070c7cc0100004110000300000134000000004d00c00000000000c04c0340c0f040c10010004040074d00010730000000000c00c0c0000000cf0000300c000c03000c00c00070cc07c00010030040000c1000000070400040000cc44000c33000000030c0f0c00000010033cc00c00400404300003710c0c401c000040000003c000003c00003cd40000700c1c3401000c003d000415000d000c04000010040c000000000000c00300100c0000d00000c040000001c00010000c4c0005004c140000cc0004140300010300c0000d5030004ccf03300c100c0000000c1cd0c1000400000c5000040c030000000010d00300040c0401000cf00400c000000000000cfc0401c00c0c00001f44cc4c0000001c1000000c000c0c00300000400c00000000004c00400c04000000300000011000000cc040c40f01000000000cc0040c1000000c370c30043000041c40003c1c0010c0040431ccc00000140c3403100c003c04000000000010000003051030000;
rom_uints[229] = 8192'h300330100c0000301041004054001c013c000040c01c001000050f000400303000043f300110000c004c000000000c3030000c0fc0310040003000345013000001001001000000300000304c10000000003000100001100010003c00001c05001050440000031000c0cf3000004010c00000000004003000001c103001340000c00030100013005000c000cc00500040000000000000000040d00000c310003000300000034003000000000000100030014010000000d000000003030300f000000100000000040003303005f000301000000f0c300000403014000c003000000f100010100c40000030107001f130003000031c5c110000000000100000000c000004300c307c00001000000f0000f030310c34000000007c3000000003c35000340400000030f0c000100c030030c00010c0c700000000003031503030103043001040104010403000504300003cc0f0040043003000c034000000000c310000300000000000003000000010d000000000000cd030000000c00100001010000070011000100000000030001c00f004100000100000f0104000000430c00440c1f0f1c0000000001000100010033000303000c31030043000001010301001004c01010010000000104000000010700000010100d10304130040300c1cf000001001010040c41000405c7400040001040000003d030d10004010000000000000c00004cc073000000000300004d0c0130000003010013000143000001011c5003000001cc0300000000510403000003000c0c100000053c0000003000000d00100343c3000c0c01033c010c000d0110000c0003000400000004d0000100c000c3040000053700030001000004000040030d010000010f0c003004050030000300000000010000041c004c003c0f0000044007c4c0003c4000000d00c5c31d00000100000010010300103330100300001c0c011004000004700003500c010000301000f1c00000000001000000000000000140030540170003033100403c0c00c0000004000c040000010404000500000003101030430030004000000cc4000001000c010300000501000300000400c44000000003107303000341030100c1000c00c005c310130000c0c0040000010000d0000000010000000040c0071300300300050700c14000c3030000030f0000000f05c00c0c10003f0441c103031c3010c3003c1300c000c300000000400c000040003300003000000f00000300cdc001c30040000000000000040303011404c0334c300047c7000c00333000000000030001030001c03100400000000001c000040140c00005000000013000000f010300c00c000d400d000300c00003100000f0000700000100000000000030000000000000004f000000c00300000000070037010010100403010c003c300100000;
rom_uints[230] = 8192'h434500f10001000010300010000000100040410041f0400003c330300001015400300003030000400000000f310003c03d4003110000000f104001c70300444014c0c3f0000c10705000030000f000c4510330c01c00430003c50073001034c01001c0004044700050001003031304c00000c03001000330403030007001100000000140000000000000c0c1f04000000300410000054010000010000070300030000000300000344070040000f000400300030001100313033000543001003c0011004104000500100400101010c4000c107004f011001030701000d00000004000400007c0101303c00000c00fc010011000000004000000000000111000f00007f1c000f04140101040010cc030c050031003030000c3c340000013110000001000000000110110f44000004030000000d0000000303d04c00040f034100030013001f0001d01f0001003340000000171013003d11141405031431010040011500004004140310f1103034c00030013c00c00001050010003010010c0504f417040000300000010c001301000c00000000050000003c0400000014000310000f00430000c0740000c0000300000104110103430000000110307000403400140000c000000000300000330000040000030f010c000f3440c04430100103c13103031400030030150000000000000f01040c0004340005030300d03f001100100014310100033400111400100000040f0003003110300000354511033430000004040000033c00c1001003c0030c30000030c0000054000400001000d0100c31003f001001103000011104003c04047000441000000c0710030300010f03110434103000300004000003033f07001004c133003040000003100014003c1c000000cc0000150003100301040101350f000501040007100000700130030404000104040c143100001400000004103000040c040d00000c30000000040404c40114003000350000400514000000001000100c0003033330130d003300000000000d00003000030000000c100c040004044403000c05003101030000003404040030530c10000044d000030003070d00040110000303003c1f0003c0300c3000000c0033103054000c000000004000554100410410000000030f001030010c000c343030100400100030015004010300000c04010000000c0004000c04030000100d000001110030000c0400000000000000000c440c3c003004300000000f0c00310004003c000403303000100c130c050705c40001013000c00030010400304100000105001c45c11403001c0010000d0c0005000000000000000700000cdc14040000000000cc000530000001001000000000000c0300000d13001004141004030c00000000000400000330340031000000000f1304050700000000;
rom_uints[231] = 8192'h300400000c00000004000010001000300c04030014000000001c0400330c04000100013c0000000400400000000000c00c0300000030010400104010f03000001000341000000034000000000000100500000010030000000011000000000000033c10300000110000003300000000003050000f00c0001300103000000c03000405003000040004000410001000100c003c003000c004000c000000043000310000310000047030c01010000f000004103000100000301000000000c00010000007001000001000300000100c13050c001000300000000010010000003c00000130000034303000000000d0000c10000c003410004400100000030040000010040000300c0034000000000014030000001100003003c0000d1400140000000c00d1300004000010000130040c0000003044d0003000000400000c00000c00000c00003000300000010100300000030011003000004400004000c0100c4c1c0000000000000134000300303030000c00000000040000130040c10c0c000010100400000040040000d030000010001d3c000000000000300003c03000000000001c0c340004000035003000300000100000000000700000000000000000001100000c0030003000c104003000130000000000000010010030003c0030000000300000003c0c1030400c000100333000101500000300003000100400000010000c0000000050100c0000000c00000100300010000c3c10000c0f000003000c000000000000000430000030000010000010003000040030041030103400000030000c000c003c0030000c00001c1000000000003000000014000040000c4000000007100c300030000000013070000300043300070100000000300f0030000000000c001300300000000c100f000300cc30000330031000000c000000001010f0000c000000000c34001f0431400310001c000c003000000000000000000000000001010000030030003000000000030000000110300c1000001030000000000000040004000f00003000c30000033404300c0c0000000c0000000000000011cc00000c00000c3000011000000000000000000c0000000100100040001000300004111000031000040000000010000000300000300000000c00300c0000001c00000c0030003000f000000c303001001000011c0000100000c00c0c000000100000000d34300c0000000000000000000034003034103000140010000000003c0400100041000000000000c000c03000000c0100144c3033300000040400343000001c0000000c0000100000000cc00000040003000030001c3000000000100003000c50010c300d003400003000300000000d00000c0000000000000c004000000000000000004400300000000000c03000c40000000300000004c100000c000034;
rom_uints[232] = 8192'h10c000000400000c410c00033000000c000c034004c3c00c05c10000c0c100c0000d003030c400c00300000c0ccc0f04f104cc40c100c33c0443000300040d05c30330c00c0c0003000340400c30040c0004000fcc00c0300103707007000000c3300cc04040000300c0340400014c0003403000c1000100074000c70dcccc00cd0c0f00000000400c0001c010000c04c0c0000000cc4005c1400000c3c000040303000c00400f0c041001c1541000000dc00000030000030000000070c040cc404001100c0004000400000000000c4f3c040f4044010c00000054c000c00000c0000000030c40000300001404c00cc0140f7c30000000000000005000400100c0000c05cc40400303000030400fc0001343c010004400c040304f004fd4c000000cc00001c004000c100d000000000c0005001c0000000040040c14000300c3c0c4034c0001c00000c04cfc00410014c0d041050041cd433004d40400000c4001c0c0340000cf04c000c0011000c33c1000000000404c0300440403c007400c0f7cc00000c1014100d000044004c0cc0c400300000004014043c04c0000000417f3400101c00c00003c000043400004100000070400040c0100004404dc44000403000000000f010c40700040004003400300000c04104001c00000404003c000c40444404c01000c033000000400d701000000040c0d305d01000c000040004141030040045000400510033010cc000104c40c0040cc01c000cc1040c040c0100003404000c0c0030c003000000405071400030c0004d0c70c00000003040f00000c0000cc00000001c000c70000c01f00400000040c00040c04014054c003030400400300000040013000c0040043700c00000c030100c00c01c01c0cc4000000000040c00c0105c000ccc000c34741030f10c0c010c000110001510003040004c3c000110c400040043c03404400c0cc00c34004c00000c001c0034c000000001c0110000c000400004400030300cc000cc00000010010c0ccc000430010000cc00c01fc30000c1000c00c300040c00400c0c0030000c004c04004410000040000103c0c0dc000040100c000000d0040004100040500000c010433000700530000c0c4000c100040004051c0c0000000000000300003404000fc050c10000cc3410003030dc0cc403000400001c004c0434304c000c0040c00000c4c03000400730003000000c000400400003c0c0000500000400370000000400f0004c00c000000440000400300c010000000404000c0c4cc0c000f4373400000f00040700cc000311000000000000000000d3000dc000000c04004010040010f4040c00c004030030000010f00d000304403404c0000c4000000c0c000cc1c4003000000c0400440c7c0c00f0000c0400030134d0300000000011311c304c00000000;
rom_uints[233] = 8192'hc0100000000003c03033000000140100c00000000310000140110313300000000134d0005000000010051c0000001c0c04407c3010100004100000001010000003d00000300d3c0000410400303070000033c0103010001044010000007030100c00101000010010131000100001000140d00307000330000130000003f30103c100000010030000000000000300300500010000300343c03000c00313310043d010c03030400030000001c130003d33731030030003340110034000030010fc4003000000300110000100170051710c00500100000c3400d03000001000001000003004d0c000000000000310400030000c733000000000c30003300000313000000440f00cc000300040003001000000133404c010000000030c30000c100400d000400c0000400c100000330000c0000300000040000700030150104030c4000010000c00000030d003300c0110000c00001110300c300dd4000000300400c3c015010310c0103040101000001000d5d33300400000303110c000070004cf0c03100034000003c010050030400000000000000110000c10510030000001501000330030030000001000010010c000000030010073033030c0010303101030d10003f0001011c000000f3000300330401000003f03100000301300001000000001341d303300033100707010000010300140000010000000003c00041300f00004401130100070030010033000f000000500c300000300100000041c400c1000100101100030004cc00400000c30dc0740000c000003c410c03000013010000503c001000300000c7c00001400c0c0334000001040003040f0c0000000300010300037000073c30000100c0030010007043000100000001000000f0010400000004000d000003301001cc03c101004440000000000000003000030000010000110000000c0300301000c000400c51cc0003010001c0043000f0034c0000000304030000000300010110010000400107c114300340000c40000c000340010100300007c00303033003103103000000d4050c0013410301000000130303000c01000c00300000110000000000013403334c001730101001000000010000010303003cc0010000000100410003010000c10c00004101000d00000110000100003c0010013400010dc001000c00d500000100000c1100001730000000c33f00030000000010003000c30010310100033c0300030100443404000003003d0300010344010100330030000100010040000300150001000c00114000030cc1000010010100c000000003300000c000003003000000c300030000c00c00000000300013000001000331010004000004001340003110004c011300000030300000004010000000030100010007301400304033000100010003000000311101000000;
rom_uints[234] = 8192'h10110404430000000000030c000000000010000003c0000003000c00003c0d00340000000400000400030330d0000030000003000c10300440000000000401000030c03000000000003000400000004c00030004c000333000303000040400000000000c00004c0000f430000000c0030300004011c0000300400000d000300000000400003000000401040000003000040000304000000c00011330000f0400003000040000000000000000000010000000001000000c0000cc000030300010000010000010000c004140000000500000100000433003004300000c4030000c3000100c01000c1003001000000400343000000000003000000000000030003300000000003033005130000c10c400000010000000100044101c10000010000300300010000000000000000000cc01100004000000000000c0000000000040040010300000000330000c0000100cc00400000010030043103000000000c0000030c0000001001000fc0000310000000030000000010f001000000c00c0ccc004040300000c0000000001440000000000000c40040d0cf4000d00000c0f31010000000000000000000400141000000051401000000000c000004010500c00033040000c0000100c00000000010c00000c00410400000040010dc000000004001000000001000001040000001c00000c110000003000000000d001110c001c054000501001003010003070c040401100100100000c000030000000040c0000000103007330040003000043000000001030003030000c30000000004d0c00101000300000001010003001d000000c000000000030004000000000540c0033000007c000000000303030300000340000c0001000c0000000000000000000000c1000000000000000033c000000000100c000030100d0000030000c00000c1030003c10003030040000040000001c0c00000010000400000fd0000000000001000030100004030000000c0300000000c0000031030000101000041040000300000000000c37000400000000040010000040000c03c0000100c000003000003000100f0030003000000000040000004003f0010400001000000000300030101100000c0004000003140400000003300100000000c0000010000000001300001000070000000c00000c0400103040003c40300c00000400c007000000cc0c04000000cc00000013300400030000c000004401100000000000000000100100000004000000000000c000c0100434300000000cc00400000c00000000400000003c00100440010001000c00401000300000300000400d04000000000000001400047030000000010000400000003000500000100010300410000c0000300010013300000000000003000000000c303000103400c000100014331000c00000300;
rom_uints[235] = 8192'h3000000000c0070000000104000c0c0011d0300003030100050010004000c003001143404000000c3c0000000101000041130100004333410400301300003100110040000100000d00003c0d430000000310014c013003030130004000c3070000440004c30d00303343000034401341000000f0c0010410034400c03053300700300000000000000000c0000000c01003300400000000000000041040100070000300c0010000300010000030c30cc00403010000c0030000400000100010c000c00300010100330000300000101100000330300000430c0cc0001303410700c0000033000040000300400313c0000000000100f00000000003c031f000000000300030400c000040000170131000c011c001d034030000c1300000f3031c41370110000313000000c0f0000000100000030c00000010000304c0c000c10c00000c00030740c00100000001c001c030cc130114113151d10001034300010100000400033d031300100000001130104000c30400444000300300000c00300030c0c1000044700000100403043404c040000040100000c000c003014000001400c0f001000430000003c0000000c10003470dc400000c0403301001300011071cf0000c41100001d00c000000d000070c0030c1000000c4c0000c03c0010334030c0013c3cd404050d1c001f000000f1c0004c3000030300000300c0400030c35c3000000410000c004401303040041000040000000003004c003c0c000c00000041010000c00000003407300110041100300c000cc100000030001007000007000450003000010030000003001110400004104000000000041c00310000000c00000003330c0007000000040010000410000300004000c00000000030c000000400000000c00c0010000004331011000430703000040300000300001c0100010110000300c0000000101c4101000300070500030041000000000d44cc130003300304100000cc000c0c001000c00f003003c130100c40003330330300000404c000000010003c00000000003000000331700c00300700000030cc0cc0001c00700004003d04001010000001040c0c0001000033400000103007330000000031144c0000000c3c01000500000000103400000430004000010070011004313000310dc300700c0003000004000010c43d00300003007030701401100031110000003000c00000000cc1000c00150000004c000c0103003003003000000f304130f0105100000000000300c40000000400003004100c100001103000041040001404cc3014c110cc011000000c0400100000dd00100000100101000000131c0cc000050c45cc43000c34000100c003000000000000310f0000040001000c40c0014000100000c000001100030000041c0033000c000c000005dc03000000000000;
rom_uints[236] = 8192'hc0000010d000033000100400030c000001000003000000154000000c3300004c0444c30000033c000300530c014c000cc0000c1001340404000c0004ccc0000070000000304300000f0000401d34000c1000704c70003c7430dd0000c00001700401304c0c00c704300c3100040f4040400c070d0010001040c007d07407410000000400044c30001300c100c0c004c007000c00000c1001d3000004c041f3d4300000000333000003033d0301c04c00f140000010000000000000341015c00000c30c14030400d00001f011f04400103000c00401c0000ccc0c0400040000c0000433400005033000100d7313000000714000c000005300403f1000031c003c1c3f33413004c3401c40004307101dd0731010003713004703011c000410330010003d000310014000000c000c03334703000c00000030701c7f00010c114051c404040000001000004c4000000c103000011dcc141c40c400031d0cd000430c0100c003c40015140430c000100030100003004030341443030c0040411000c1d0004100110f10040010dc0010104003000c4004f0c0370030c400000003d00030c4000000000341000001340cc0c00001c1370c1704c00770300fdd40003c01700110300140000004c400000044c0c000000c0334700003c00000c4f4000000030403010d10cc00003ccc40000dc00413c5c0003c00c000c001100c03033000dc000c04d0004413040030001030d7001001404c0077001c310c000d010300440073030000c0000c300110101c170c7cc0000001435304701fc4000c7c3040010000000c00000000030c0cc10400050001d0040c00001c04400c07c00705c00304010000004000040400004c0004001000100000003303013c74c4000c00313c000c700045001010000f0300103c00c03c3c140003031000000c13140043d05000300f33003001704314040100d10010307000000c434000010004c030000000000000000140100c0d00040cd30000301c0011000f0103c0047043003000000401fc0300004f0000017c4c4003f13001c4100004400001cc300f43331103000c10000500030010040cc40c401100143040c0141000003303741000301134c000010c1000400040000110c4400c000000000044100004041101100700c000cc0030303430300014000014030c3c0c1dc0400000100c00400000000003701304d0340c030000040034010401c00d3010130c04004300300f700010c40000c03c0c330c03070003c00100d00f00c001f0000000c0340004300d3001004c35410300050c30f03410430407010004000000c000010000d000101440005c0401001000c0d331040100000c00c041c004000001c40000000140371413007400c0c0100000d300cc050030cd001103000000300c4c404043c0fc0c040c070400400;
rom_uints[237] = 8192'hc0000040004040000000000000cc00000040000000c0000400400c4000040000000c40000000003c00000000444000c4c00cc400004000000000400004c4400040c4c00000000c400c0000400c00000000c000c700300000c00c4000c000000040000000000404c00000040400000000000040000ccc000000003000404003c000400000c0000040c000400000000000000000000000004000004c40000000c000000000000cc0000000000000c0004000c000004000400000000003000000000000c00000000000000000c004c0040000c40000000cc000000000c00000404040000000ccc000000004000000000040c00000000000c0400000000000000004400004000040000000000ccc4000000100c04000c0c000444004000000040400000000c0c0c00000000000000004c000c04c0000000000000000004000000c0000ccc0000040000000cc404004c700000400400400000000c0c40c0000000000000000000c00000c000040040c00000000004000000400000000c0000d0000400000010000000000c00000000441440000000000000000000000000000c0000000000000040000000004000c0000c0000000000000000c004000000000c0c00400c00c40000cc00000c0000000500040000000c00040000c4000000004004000000000000000000c0c0400400000000000000004000040c0000000000c0c4c000000c0004000c04000404c00300c40000030c0400100004400044000040000000000000000c0000000000040000c000c0400000400000004000400000004040000004c000c000000000000c000000000c4400000c4000000404000040000c000c0000400c00040cc4000000000000000c000400000440c440000000040c4c0400440400000000000000c00000000c0000000000000040000000000400000000040c0000000c0040000c00000000400c0cc0000c0000c4000043040000000000000000000000000c000000000004c0000000000100cc00000000c00400000c0000c0040000000440c0000040000000040c0cc40c400000000000000000c500000000000c0004c40000000400000000000000000c00000c00000c0c0000c00c0c0000000000000000404c0000000000000000000c000c000c0c0400104c0400000400000000000440000c0000044000c04c00c00440000000c000000000000000c40004000c000c40000000010000000000000004000c000040000000000000000400040000c40000000000000c0000004c4000400000004c0c000000400000cc0000040c0c0000000000000c00000000000000c000c0000000000000000c0000c4000c00000c00400400000000000000000c000004000c40040000000000c0000400000c000030004c4c000000c000c00000000c000300000000000000c400;
rom_uints[238] = 8192'h300300c000000400030000c4050013000700f10000003000004103003c01000100001f00c434000c0c50000003c000c044c000cc00040c04034cc0400000400000c000c0000c00c0c000004340000301c74000dc314c0000f00d00130000dc000cc100040000c0000003000030c04001010100150000011f004000c001c3030c7703c040c410000c00000100410000c003c0000000000cc3dc40400003c0400000004700001c00000040010003cf0015c00c40c000030003000000d0c0030003000d004400000000040040c400c001000300310000c14000c00140130003000000040000004c0300c30c00107001c0003dc30000010c0000000000000000000000c00000d00041030c00c0c00103101400110450c00d4d0400000f0001300500000c100000c041c10000000c00003c004170000000500100004c01c0c0c104d00040003c030dc000410d17ff0c000000103f001000000c00c0000300000140000003c313104c00400c0030333305044400507410004c000c000d0340c000cc030004c1c0110000004c010000000050300f000fcc0c00000cc401004c01010c03001400000005c04000c00370000cc00d700000f150101c0c01cc0c0100c00040034101173f000010c340444040000340c0d0c00141014331c003410010040101000003540d0010c0050cc000cc4300004d0300000040004340030000c4001400313000c030434001c0000c07cccd004f500c03000340c00031034000030c300044c5047c4000000000000f00dc101000300c000c0300c0d0000003c015000c0000704303030cc00000000000cccc0f037044c1000014400050d000000c41345c01001000041107c0001000503f000c00300303000003000003ccc003030000030000000100030c0000c000333c010000011c5000140331010003c3000d00000040d0703050030300114cc050004c1050c04400000700c000000040c0c001000000010040300000c34340030000001010100cd4c330c0530c4440c000cfc1714103000c00c00000000030003300c0004040c000c300000000c044c50000400f00c1c007710704cc1300000300000003c003510f000000430c00303344cf30004c701000000000c3404343011000c001001003003000c04003404407c40070000000c0c1cc0000010341c0410014000300d3440f040500c4001003c00014100cc40c4044000000014c0c4000040c000cc00000010001000000030044d300003d00001100010c0003000000000040ccc000400007f00000304000d340007c000070035030000030c0030c00c04c074c3000000c44c000000000000300000001030401301c03000103c70040540003010040000340300010c44100c300300050000350004013445d0301330000001c00030cfcc0cd0c0004cc440dc000000400c300;
rom_uints[239] = 8192'hc44000000000140003c0000040003010c000c0c000000400d010000000d0000400040043304040000000003000000033000000c04000007000000000c00000000000d0c0100000400100c0140000c040400000c0c10000000310004000000400c0000074c040001000003000003030001000c030c0000000000c0000000000d0100000000000c0c000000040010000000010000000001000d00000004300c04010000000400000101000000004c000100040400000003000000000000000003010c00410000040403340003000003010003000c000c00000100000c3000300000000000000c07000000000300000000000000cd0000000001000100000c0000000430000005000000004503010c0cc000010003000000000100000d000cc10000000c0000100000000000000004000001030401010003c0040300040301000100000c0004000000010000003141000000000000030303031c000300000d0000000c000c0f3000010000000000000004000c00c000000350000000330101010000030c030c30000000000c0000040005000c000000040c5300010c00040100030f0d00000000010011010c010300c01100000000034c40000c000d00000000100000c00003000000000407000000000c0d0030000d040c03000001000001000c03000000010700041000c1000000000000000000000001000f0004000c0c01054f0000000400000c0004310000330000c000340007000c0130000001000c0c0400100c11040f000c000c00000f000004000004000004000d00000c03403000004c03300004010dc0010000003010110f35001100000003000404400004000741004cc0000000040d0000000f000000040c000004000d0c400000010004030000000c000000000d00410000003000000000030001000000040000030003700000000c000c4104030000070740040334030f40030040000c040dc0001100010000000007000000000100030000000301000000000307000000000400000c00000000100000000000000000040010f0000300000c300004010300000100000000000c000300000040030000070000000000010000000000000c00000000003c1000030dc00c0c0000040000110103000cc030000c03340c00000400040c0401010000000d0000000005000000030010030c0001000c0003000000330000010004004000000003000000030000040f000c00000040011000000300010000000d01010000000c0000043004100c000000000000004c000000000c00000d0104100000000000000c030c000000000103040004000c300001000000000000000000130000000473000000c0000003000f0000040030031000000c0d0000010000000000301c000000001000000c00000000030003000d000000000000000c0c0c0000000;
rom_uints[240] = 8192'h415000000000000000013000000000000000403000c00010c000004c001d000000c010000c0c000000300300040030104100440030f00040000cc00340000300000400c400040000401000011033004c000c10004000d4c0000f0001000000c000400c030000400c01300100010c043003000000000001cc00410003c00c00300000400000300000c3000100c00000000c000000000340c0400000000c00100000f5040000c0c000100010000000003014000c0044cc00100004000040010000d00000000000170054003c1c00000000c0104c000030101000300000000f300300410003d010700000c004cc4400100030000000030000000000c30000000c000400cc0044041000010c0430c000c033c0c04000c0140400000000000000000000343000340110c040030000f301000000000c0100304040400010537000010000040c40dc0004040054004000c04000004030c0000000000000010044000000037000013040c00000041c04c0c300c0031030c00000000100c000c0000440300004c000000000004c0000000c4000410d00c00c0004050000004000040c5000000004f040c0103004000001f01070500004030c000103440100443400c00000f10003050014000000c4c000000300c0cc001c0000c400005000000410001000c000cc4030000c0000400040700000004030000040c0013010cc1003c000c100001100c000000000c0551040300c00050c0c00000405003030403010040040007c0040000001001300000030000504c00000000410000003100400c0ccc000000000040fc004000000c000040004c1003010140100004430000c7004000c30000000010044030044100c0000c000cc300000040c100000c00100440010000c00403400c00c0c1004000c00400010000030040c000100400c000430700c4000c00040c030000000041430033000000040c0c3030400040000c04000c3000000c030000c0000000004000000000f0344000c14c030cc00c030000c000000004000cc00c0000000040000c000013c0000cc00c00033000030040000000004000000c040000c000000000000c0c00001c00004c010cc0400300003ccc110004400000000400400c013c00050000c000040000000100d03000000d001000000000000401404340003c3cd004000000c000c00c040cc0f00001100001001000400000000000000004c00f0000401cf0400304000104400011003730004400000c00000010c300000300000004044000000c0cc00300004100000000c34c000404c0000ff00000000c00cc000000000041400c0001000c00000000c0000c0003000c33000430000000c4000c1000000000041005000010010100100030000c000c01000000330300001040c04cc00300330001005001c03c00000000c;
rom_uints[241] = 8192'hc0400300c340044000000000c500030303000000004d000000c001004300310440c0071f00c000c000000400cc003000000c400150c00110c0c000004c00440000310c004000c0c1c30004c044001131c3400c00ccc000c303f013000000c30c03c04c004440010000000d00c013400c0000f300c0000100001c50c4f0000f0000040400040100c0000000c0c400c10000c3c00300000000403000c000000040c4004000000ccd130340000301000000000003000000c000000000300103000301000043000015400c004001c00c0100003001100005031c00c0c0c3434f000001000000dc0043000300001103400100c104c1cc0030000000400000000000c04001000000cc10400c0000c0000c04000000004300440000010100c001004c01050d00000100400000d10000c0000ccccc001041cc44010000c0400000d001000100c54cc0401cc303440030d1ccc101004004c043010c0000000540400003000070400040c040030c0440cc4004c10c00000000c00104c01c0c0000000000c0c001c000c0c0f300400c0000c0000440c000c004c0001000000000000d00c003030700c0c011c000000003000330051040c0c00000c030000f0cc30000110541c340010000040000434d43000300c000c4000001c3404001300c413c0000c0030c400400c000000cc4f330c40c0100000100004004f000c700000001c700001c04000dc40c4110010003034013c013c1c40c0c0000000000c4000000d33000004000000f100c0cc30003c000300040007371c4000000fc0000000004000000000f7003c04c0001000003c40004100300400000000d070d000004c00000041001c0400000c0010001070000000041010000003010300000c44000010030c00000007011001000000100cc00400010c000c10300000030000400400000070300404303000c00c00140c4400003cc471c03043100004000000000c0404c00c000c051100000000000c34d040400000c0047001000010cc0004c4f3001030c0034030100000000000cc0000c00000c0000040000c00c401000400c000c003003000003000c00010000cd05034000004100030000000c040000000041400004c3000d0400000340014d3c0030c0000c0d003c0000014d010000030043c000001700403041c0c00000401000c0c300d4c1c0c030004041c100000dc04300c0030700d3c0007001000c000c404c03007000071103000100c3c0000000c0003400030000c0c441030000030044000040000001000007c50343014000040000004000010000c1430031000000000c000043c00510000000004c00c0010000c00000000c00001d000300c00013100104000007c001000340004040000cc0130000c00f000007000001500000c00104041000010c000c00c0000c0c00730c000000c3c00000;
rom_uints[242] = 8192'hc00000000001400040004400c000c40000000000000cc000c0000010000400004000c00000c0004000c000000c104304047004000040040000000000000000000000004040000000c0cc0004001100000010c000c04000000c010c700000004440300000040c0cc0000000400c70000000000030d0140000c00030000000c00c400000c000400000000000000005000000c000000000010000000d0000c0000c400000407000000c0d00000000004400070c00c0000103c000c1040000000c00c0000000000000400000c00c700000000300c000004c003c400000400000c0c40000c000c000c03000110000004000040000c0000000000000000000003000c00000c00000000040c04341000001c010040000000000c0d00054011c0044040000004000000100000000c000400c0403000000c005000000400000000400030000000000cc00004000000c00c004001c00003000004400004000004000001c043004c0c0000000c0000000030c00000000c00000000000c0c00030040000011000000050000c0010c0004000004c0400ccc00000000000c700400c13cc403044c0000000001000000000000c044000000031040000040410004000000400305c00000c0000000c0c00004100040000000004044c404000400000c000c00000040004000c0041c7030000000001000c000000400003000c000000044040000000c004000000000000000030c0cc0001110030000040000100c50040000c00014000330003c0000040004030c0100000c0000004c4004000001300000000004040c00000001400c0010000044100000000000c00300000000000000040000000c40000400003d000c00c1100004000c003300000004000000000000000c000004040004c0000000000000c1c1cc000d0000010000000c00000300040003000410000000003cc40000c00000c04000cc00c00030000c0400400400c0000000040000000000000000000c000c000c000000000000300000c4c000300104000000000c00055c0000400c310000c004004000000fc000c040000000000f03000000400100000d0000000000000001300000c0404c000000000000000000300000000000000c10000000010c404000040000000c04c0001c000300c00c00400f0c004000c04000000000000010000c04400c0004004000c0040030000000000c00001000000000040404c000000000000000400c04404c030007000000000000000c00000010000c0000000000000000cc0001c140100000000000000000140000030000050000034c3000000000000000000004000c1000004c00000000000034000003400000000c0000000c4004000000405c0000000041c000000c300400000c400000001400000000400c0300440001c00000000030100000000c30440c000;
rom_uints[243] = 8192'h40300c003014000c00d300010c000c00340414310030040300040c000000003400d3400330c0000cc0040c30c0004c0003104030000000c0044330c430000014c00c1c0c1003003040004f0730000030000011c3c7c700010cc70c0d300000cc0c7fc30000003300041c0c000c40300303000c301000c40040300103f0001300c00140c0340400140000c00c34040070000c0010000c04300000c10030cc04000100300000c00c000c00040c00000100c000010300100c401040070000ccc1cc0340c1c10004044000100007000c0c0000000044000400c1043300141000031000010040033000000c0c0000000404000340c003004000c00000d00000400001304004040001050c00433000440c000cc0053c001000030010c340100000f0000010c0000000c00400c000030034d000001c00c0000030000c0430004fc00004000040010c00d00034070d0c0400c40000c040c030c40014c704c140ccc0100130101c3440141c00004c014010740d0c340430010c000403000300030c004c700344c4003c000400c0c0000001c4c0110500030400004000c00003000000c000403100000c00000400001000103404040011100401403000000c0c000001f7071c04030010c00c0000d0000103000000003000c404300300001c0400040001f00c1000cd40430000010011c4000c070c0c00f4005c0000f0110c000000005c5104c00c4703004030000d103c1c00000740101000cc0000f0000000000c0001010000c000003345300100700001000300004c0400303000031043c0040f004710c000410010000300050c000c0044100c00311001c0c030000010000c0000000f7014c10003c00c707100040100040000c000000000004000000400000ccc300d000040040000000c00005c004104000007410000f00c011300100304c4c03000011000c0010130300004043034440134010000c000001030c000c0000000001cc0003d005000040c0d0c000000cc01000030c0011000cc100100c003000001c404003010330000000004c01003000000000d00cdc00000000000000033c4100003000103000c000004001003000000c1cc00000c00c300030000001030001c0100310000000c4c0c3014000401103000c041000c003c0300c1cc1130000c0030c100101000000004070001430400100c31c1400004000000cc1c300000051000000c340300c100c0c00000400c000400000105040000c300004000040000000c1c0400100000cd00030000010000c00000004400400001c07440431004c30c0040030c0400000000000330030300000300c00000030000c10c000000000401100000401000000003c0004c00003000000000040c0c00000000cc031000000c004000000104001cc00407040000000c0c030033001000c000c334000000000c00;
rom_uints[244] = 8192'hc00c00c40000043400000000c0cf00c4000003cc000c0010c000000c3000054340000000000d0cc000ccc0004334050000d4c0004000000c00030003000000000c000d000100c000c00cf0000d00c3c0003100100c00c000c40000004000040334030100000300c410000f03310c004cc04403c000c04c00c0c00404003c0300000c05c000000100000c0000c3000000c0c000410c0403040c000000030000000300004000f000000cc00400c3404043c000000000010400000001000000015c0004000c000110000440000014400050f30404000001404310044c00700000f00000000f000005c043c00400000000d101033040000000c0000040000000440700330c0f4300700000404130001000430300000003c1f00001c404f03000004000044005040100040004c000400000000000cc0000000c040000044d400000030000000400030400c34100f100001730000000000401441c10001c000c704100c010c0040f34000000040003000000031d0c0040004c0100000300010c0c3001c001000000000300000300004740000000c0400d130000f0407000400000cc0001030000000000c3c000010000c4c044000000144001040c0c00031000140c400000040004c000000001c0400400cc100000003100c00400000000000c03000c00c0c0000c0005c70c040f4c030c000040c00040c00300c3c00cc00014011007c000030003010c040fc44c00000440f0000f300040003000404c4007130040c4010c41000c0000404300c0c40000c00c100000c00400014c0000400045030000003100050304030003c011c30c000c00400004cc000000400c00004cc1c300d010034c03000300c03040cc00000d0f053c0004000100000c0000000ff00034470000000400000000cc000003d130000c0cc430c000d00c30c00004000000f0f004000000003040000c0000100c0017000c100003c0030300c0c000000034000000000004000303c00100000301000c0700100040c430000cc000f00c0f004000c00c300000400333405000400100005c00030400c000c003004fcc000000300040004000c003130000c000c3cf0c0000300c000000040540011c5c010110cf00030400c004000d001000000c000c0004c40003cc0c0010c0400053030c0d03cc03300030430c0000000c00001300030c0004013c030c440c0004c040c00400040c010001000cd000000300000000010001400300010400000000030100c000000d00000d000700c00313c30000c0404c00300c400000010100000f00000140c7304c010003000000003000400c3001344c050000000000000000c00000000140c040c40000030000000c004000000000000003000403100405c043000fc00000030001030c340040c300500c3c01c00000c3010400403301c3c0c000000;
rom_uints[245] = 8192'h333400000004c33c040c0000000004300c070000000cc7c0c0cc03003050c000003cdc0400000000c10000c303c0f130f01440500100000000c3c000451000c00001040001d00140d000000d14004100005c4000000300044c0d34110003cd15000000c0c4401300f00c41000001000400400000c00004100000003003000000c305010000000003c030000430001041030cc00000007040c3000104c003004000000000c04014c0410000000040c000100dc440000040040000c01045000400040000cc000100540000004c0000c04130440033c00034050f03c340f040010400000000c33000000000040000015001c3c7070001c000c30000000c00030000104400030d000041003303000001c0030d4300d13000300004000010010700c00444c0001000c0000000000110003130c001c0041001000040430df0004103414500300000300000cf014000000410000050001043000d3c4c0300000f30010c000c0030100c41004041000000c0400cc000cc04004fc7010c340000070001c134440100100c0300010cc00044c000c000000001034100000014c00000040000f0c40c0d00c0400300043000c3430000000000041c004dd3301007070001d0000030400033c0c0c3014d0cc0c000404000050013c045d0c403011c00001303010c003c10000c4301d40c05034d000000c341444c000000004104000cc7000030000c0c410010c0c4000401040040c04000000000c0004100c003000cc330400000040333c00c4000000140005400001000403000c000030c00c0001040003314c4010f0101000300c0000cc40004000000c00c400c040001000d00000000030040400000c000040403044000000001411c0000030104c003c10043c00010c0000400c0d000000005030003003401c000014001cc0010300000f0000141300044c00003c000004040cf0141004fc00000070300000030000104000301000000000fc010000300cc0700030000000f030000d0cc40000d000100000300040110030c00000c010305040c000d4000554ccd01010c00000c00004000010000300d030400c100000c03c0030000010440000100d040003400000000004101050c070154000000c34c44030003135000000400030007c00030030c0003400000c0470031144000050101c30013030404040dd300c30c40d00040000c3000030300c007cc0003003570104101030c000000c04034001001c00301c4c1c400400c443400330f41c004000c0003c0f00c034c0c0003010000c00170003004300c4000030033c3f0034c014004c4000400c00043c400310105010010cc004017000c0000100c4c400c00d404f0c000000000400000010000000003000c00c0000000000001c3000100c3100000c0000000001010000400040c3300410d41c7d00003004400;
rom_uints[246] = 8192'h350000030003050104c000300000c0c0370000f05c10000ccc3100c111d0000300004c3000004000017c3300043003070040d100c0003100300010410000d0000000000000c03000013010c0000174c000007300005100d3d400000000000010f100700014004340000c30344cc0031310cc001100033c4c700c000004000000c04040400000f100c4010000010300c03000dc0030004003000000c0000000c1430000cc010040000f00000c00000000c000000400d0117300340dc4000000000c1010000c0434107400400140340000103010c71001c470c010c00010f000c000000040c1300033f040c00430040000000000100000300000100000000cc010f0000d001000c10100005c30f010c430034000c00000000c00c100000000c040c0100000700000000004303310004300310040104310430005001000000f4c100000000c001c03010000000334000400c1d0f14000000034c0400c0040000003c300c0000040100400000000000000401301441000d000c0c030040434003004007003c410000040f10101004034000040c0400000400100400003f0040400d0000000c00040000cc0334050c051c004000000114c300004c00c4000004000d003f0000000403c00100011040000c0c00001401cc00010000040103700d0003300c404000000003100000000001303003300034010c010c0f4070c030000f130d0000141504c031113c1000c13004001307010000100001004310c0fc1c0100000400003000000c0c140004430c030713003000040100000c4c0000c0100000030000100c0013334c00040310010004c000000c1303000c04c50340c0d003400003040001315103000003043000400300004000070000c0003374000c40000000010c000404030f43f4000c14c00000004c400c010000000400700000470c0000040054401300000011313c4307c000000c140004000c0000300033000011000c000000000c0000040000000004000044010000070c0300040c300000040031030f0307f000000c1c3414004144000400000c40413000003dc0000000034cc300011040010400001000000c0cc11000130000c1000000400d00400c000f0301040100c0000000010003c0cc0050000400004f00001c040504d0001f0304100004000c0000300000034101010000c00005070001040000000403000103040c01000c0000043040d003030f00010c00044c0c14c50030c3030c1003400310c0000400330000040400000010c4000303040000044000440c130000001c0000040001044c0c0d00c3010010000d0110cc00010000000d000003300000010300000c0130400004cc0c30000000d000000001001c00003c00c0000740000000000f0c000131c30401004c0000000500000043100003010137400004000;
rom_uints[247] = 8192'hf4400000001c000000f0000000101330035c00141334000c30c0000000000430004c0030001c0000400000000c00000c0430040c4030001c140000400000cc000000410c3000000000000400000010000000c5041c00400004000000001c0c0000003000303c0004c01c05003c30043040343004003000040000004010c0003c0c1c00000004040c001c10f010000400c500000000300031f400000cff100001c40004000000f004000c00000000c0300030c100000c000000003000304c0c300000c010000c31c0cc00000000005c3000c0001c303c00f00000100000f130c000100004103000000c300044344010003030000c000500000c000c100c00000d043000c0040c04000c000000404010303c30000000003000f00400100405030700701000100c003000340300000000f00000300c300400043010303034001c403c00d004300003000000000000001c1000000400104100044000c41030000c040030c003c000030040500030c03c0c000010c000001c0c04001c0c30000c000000300c004c1030c00300040c300040014c003c500000010000400000c0c00000000c0400003000000c301c00040c003000c4040c1400400000000004000c0700300c00000c0c0403030110044300000000003000100c040c000000000404044c0000300330001000040c301c00c00000100430d0400f040001040c1003000430f030cc040c00300000c00004f00c700c000004f0c000440c0300140000c04100040c1c041034000c00000000004000000000c004045c00000030400c3100c0700000041000000430c00c000000100c000050040000005f10c03400003000000050040000c44c0037040010000c004c0004101c0c1003000c400c013000000000000403000300f0310c00000c3000d00030040c04101000000c101000304cc0000c4c0040c01000100040300cc000001f0000003004000000000040444000000100000000c0000000000c30100030107030000c0c3100000400300c404c4304101100000040c30040000043040c40000400000cc00000003000103004001c000003000030004000c40000c040000000001d003c0000001c00004000000c040011c0100000340034000000040410340c10040400c00c43c00004300000c4f0c034100400354000000000300000300010000c300010003001044000000000040c10300040043f10000431000035000030404014100000001c100000000003000c0000000000000040000c000030000c000010300030044c0010003000000c1400003110001010004c0c03453000040c0004004f000c34000400000040000003d410000000c00c3d3014001010103014301030040100300400000000f0000334000000000000c00000000000010000040010000140000000400310f0400000c00000;
rom_uints[248] = 8192'hc001000003000000103000c041000040100000003010330000f10000000310400041100c004c300001300000000040407000001c00000040c0000040d30000c00000400000013000c10000410c0000540050000000005033300040100001110000000000000000400000500010c0d33300300010000c00003004003000000000400000100000004100000003000000c330000000000000c000000000100c0043000010300041003c0c00000030c0000000001000000000000000001000000c010404005000040000000010000010101040c013f00000c00010031000000000001050000010000010005000cf0c0f0034f3000001000000000000300c000000c41010000c0000000000140000040010000c000000001000c0c0c00001d000100000000000010010c0000c1c00f3003000300000c00c100000000000000c400000030000000000103000c0000000001010100001400000004c440c000c000000f004f0000000000000004030000000000000000000c004001031004010303000003000310005015000c000000000000c34d0001000100000c000f104100000c000001c501040000001000c30000000000010000000403000c4c010300030c4100000040000000000000000500c400410c01000003004040030301000001000101100c0000000c150400000fcc0c05000301400c0001000300000001000303c0c0c000000003010001000400c0000c000000000000000003000c04014150030530000703c000000000040030010040001000010100000413000004c10c003000000000004c00c00c0000010000001300cc000000000000c1000407000004304001d40c00000045010001000000400f01010000000c0c0003c000c0040001f00000100c41c003040c03300300c001000c004c3404000004c000000300000c0000100303000004040010034015300c00000100000f0304000300000cccc300000010c0300100000000030001c000000301010001000500c111004000030000c0c0400000000000010f0c000f000000030000000304c0300401040c0145c1000001300f0004000400100300000000030503c10001030000000100000005c0000000050c0c40000c000305000c30000000300000030c0000000041000004340c000001030c0f0004100003300c00000c040001c00000cd00400000f400ff0000c40c00400001c00000000c003100040000030000c00c7300c00300010030000c003000c3000500000000c00f0000000003004541400003000000f10f1311000104010000000400014400004000000000310040000000000c000034000000000000000000004c004000000000010c000000000100000c040001000430000c00050301000400010000010001000c0300000c050003000c0103040300444c4000c00300000;
rom_uints[249] = 8192'h441c000000000c00000100c0040c040000c00003000cc0f0000334000c100440040004f000c000001010040cccc00c043000440c100c0f010030000000004000000430000000003540000040000000000000c1000c001033c700f000000000c000700000000000c0000400030c33000000403530000000000cc00cf00c00000314f4400440000400000000440000000c00000030000c00010f1000c00030000c001000000330000404004c0010c00000c0131000000030c03440c40003040430f400101000040c0400100400040c00003400cc4004401cc100010040501000040100000c00000000040000404000010000710000c3000000000000c000000000c0000c004c00c000300700340400110c04004010000340001330cc4c0f03300000004000c00011000000010040001004000cc0000c000000000000f0400100000c10300c0000300010000c003004004010104130035004373041c7000f000c00000044044dc000c003340c004444000003c0003c0c000000c40000400003000037000003c00000000000000000005410000100300000700000000c000c10c0000040000000003340040d0cc040044000500030000000000400c00000000400000cd0c00c0c00333cc0100000c0000005300040300c0004300c041004004000000040001000000c03000440c00c40000c0c00000003c00c001003c40000c7000010000000000000000000c01000000c000cdc00cc00000000c000c000c0000cc00100400c0440000000003c04300010c013100000001000041000100000000010301000001cc0000010000000003000c0c0000000000c0000004000040403043000047003c0003000c44cc00ccc000000000c01000000c400cc400c000000000004400000030c0004003004001000403000000c000cf044000cc03004c0c000c0c3401c040011fc000c144034c4cc0500000000c00033004c0c0400c0000000000c000400000040f000000030040000c0000000400400c000d00c0c0000c0001000000003040040000000003000300000000000ccd000000000040004000000000040000400000c310000000000000000c4300000c00000001000000d0001000011c0000114c0000000000000d0c0000000000430c130000000d0003010005000c000400000cc10c00007300001004030001c0c0003000000000d0000000000000c0344d000000000c00000014004000007000001040004010c00040100c40cc0000000000000c000000000000000344000140007400c0000003010c00c304c004000000003100400300030000000040000c0000d000c00c0140000000000c0000c0044000030cc0000030000000000004000400010000c100000044400c00c130000000004400cf0004040c000403000000000000000c0100000f0003000400;
rom_uints[250] = 8192'h41c00000000c001c40400c0000000040004040303000000000400400c50400100c000000c0400004f400000c00000040000c00303004140400000000c0000000300c1c000c00000000000504500cc0c401c00000000000c0000000000400d00000000000c0c000000003c0000040334000000cc0c03000000044443000100004000cc00c000000100c40000010000000000000000000003000c0400c0004cc40f000000000030400010010040000000000040000000c00000cc0000030000c0003300000000c0400000000000000c0000cf4c000c0040004cc0000003000c00c0000003000000000000001c0104000000c000c040000000000000400000000000c0034040000000000000c0000c400040000c0c000010c00000c00010440c00000001000c0d000000000d0300410000000000000040c000010007100c000000000000034000c0000400000c04000000440000c000000000c0003000040000004000c00c0c0400000700000000000003004004000000040c30000c5000040c040c033000c00000000450000000300000000000000000c00f400000000003400404c000000000000100000000000000000000000040c000000f000000000000401004000c0400000c0000010000c040000c0c000000400c300003400c0040000c000c00500f000100430000c00c000000000000030040000400000000000000100000000c0100004000001000c000000c0141000c0100000c0000004001030c004404000101c000c300000000c0000100c30c00000000c0c00000400c0000c000000000000000000c40c0000000c00000430003000c3c0000100000100100000c000410000c00000000c00030000000000c40000000cc30c00000400000c0000c0c000000000c0000000000000501040000000040000c0050c040000000c00000100040004c000c00cc40c000000c004100300c004000000d0000030c3043000000000000000000c0030300000000500c0000000100c0400c005004cc00000040c10000400cc1c00040700c0000c10000000000c50000000000000000010040000000301ccc4000004400000000000000000c00000400000040000c00cc0400000fcc000003000340000400000000c0010000000000000000044401cc40000c010000000000004c0051c00000c4000000044c0f0000c70000010003000010000c5000005000000043000000000000000000000c00003000003000000000000000c3400105030000000000000c0300000c4100000c00000000040c400c04000000c0c0000000000c00000000030000043c00c000c40700000100c000000004000000c0000c0000000000c0c00c00000000000040400040004400c00040000c000c40000c000001c00000000f00000400400c0000000000f00c00400300c0000000;
rom_uints[251] = 8192'h30000c30000000c004000011000c3000040010100c0000001340030000000004f00300cf00000001000c4fc00c0d0034004004130c0010000f30047c0d0400000000c40c000c000007010c0004000000000000c0030000400004000104c0000d0003004040030000000000010c400c04001053100440000140000cc7c0cc0030003100000040000004040d00000c000000040004000c040c0500cc30000f00040000003404c30300000001000c0c4400dc01000c000c40000000000000c00c00000c00040010300110000010001000000c0001010c000101fd0c04010500c00000000c0c3300000dc1004000140004010c00c00000000100000054040000340034300403004404013c0005300000003c0c0404004f00040000010001400100045000000414000c00000c00c004c40000010000001c03004c00100304c0170c00010c0000041003700004f040c0000d0000030000400004c411404c00000000440000c444000433000000f000000d0c00000000000100000c040c300000000400040010c000000030000d00c000304000010000000c00430340040c40000c000fc0500c0000c0000000cc000d01705100040000c4140000100cc00000444c44310004c700d0034004000000f00000010c4c0001073004000433100004004040000c0400004400001400c004000c000c1043000401000c400040033001c0440100010434030c00000c30c0040000c001c000000013040000004c114d000400400f0c0000033c0cc00001000040004400074110404c003004010c0000000300c0000400341404000c0400ccc004c7c000404040c00003004005000004010f30000040040c0f00001000000030000010005000000003fc00c401000004f00c0030c0010010c0000000c403c0c0001400000400c01c004407300004040443040f40c40c070030040000c003030cc10005000000c000000004cc0000c400004000030c004000400300cc0030000000004c1000d00434000004040000c0000000130c40000001c00404000000040d10000000040000f000c0000700c30c400000300000030104f0003000000000f000430010010c04030000000004c0003d0f0300004040000450104d0f00304004000c40c000040100cc00000001000c000c0040001444100003100000070c3c000404c000cc000440c0000470c000000000400000000700000d000040040000000c0003000000400c030c0c0500000cc00c30400000104000400300000000074c4010000d140040003540700d000c140300400c0030c4cc0005040c04030000000c010cf004c30004000400100000000300001010000c041304cc40000400d00c04c000040030400000000c00004c0400c00400cc0000000000000c144040000010700010300c000300c404044c4cc0c01000000;
rom_uints[252] = 8192'h1f0c0c00000104030000000000000001003c000fc30c00041d100c3000003541110434d000040003001c0000000c07100007010104340f34000c110103100000010c0041100000100100040c7000c004003000c04c0f0000000001003301303c0000001317000004000c010c04cf040005000c04000c0433011000000c03000c3ccd0000100000000000000c000000c000000000000000000003000d0c1c0001000000000331040004311f00003000050004c300000c00301043000101000040000000030000000107000045100100400000c01c0000040c0030c0010d0c000000000000c00003000001000100c1000030001000040c000000101c001c000030010000304000100100000404fd000000000504011c10010030011c0c033c030044000000030c000100040c00000003041c0000003000030033000103000014010c000010000003000000000f340cc00000000000010c00f4010f3000000c04c30000001c4100141d01000003037030000010001d000000000001410c0c10000000c0010011001d00043c0000000050c00400000004000704301c003000313000000504000000041300110c0300000110300400f003050100c000010043003c400f1d000c0c1c030004311400000000001c411000103337000c0c0010000d000c1011000011040c0c00000004001f03010000003430000003000000000004c40000030000c330000c0000340c04170000000fc0140f0000040413d0100150c400c00d0c00430c100100040100100d0c000000400c00100c300c00dc00400001440c0c3000000fc40c030d000141400c0c03100500100000040040100c000403410101000000010000001d000c3c000507130000cc030100040400cc0000000055011c0004000c003c0c0c031c00411c140004400fc0000070000f00001f0403300d000f33110000000000010c03000500540c00000c000f000c1c400c010104003404340100000100000000070cf000000010000000040000c0030c0100041c000000000005000001040c040000040c000003000c00370000000000000d0400001c4c301c1010fd0f00000030003000000c0100004000000c000000010100000007010000013000000c30000400c0000301000c00000c010000000fc0c3000c000c0000300d00000010040000100c00000000000300040004053f000000000010331003000000003c00300c300c0c01040004d30100010004000000040c111c0c0004000001000000030000300c011f30040300000c100f00000004003000040000000f00000334014500110c3f00000c30010000000000000004010000000000003714043015f013000007004004000450000300000100c10000300c040c010c10c0000004000c04001c040001010310010c0040000300040000100011000000;
rom_uints[253] = 8192'h40000000000000003100000300011001000001300000000000001000010000000010000d000301000001000010010100110303030000030300041100000300030001011000000000000001100000000000000003010000000000010000100300010100000003000000000000000130000100000000030003000100300c0100000001040001000000000000000000000000000001000000310304010001100001034000000031c11011100100003300030003030000000031103000000000301300000300000000000000000000034001000000033000010003010100003000000000000001000300010100340030000000040001330000100000000303000001030403034700000331000100003100000000000000011300030001133000310000000000100003300000030030000300000001000100000000100013010003000100030000000000030000300000030003030000130030c00103c030000000330000030307c00000000000000300000000000003030001030100040000000000000000031030003003030030300003041f0000030000010000030100000100000100000000300000000100000333000000000003137400000000000000000300000003000000000000c000000000000307001000000040000001000000003030000303007001010013003100000003000000000000100003010000001301000d000c00000100000000001000030300000030030000033001300100030110000003000c010000000000000103010003000003440000000300001100030000030300010003000000000000003300000007000000000000030300000000000100004104030000110040000001003101000001001000330101000000030300000010000330000010010100000434011000100037010300000013000000000c03000000010010101100034310100000010000000001100000000103000000000000010000030000000000000000000300000000110300000000000303030131300000000000300000000000000000000110000000030001000000000301000100030003000000000300330300003000030003011000030000000100000000000013100003000030000013000000030000000000000030030003000000000000000000000000000001030100000000100000000303010000000030010003000100030100010001100000000100000001000000000033000004030031010030070000000000000000001300030001300400001100010300000030000044040000000000000100010003000000000000310000000000030000001300000000000000000000000003000100000100300300010000030300000000004000003100000003001300000000030010000000033100000000000000030100000003000100000100;
rom_uints[254] = 8192'h40040c1000000044c0003000000000000c000c00c0000000cf0044000003000400000000040043000000007000000400000c00000004000c001000010c0c4100c50005040000030c000000040000040100000000c70c000c00040000400300003000c000c0001000100c4000000000c000000000cc0000000c00000cc30c00000000000005000c000000400c00000000c004c00c000000c310040c014000c000041cc4404d00000c0000040c30c400000000d40c400000030c0000000000c0000c03404004000400000100000c030100c4000cc40f00003c00000000000000043c0000100400c3400104300030004000c300004f0000000300000000fcc0000003350400440004140000300c04300000000c0c00100000130010103000000000c00040304c00000c000d000000000004000c000001540000000000000d300000430c000c40000c04000000150004000000c0000c04000c000001040c000001000000004c040000004f0f0c001400400c00000004003000004c0401000304003000c40000c000000004000c0c00000000000000000300400000000c00350407000000010c0000000004440400000040300000000400300000c01c01000101c014000000041c000004000c0000300004040c170004000000000400100000001000040000330710cc000c00000000000d00000001c00c07000c34040404c0cc40000c000c0000040c01000c0303000440004400000000c0350c0cc000000c0000100000000000c1000f00000000cc00000400004300403000400030700403c0010f0cc70c0000cc0000140c0000000000c00f00000c00000700040f0344030030000c00000c000000000000000000030c0f03000c000dc000000000c000000cc00c0000000000c0c000041c000003003010c00300010000001f00300c000c0004040100000c04034c000004dd4c0004043000000cc00c04000000040c0000030000000c3000c00c00000cc0c40000030f00040c0000000030d400004c00000000040c0000000000000000040300000c030c01000000c0cc000c0040000000300004c0c00300000c0000003c00cc300c0041000c00001000000c00000430000000040040000c0d00c4043c00000000000000400c000400c00400040c00000000003044000000000000c400310c0c3000040440000c300c0000000400c0000000000000000000000004000001040000c004400010055404000000000c00000c000000000000000c00000c000c0000c0300440030c00040404070000044040000000010000c00100004300010000001100c010003000000c00000040000c0d000030004c0030010000004000000440000c00000000cc0040400f000004c00c00000c00000c0c000c30000000300004000001050044c00000000c04000000;
rom_uints[255] = 8192'h10c100000000000c0340040000000043cfc00043c0400000004470000000f0070000003030100000004103c0310000f03330d0d000003105000050300001c000fc0033cf40100000040057400000d30c01c100100410c0430001f30c00c03040004340310001000fc00004000c000430004040c0333000000000001740710000c1cc000047c1100c00c40030d00053040071000c0040d000000000c0c000000cc0c101000040700100c00000011000030040f1c400101000101040c00100f000c01000d0c0000c34c0c000c0c007df031010c00000503000c1400c0011304030d004000330000100000000d431100001000403530140400000c004400000000000033000c400000030c03000c00c10cc300c303000c50100304400044004cc700000300000000130000100003300300033050c030c104000000501400040000c00c5c3140100d30030007c7c03010000c0351000100000000000d300000000430000c0570d14f300c00000414f10000000010004003000001011c030f000544c3403404044513100c3c5003000000040c0c00c040000d0110000c14000c10c40c5df3400003c007000c0d000310cc3000000000010c000f004400010300040144cc5040101140300000000007100111500104004001013030030100c10c000310c1400010057000004040c40000000c340c000001301030000c0000000c000f010f0f34300000030100000700c11c010144130044001404000003310c00000c131010000003010000000c0700714000004000000d00140300400010034001301c001d0300d40370003d3000c000010000014000004c10000005000004cc400100000000040704000000431300c0003c30410054c0030c00030000001003300dc3000004300700070c10f0cc10154c30033010043c30000c1000c100050cc0000310000440070000011000cc1100000c010c000404003004f30c03c43c00000c00d0000100000304300003003000c10040043f30000003100113100f033fc14010000000100c0c14c00403000000300004000cc0330310040001700100c053c0000004030c0300040c400000c00003040000000000d0f003030000cc4d0000004c1d300003010000000c03000000003000013c5033cc100000001010340f003000100434000404400c000c4104043107c03cc000000050300000c500000d00c1001003cf00000000000c0404500000040000400c43000030000c0000000001400c3100c30000001100c100f40cc0c0014c001470100704000d050000110400011c00031414000cc010000000000c0107000cf0000000000000000f000c0034000004310c0000c00dc300000c70003001410403101000c001c00c134001f70001000000030001440400004301010035000040043000000c0f403c17430000000c1;
rom_uints[256] = 8192'h4cf14004f1307003c030104400c1000cc300c4003001f00030f0501cd0f010000004007044700000c1400137003003000010001040cc700050c0000ff000400000cc0040403000c000000050304430040cc00033030c000104dc00c0030031000400510040040413d1000044040c04400143c010c00110cc0030404c0440103005410300303000000c000c00003444c0300000f00041433fc03c0000001000000000040cf0001000704f000040c0003000f0c030000f003004c30cf034c3003034400300100371314c0000450030f0c40140005040dddc0030001400c0034000c03440013040003000f000d00000005cc0c0f000404000400030005470001c1030310070f01070140000040040f04c003030000c0000c0504410c470c3303400c00300007400c0c040c00144033301d003400330c000300000407073c3d04030404f705000013030000070500043003510010033c001500003cc4100430440740010c00140130c3c00c0000050004c0030004000cc3400d00400100000000005f007104030000043030000010f343c433030c0001c0cc04370f000003300f400733f000140500f1040c003000000fcc3f10040c44cd00c3c000400104cc000504000130c0401300000501007000110c440400030c4f1f400c4cc00000cc0d371c00c03c000c44c1440001400540030055c303015d010c044500000040c3040d0000100001000c400304000f10cd0300c1c030000003005c004d7005040141070c0ccc03c70f000c00000131440c00c00f10c70340030000400f34003c00134000050405000c0030030c00c0000000c3030304000730000513440000570c004f5004000c3004000300040403f4cc04000f1000f00c40000003040000cc00000003f00d00c003000047c330511c4fc3001057cc0300c0100100c4000414335000cc040c040c11140c0043007034540403000c404004001040c00033d0c0c3040c0c040000040010000400000007000c0000500100000004040dc30c0c430f0c00000001000300500304000070071403400440305c010c3000010501001000000051000d004030031403c0000301c011004010000c0030040000cc31000404c504cf0130003f041c0303070f03c30000040300100100430001c0030103040f40400f140100014c0c010010404fc50f510c010001010c00000f013c0000004740410003103c0c4c033300005000010100013013050334000401000c000000cc01000400cf0304000d000c040001030017014400f0544c0001033c04f304ccf000070c0000c5300433400cc004370c00001c0034000f3c0054035700040000505030000c50040003054310110400110001010540000ccc3f0c03000c000003100f0070001007000001000333000340000000300400c000070c0000cf00100c000c00;
rom_uints[257] = 8192'h10c03000050d0000050000c03040000130000d13000c00f401000010500c000000cfcd300130000410d00d30000300c0030c003c013103001c00c04040004c0100003103003d0001000d000c00000000000000c0103c0430033ccf0710c0c570cc014c000000c0030000300000c1040400040c04000000003c7000401401040344031301040004100000c00440001034f050043000041100c000000300040040330000000030c41130000c00040031300010300000370f100000000c500000301d1100000100310000044d0cd0dc3404000c030040000f0c4f5c0cf4c000040c00300c0000001d004c00033f433c04400f004400031030001110000000c000fc00003000c40c00730044003c010000001010000c00004003003c00001fdc00f10f03400050000050f77c011f500fd304000dcc00000c000011000c010414040000c00000fc410100ccc30fc0340030001cf1400f300004c0101d003030c01c000c00004c010c000003410030001c03040000000010000030cd3c000c0cc0f0043040004000c40400c0014000cc00007300030c03030c00301c30407500734400c0f0000000c403000c0004000c500c40c000000450c004003000c000303440000c30030100413000301000001010c0041c340c0701c0000003c4000000f73c04000c3013000013403314000444000c0300004130000050fcf0303004100c0c1454004c0ccc0c0301c7000100077c0043000c00013000000d00004000014c7003000c0f00100004c0000f0000000010000000004c3c000004013c0cf01001104c000c400050001004100000300040000001d000300f0040404000100010003100000400000c001313010c000ff0040100d00400004400c00300c00004c104010c30dc0110710c0040000c000f0000cc0c000c04000f0300000c41c00331cf43c01040000010000c0000000010004030d003d10c1000300000100c7004c0000c000003c5000001400031000c0000500000410004000003300c04000113000140514000040c0c004010001000340c4c03044033c3300100400c3043c0f05100c000c0c0041c0cc05410d0000cc304004003c00c330530f400001714004cc3000000c00010f01010500100c00034c30000000c43130c0001140010001030400c00001004c440300300304044000000117710000005cc04000f000c51000177003000cd4000cc703c0000014000f300041033c000570030513030c03000005000100510d30004300d0f00c01003005104043c0c001f1c440710004f00c0c0103000000000c40100040104540045001c0000040c0c0001100000101013000140400c0001130c11ffc003003000c101033101000c00000000130000013104001c4000003014000150001d3010003c0304d0045004003403000cc00004400d400000040;
rom_uints[258] = 8192'h5100c0000c300c00000c3030c0c00700000000040c300140030c40000030300c00c0000c00fd0c0001000c004c000004c0040440100004403100000c040000040c00c30001c0000d0000031f7d004140004005c3005001c0004c134000000c0000070c3d010000730000030044c030000003030000014140000c0017040000130c000c040c040000000000000000000000710000000430304400000c0300000003000000000c00c00000c0000c17c3110145400000c301030041000404400000340c40000c000000c00c000000000000030034c0101000004504c0001440010000c00c000000030000000041c00c0c0344cf0003140c100c004000c000000010041c000040310c040400410003c33000d001000004300f00fc00000004070c043404000000330010d301c03400404303000000000400c30000000003001c00304c00030300f00000000c0004000c000c1003c03d030100cc0004700c004c0000010000c44f0000c4c04c00000044000400c03400031004d304fc00034f00000000c000003000004044c00303003411000c004000000043004c0000c30030000c000f00004ff0c0000c00c000010f000704410004c30000c0c34cc0000300000000000fc0040003410013c0c00000d0000f00000000010c0340000000000000000c010c33013000ccc0010300000c0040c0011cccc0d000000c00000000041041000141143001040c00040c0d000cc4c001003100301001000d0c3401cd000001030000c30c4540000040000050000341040c3001000000043c07030440000300000700000c03003c00004703000cc30300000d0c04000c0c40110000000004000100000c0c00407d00003c071013c00101070007000c440f0cc0310040000341c3c1000040000c0fcc0444300c00430444cc3c000030000f0000001c500004005c0c30307c0000040100370c0001030c05340000000c00c001004c0c00010040000c0103000001004c00c3c00000000000c001c0003c7c4c0400030c0400000170000000040c4000000010c000c003000040407c030c40000000000300011c4400000c303c40000d40000c1f000003cc43000d4110004c00000ccf0c44003000010000000400340040440400400003c4000330c004c000000700310c01007c714005004c030c070000004400c30004010c3414004510014400c00000000cc3004d01f00c3c00000c3c0000400403cf01003030040040f0c3dc4304400013400000404c03000001c0000000040040000000000041c0c00000000304010400001c040000000c000c000cc0000004000010400c1c0004000500034000000d00000000304df10c043307000cc30000030000000005c003440040031000000310700501030040c0010003000500044510004004000000000010040050005000040000;
rom_uints[259] = 8192'h500000044000031000030310000c05303cc0001031110000033010070c00c40000100001cc31000104100033100000c000000c04c07000c00000300010000000500cd0000d0000300000331000043001000044010000f000410000000c030d0007000010014003000c0c10030c03073000003c110030c000003001c013070000000030010300000004300000000c104000000030000000101000010300130f000d0000000c00c0430000010530300c10000000300001000034500c013310c0004010000c00001000400c0c41010034cc000000c50000100150000000100000010000003004000010000001f034113300010c043410400010030c340430003000000cc010d01030103030003c04f00007301c13003c4c1000130000400300f0000000100c000c10003004000010000000003040030001030710000003400000c303000040040000040cc000413000100c000003700c3c00300000001030000c00010c00103000330300dc4c01107000004c30040000c0043c0c3000101000000000311030000c30030100000003000000100c0403000030c000c10400400000300d03031010c0c0c000001000000d3500104040000000103000410000050d00101c0034c000303cc000130004000c000c030101000053300000c111300c000300010400410100000004030400030030130030c01000100370400014003300000100000040000c10c4304000130c40040310400301000000040c043040400c110c00000000c04040000030300331000400035000000000000c04300000100000d000003000c30503101030003005003000011000000000f0000410100c000c00000c3040c030330010010000000000340010540030043003003040000000000000000000c400000004cc10030401c000000010f004c4004c000c100004001d4c300d30000d0c1f0000103c03730000035000130500103003000007000c1030030c00c300000000003300000030003000030000030003300d50000000143003041c00031003c000003000000000400000000c000d03c0003000001c1003300c0000031001011c110c410001000000d0000110003000100c10031700001310100000000001110010301403010000000dc000000c00fc0100140010003c000000000311100000300000000d00400100000c05000d000013400013030c0000030031c00c0c0301c030003c0000003c00000303000000007034000003c0030101040c0310010000401c0001000300300000501001103031300430003000300000d00000035310140407100000000010040c0c0004103100c0000000030000000030003007001000300301000003c3300000001100004000000030c000030000000313003000100c304000000000001001030000000303000304c000000000003300000;
rom_uints[260] = 8192'hc04300000140000003c031000141cc10cf0140040000510000430c40c0300c11000034440004000000f000440500004c4007333500c03fc5433c1000030004040000000d00c00051100000d3410040040000404003f0000000c7c300c1043100000c0304f300c500040307c0030c44d0004c000040c0100100000c3cc40014004cc000c010d300c000100040c0400404fcd0314000100004c0400300004c00c001040c0000cf40000001034003c44c3f3040c00000c001700000004000040700004104300000c4cf704c003cd01d0040d04fc1d000dc4c00005000c744c301c0003000000100c000f0400c0000550f00cc400400007cc0000000003000000000c000c0c1fd00cc01f010040307700050300444000ccf0000d00000001040c7c00003c0004d3400004054c4c030000010c0000340103fc70007c050c0c0030d00000031050073c400300300ff5f11000c0cd04000000cc0304440031000000cc404c0c4c0c30f400040403500f000400c0000c000000c51cc000000300000c3400000100700c300003c0000c04040f000c0000000040000004dc700cc3000100040400000400001cfc0c0c100000405034000c0500f000400f3000f3400300000cc104c0010000441c00c03004500cc00300400013000170000c000004c00040300c00000100c0003c0110000c0030f40f100003c03c00c00030000000054005c0000c004033304003011004040c3c1004c1c34c040c000034540c0c04f00c4000c5005c030cc00d1000000007440c1c40000000000000040c100340030c001c430c0c0000470440c0cc43c03c00c0c3000044000c000ccc0005d00010000f04051c00003004000c103c0d03c00c45000400000c4cc0050c000cc14c0c0f00000c047004000004003c0c40c405400fc0004501cc13000110003c430ccc4f034d0000d0c000cd04040033004013c30003f0c04140cc000000f440047d1c0003043140010000100100c030000000000c00000000c00c40004314003000400013004050000c0000c000c0001007c007030430000407c03400040034cc00401100cc01040001010cc450104310cf70cc00000c17c04041d01334004030c00c5001400443000000170000030c70c0c30014000c0c44500003f000000403410000cf7d0000400c000000f0500007ccf0001000430ccc000411010c0403f040013d0001c0144c0c340400004c310c304c000c0100000c3400000cf0c0c00000300cf400100040040000000c0c0033f00c0c0c0105000001040ffc300000cc00004c040c00fcc0040cc100010030040c00400c00c000c00c01300033000034f00c0100c0c0010f40f004c00f440034000000000430000c30000c050010100c4cc000400000fc304c000400004001c0401700300001000000c0000c330d00030c000003000;
rom_uints[261] = 8192'h41000000140001c000d40400c070cf03c01c400000000000007344c0c50000000d10c5001000003104c000c00c0c03c070c104000000c0c7030000000001004010000f030000040000040c30c004c03100000cd01c001000150400000004104004300133000003330040000003c00c00c7c0000d00074000400413d075c50c0313fd040105000103030000004000050c0041000003c0c1c00c010000003031c0c5000003443430c3cd0030c400073c031c0c40c00040c003730004c00c400000c404c314c001c0c00c000410000c3100c00c04c0c04000c3040000040dc00c0c0400004c0c0d00001c0030110c004010400030d37c0000c3000fc3340000001005cc0000c0430000c0010c44c0000000003c0040000400000000000343000d300004d00300d010000d4ccc00000404000000000040c4000000100330cf4c000ccc000430c73d40003000c4100000d0003c0f45c43c301000f005001000cc0d0004044000c37c30400010000030c4c04010033410100013030040c0401c130000c040003c0400040340004000c0001c3c000c0300000054c001140300000004000f503000cc300cc00034000c04c010017007c00004530c4fc0401400011010c000c00004031004000c000004f000000c3cd000c304cc000c10cc0003cc4400d400414c30033000400005c134f700000c400c13c40c00430300c0003304131c5c0030101cf400000000000430300004c03c0000c300107c0c001501c3c300c0c0000003c3005000100000070dd000041410c400000f04304c40d0000140cf04037470000037000c0f041000100c00000005c00000000fc7c10c001c0401000c04c30cc004403000404000cf10c1107c00330c01c004c0000d0000300040d000000430404000000443110030004000c034400c00440000500000035404d0041f0070cc7f003c30f00004301404c3030f030d14130c30c007cc00001d0040040c00000c4010000c4000000c010c0000000c004370014c00c000000004500c300011d00000c3003010c000001000c4100000001010d00000000004000100301341000100500ccc00cd0110c0440003c000101330d11f13104400043f00510f3400714310400003cc4cc04df70300300000c005010340040010dc400000c03001d0c0d0c000c0300c33000103400c3004c0000003010001404430000000c00000000400003000c01000c1c0000000300400400014c400100030373000001030504c000040c00000011310c030004004000c000001d0030005030000c430410c000cc004300300c004c04003000305c304104004c400107000000dc34030000c33000000011040043000c0040437c04cc00000c0c0000003000400d04000c000001400c744000303c340000000043040c33010400000001cc100cf30100000000004c;
rom_uints[262] = 8192'hc1400000007000000000f0c0cc0340101d03000300000f0d00300d000303030000000005111c0040071010131101c414cd0000040c5000170d000c00000000000000141d00cc04f00000000cc300000300300100044c0703000c14003004010000000cc000100c00000c0c03400c0000000004cc00000c0f0040010404303000fc0ccc040c04000000000c0300000030000400000040043040000440430400100cc303000401040400110000000400c000340000000c113c400000c400030000000c1c000d00011c1031001c0c000003400001010cc430004500d1133003400401000030cc0000000004000700c0034c033337030d0d0010100000110000000030c10100004c0c041c14710cc003000c04000c005441070030cc000000700c000000cc0040150c03003c0c43030040c001000000c0040000003c3c0000f003000c01000000011000c0010040c001c00001014f00001111cc0070011c10007000cc01034f0411f300c0001000d03c1040000441714007730300d10c31030c1000043c0c400011003100040c000c0040d1070077000000030000000010000c00c004df0000000c037000000000c10c0004300000100c000040013cc70000003010010300030c0010000000000030c00d04410d01004300cd030000c10000c30c0f133000330000c33c0000300c000c0030100f00dd0300431dcc00004003003d7fc00000410d0140000341c0030c000001300100c0101ccd730000000c4d101d0c30044cc401444cc00000000000c0010c0001cc000001c00000c40004f000000011c40cc1470000000001400000001000003010c000000001103c1030fcc30440000000031c003dcc04cc00511c4300c00440c410000304c0030c0f040000005cc0c00000000c0300000044f3c0c000040000c7440c0030c000000c00010000103c040010031500000034001dc1004c0434040c03400003400c404000000001070400c00c00000004430c000100000c0001000d401ccc03013130070c4000700000000c004c1040000000030300c00c14000003c000c00000003013c100000000000030000300c00d34004c00005001c0034010300c000cc000c0004c01000040000000003000000000c1c00004000004104030000000001000c040c34040dd0300c5c10010000400000001013c000003000040013000430000000000cc4340c030100304030c000001000000000070001000c101d00410000014000500343c004c0000000000d0001f00000100010147000c3c0c000000000c030441c300040054010000d100001c01000000050c010c0011c10c70000c00010c4d0000400004030c311cdc0c04000000000000c30000c00c330700070c0000000070004c3344040c04003c00014c003000004000400047013c0401000404003050c00000000c;
rom_uints[263] = 8192'h44c00001000c00003cc41000c000003330c100c1000c040004030c0304000c100000c70300d00000c0103300000034000014001c04d301000000c003400000cf040300c400000c0c00003c000000c00100c410000004000404d300044000015000c010000000000003030000000000440c0c0000c0100030040303030044000031040011c14004000000000c100100dc0c0004000000003000700c00000000100100010003000000c000000c5000003000000000030c03000c0000044403c000011003100000030010000c0000c4040000040c0c41004000050c03105000300f10104034cc0000cc103001340030c30100c40c04000000004300c000000000000000000014333104d30514c330300010c0fc007000000001070030303430000005c3000c000c400035443c040000004401c01c000000c00000000001cf4004000c00c001c014300434c404c03040c00000c0051117005c1c3c000040000c00c0000c5010300c03074010c000100300000c000c00040c040f03130c0040000300000000014030000c01000c104000130000000300000f004c000000000004000030cc030c000004000400110030c0000401010c00000310000003001300001fcc044000c040c030000c4400c03c03400c030000000000000001f0040c0004700510000000307007400000430070300304000c000000000000000100300c4000cd000c000003400100c10000001050c1dc0f00003300cc0004300010cc000030cc0500c0cc00400110004000043c000004104c000031c3050d40003400000f0c10004c00c0040000000010000004003c000010000000c030000c000c0c00000c0040000003f0000071000703d300000430c000c71d0407cc140005c000100f000303000c30000000000c1004001133000c7c0f3000000103000310001f17c000000c0c0000033004010d00000000000413c04040000030c0c00000040c040000c430014000000c00003000000000000cc00000100011000000c00444c4c1040c0c0000000c3cc0040000c404c0c000010c0000c40300000000f0004001c00c040d00c040000330005cc0d00400703300cc4134d010000000400400cc0000cc0000000000010fc100000000ccc001c00100031c4c040f00010c000c00000c010c0030c00c000004300c300c000cc0f04510000c014100440c00000000000000003003d40000000000c4103d000410000000000c0400000010c00c000c01000001000c300000000300c1d4000070030c007c131c010cc30110000000040313c000000c000000011000000100c000000c0c0000c0030040050000003440000d00300000300101c51c00100000030000f0000040000c0004010d00cd100d004f1000000000000c000007030000040003303001400000040030fc17000000fd0000010;
rom_uints[264] = 8192'h5301300133c04f34300f03ccf004c04003c040000005400000303040c00c400000cf4340345000010d00034c0040c4470340000d0403c010f005040401c3cc007000c0014000400400010570000cd001c500000400f10d0030f000c000110100c0c4110f400703000000c0030540033000003043050d030007010073c00c013f700fc1000dc003f0000000000003171007300000004003c043310703130713d7c00c01c10103100030033004404005400c43c00004c3c7c50c3000007000003300000d33c00045000fc0013000000000400000034c03c00c434001c100434010c01001f30f00000004c00100cf01cfc04c01000c4c1100000c0013410000040000030c41cc133010034000cc0030000000c0001045c0000000c30cc4003000003003300d0c010c000030cc004fc050fc01000007300400c100000003034004c0000d00700c0300040030c1c1044001400d0100103305451c00700474c040cc004074c00100700d0301c13734504004f00447c503c1f035c033303130030404750403301300040030c000010000013c101003050c4400000433c00000430000100030c1000f30c730034001c30d040100c700000101310100000d310044ccc04100c04001c1003000004000000004c00000c10c00c00c00300100f300000530f000000c04043000014d00c00031300301c0110010c4700004c1000d51700043f041c03f03400101004000cc0c00004c0c40000401300f300003d010f7007330c00003c1010004030100c0001031000cf003c01c0f053c030005100c000003010407c0c30000004004f4000004314370000010000004030000014c0000c104c73000033004c4030300000c00004c000301440107c0c1004000c0c05000c00003c000003440054000000500f000051700103d004141000c10f001503040f301000401000000f0400c0c00430ccc0d3000f3f0c00044014c0134070c3000703000c011001000000040000000040103010000011c0544030c5c0434cd010000cf00c30003c400000d0c000400004c01300004000140c00c100000c0c003f3104103050000c000533c0401011004cfcf40310030f0100740000c0000d0c00f3c4004ccd300010000100003030140001c00400000d00000003c41000007000004c0000cc3300000000100c00003f5043300000030c40753004000c0013030003000500c01100031000003101001040c000f00010cc000c10f00c0030000c0040303350300001000000310011040c0c000001415404c01703301c00fc4001003c0300400000c0000005d517001004c00303011300c3103004000000035000000014105000f000c000400c003c0c000c40005000040000000c10c03c5054001100143cc100c3f50c003f1000033013000404041405000c00f0c01100000c0c0400400000;
rom_uints[265] = 8192'h703510cdc0003000c003c01410013001cc31003110503c000100d00301005040c000000000100000003030cc01c000013c00300501000c0130003000c000cc010000d43110000c00c0030100c00410d031c0410703c5100c300cf01000304c40003c01330010c001000dc0000000c00010100fc01050c0000000000010d400c3c3cd3130300000100300000100010300400000c003005000c000f00344300c10000043000000304040000031c130c13000413cc000c300000c4143000040031000400000f03003f0010000c000c4c4114c0000000c40037c3d010d000000000003c000ccc000103310030000000400f14030001070000cc000f040003003000030003110000c70001f300c4c3500004007500131000170cf0013030001c0c0000410f00c4000103c3010000c1d4030d0000100f01130c00040dc033343c0000c050f3000301c004500f00c41f040c30040331351000c30401031f011000400303000040cf10030000c30c0033100c330017403c00301000000010001c041f0301000dc0c0d00400004300dc300340cf0300c04c000000c0c00000300115c004d03010003f1001c00337330000d000003300c43400111000000000030c1c0d000000004140000c4c0ccc00c317000000070c000400c0433c04100000f300000f00000000050010001003001fcc0400001000c303401f04331000010014df0030170003c700031005000440013034004000030030fc0c00c40300f040d000dd04d140300313c33300000d0c00031114400103c0000c030c00d13f00000100f0000301000cc7000303033003010c000100001400c00c300f000004d01305000c030c0c00300c00f300110f1c00cf10000c0000004d11400c4c40001404013331130cc031534c0300fc00c1c033001030fc5dd0001453c0143c00f103004f0000130330400100003010c000310400030c00001c01005040000f10040cc0c10000004040433005001300c0100f0300c401000300d310004110f3000430045004f000c4003c040f0c0034000c0f0000001c003c0010c30c0007040c01f0033400000003011000751033c41000000c00c03f00c300100005c30cd04070740001333f100303000010c014044cc0070403010300001cd400000cc10730100400f34700043003333400001f0000000c0003040c310c400001007400000033c003f004c3000400010f300c0030cf0f03c43110340001c3c314310c1030074500c004f300040010c73040000000f10c0010033303c11000c30000101103c330100400000141030f443c4013740030004340010133010003330c4100150c00000100310307000053c0100004013c003c0c000d3c033c00000000003400c100000c0001cc0440000c0000040f0000003010000c00c700030000003004000040014ddf00000f03;
rom_uints[266] = 8192'h1c00000c14d0430004300000c000300c300f10010703d0000000000000004c0004013f34cc7400001000003000000341030c0040d1300001300c000000000004c4c4c3c0000000010004c004c00c3000000000004c4010010440070001343c500140000c000cc4c1104c00f4004c005c0000f040c00c07000c0000740c00c0c003330c5010000740000c3000100c3c1003000000000100030c000040030d00453300040001c00500cc0000100000000fc0000000004334700c4c4000d10030044000003c00003000040000300310c40000c40100001c00001040340c4050000040000144cc00000000004c144c010c0c130104400000003100f0000c0000000004c0100003400c103000403000c0000d30000cf00041c04700c0044341403400001cc0000000131000d0000000000505c00d4c04cc004000000511053d430040d4030000030c100100000150001030000cc000000d00500ccc07004d0003030300044040c0310c000c0cc410000000400441400000c4c0000cd000001000500001043c30000004c10300030000003000000000000000440f004000c30300c10701c40c0cc000010000cf404c0c3500000003041c00540045040c03004040040cc530003340700000c00c000cc00100000000040030fc30c04000000300001001400f1000d0104043000f4100500001003501433001000031030440401d00010050000cc0000c00cc30c3c0000d50c0030c1300c300c0010f01010c3cf00044040010000000d00000000040033430000413c000000c33000400c0300000c4c4010340400c0103100c000100c0c0040001000040070000f00043d30304c400c0000104000d000cc04404cc000000c00004003000033c0004c5040010004c0040c10004431c00004100c0000c4d50044c0404001000300c15000d0000000500404dc00004300cc00c0013c0010c00c044710044f10d00050000c000000000000031c00cd000000cd00c00c0000040030c00000c3c41040104c005c04100440c0c000004010f0f3000000001030000000400004df500304100010000700000000000000004500cc004c500003030030c000733014114000c43c010000000010f40cc004000001c01110000c00c0003c00c001000000131300000c000700030007300330f3000070014003c540000400c04000031c003c05100d0004c0000000000000f040fc0d10c00000c0c30004030001003c3000040003c04010000000d4001030c0d0400000001034c0000dc4300c10100400c0113c010304103040403000005000000530d00cf00c40c030004030c0003fc07401003c4000c40c0007000300103130cf303f10c010c0100c0703000000000c440011300000c441003c0000cc0034cc0c00c004c0000c1c030040c000c0000050000c10d0401c00cc0000c130;
rom_uints[267] = 8192'h40000000033000000c0f0000c3040000c011c0070000001000c4c00030000330000000000cc1c010001000000000c04000503000010000c0040000010000000ccc40300000070003003100040000cc0040001000c100410000400f000000000000000000040003300004000004c0c3004f00cc4000000000401014003040000cc0440030000040000000c004441001000110000000dc1000c000c714c1040100010003053d00400000ccc1400001030030c00040f100400000c100500c0030c040000440500000000c0300340000004000000500004003cc0040400000000c4000004000000000c00cc104c0c04140001c0004000c00040100000000003c0c00400040c3000000c0010c04040c0107cf00030070f00c0000000744c00c000043c000000070030c04c00340000000005000c000100000000c000c400010030000000cc00c0000040c00c000033c040c03000031c04034cc1cf30c0400cc0005000c000040004030c14c0040070400010040c00000c03c000300441000000c0c40010500cc00005000000070004001100400000004000cc0d30040704100000700004000f0f0c000000100c001d400c00f01000c0000004c0c04000000c001f0c0c4040000400004400000c00c100000c0000c040033c100043000044303c1401034003030c00000c400001430030050c1cc40003c0400010000010cc33400010c7310c10000010cf0c400001c00c0d00040010000000700001c0000033cf00100c00500000000000c000000004000430000000100dcc1c0004000c000cdc00c00c0000040000000007c300410000c0401cc000000000000010000000040340000000004000440c003000000040f044040400300c0003400c0c0010040400400c00044010004c03300c004c00f11004004c0370000040004400100443c0004dc0000000000000100c000c30004054c0100000000004cc400470300304000103040c0f00000000c3000030040c034000140040c000000c4c0c0401400c000c0000c0003000400000cccf000c00000100c404c030401400300000c0100cc00013000c0430000cc00d00001000004000003014000040000c0013000c3000004001000030c4041000500c00f00c0000030c04400010043c000c0300300013c400000d00c4000100f04000000cc00010c000170030400000c4001f00000000000c0004000c0004001cc0000034040000000001000f0010040010000c00340040c30c4040000000d0000300000c04c0004f004c30000001c000c04000000c04400c0c0000004f1004000700c40c04040000003330004400c00000c000000071000000004003c0000f00c000004000c004c10004001030100cc0c034000400c4000010000c00000c00c4000007000000300001000000303000cc4000000000040000;
rom_uints[268] = 8192'h105000000010010300410033d00c00000c300003000c1034015f000c300000103050300000d0000401c0014030000730004004100014443410340c303000f0033000750000110000000000033000d0f1d03010341001f001110070003400010407d000030040400c0000340073f004043004340000d30cc0000000f00c300000407c40c4004c000000000004fc1400c00010000000040000c0000000cc730430c40004001030330000101d10100330000040f0000044000000001030010c3000c5100010000004013010040100010004000f04000f0000040044c1f400c0000140c030301000c000014003f1011104003300000034000000000400003c0000040000000000c00404c00014130030001003403c7c3000400c70000410cc40301c004c00000430000d00d000100031400004000300d000c0044000000000f4000400330cc0c01040100030000041c01400003011d00001f01070471000d0005000033000703030c04c4000c100400010300c3c1000400f04140003007400000004c0c00d40310c10003130000fc11c0000040c00c4000ff00000400010300000c000c0303000400034305030c05010000044d010d100300c0000f400fc000030340010c030040000f0040510c33000000400000040401c303000040c041c00c0d3000c0010d0003c403033004d30f0004c00000410304001301000000cf0013d10040c3f00304c0414d7100000050c00000440440030100030000cd010000040c041c40007300c05c000003001f0f00000114c0000011330c03c11303f30043c300300100100040000300140107ccc070014c400040010c004311000343000007000040030c0304100040c300030000c0431304f0001c00000371c00300400d04c00c01000303000c03f4041011400007034003034000c1d003c310100000071c00c00c010300040003030000003f03030053c113000000000000c4c03131040000004d0000000400000007010004003c030d4040000c0343d003070cc300000003004341000103000030010c404400400300004c0000000000c05100010000001c00c00f01c300010000710c0004000c00000000c003000000050000030030030c4c0003000100004300000000c0000100004000037300000f05040100030c440d500300003300c30013034040401040030c00cf0001c10100c3030000000740010007070c1d0c3c040000c1300300000000000101004104700c000dc0100f054003cc004000400c0d03004dc0d000000cc00c000c474c00011030000f07000000400003c0300000000030413101013c00440cc30000430300030300c14440000001000401c0071100400c400005014cc40004010000004000c10c4404c010300c40000300000c0000010303030013430003000311004103c03c000000000300;
rom_uints[269] = 8192'hd140c3000140d4c0c000c0c00041005c33404043404011030100cf33c3d0f1000030c041cc03000044030040c01000000000c0010330c04c0000000000c0303001403031000013310000c0c0030001c0f0c74f1001d04130c3c0d00000000303000430070001000033d001c0c0000743c110ccc34c01d0c000c00d400000c001f01000000000000000030000000430c03030000000cc41c0d0f310300dc340010401110000c14300014d40c0400310440040000300030044000340001dc0c0003044c00000000004c0001100c04040004dc00000004030c0015100c74040000c30103300d00010c300430310f00c01c0c00041c3103000031000000000000030c04133c0300c410001707031c030d000c040c1c01330300300310001c004034f0031110011d10c43c14c10001000f003c0c304c03c03c3c000f040c003540040404040000001cc000c004003c400005c00c0d37c0c011000004000c330000104d0d3f0000303c0c0003310000c00003301004011c0c040004304f03001c0030001c04040103f0c00c003004000c0c040000004cc0000040003c00000400000000041400000c30040f00000034041704140030040d3030cf00040c0000303113400c044c000cc431c400000c00000f04030f000001043c00c0003004044004cc000000f0d01003334001300c303c000f0c0c04030c00300c0301000111c4001304000101304f34011000c00c300c30000000c000003cc3000ff31c00340c03c000c4c4c410000000d00100400f00010c000c300100c070070403141033000c10033000c0040c000c34030c13c00534100c051131040014c00000c000140003100d04000c0c00c01d07300c3c0c0000c0011000c40c000503000014000f300c301c3003010c343000430c00000074d00c000035051c0c000000010c010c0cc5140c041300c40c03000c04c013311100033cc00004c0040c00340c0c00c011100000cc70040010003c3f00047000000330000004000c430000070c000010040c3004000c3000c33c0c010500c0400c4000000000134c3000101f03040f04100d00103000cc0410041400740c003c000c0c4410000005050c301000cc0400000004101001130c07103300001c000414040c010d3d1c000d0c0c0010130000030c3300000f0410c3040001100d000cc41c04000004140d0433001c30f10003001030d300000c04c30034c04c430f0c010ccc3000111400140c00040fc400400000340140011c3000000000c100040410101cc000411d04000040000c04100404000c10100c040404040000c00010101c00dc0000cc000d1c0000000d0010000013c000000c4c1300030cf30000400c0000001000300000051000000000cc04003f3d000101c00c00400f30000c00430431011500030d0700031004d000000d0004303;
rom_uints[270] = 8192'h1701410410d000c000100000010014070c101033340dc0031410c3370fc000c00000004c01c000100440434003033c000d4000003503c041000030034d000300040043c3003040d0000f40f0001cd10d0034cc4c30413c00000c03030401000030000130300f00000040400300304003c0c0000400404300101003004c00031c30000000ff00000c00000c000000000001c00c400040000040000043c3030040013000000000f000103000300c0c00300001f30003440001000003070500000001c0c000c000070401c010010030f01010340303700000c3003033013000c413401000000041400000000df0040040101c005100030000000000000d0c10c40340c010c00400c0010004040fc005f1000100400001f4333000f013400c05c0300003c0001c4300f03503001000c01cc411300001053d700040030000c3010000cf03c0c030c41c04c00000707c50c040c00004c40f0c0103730f3c7001c400000c00003f3440334301001000070d30000007001014400070000f73030c00030400300500c50401010000000c30cd030040001c71300c4030cc1033300c00000004c3300000100000000311c30000000400010c01c0400d50070c11000000003cc400003d4c434d030004c00d0cc00cfc430c0344133750d00033c00c03044401100334113f0c03413c0c3000000300011c0c0004f00310100100034d00030430f10c0f0004000531001430c0c00310000f01000c401000100004100cf00731401413400003134130340000400c0c100410100000003304c0000c030f400f10043c0013050010000c040100003fc303570013470434c4c00030c00040c0030c003f00040340000c0430044143c04000000f01000c14c01010330540014c100400f0c040040000034300701d0fc0f0004ff4fcc01000c10100034ccc000013300510100404d033040c001004d3f000400011050f0000c00c35f00000134003301504040d00000000034c300c0033c0003037c0f5004130c3c0c41f004334c3114f10040000c10c0410400040440cc000000001c03030c0100000000033d00040111000100000c00003000070300f000510140d0c0c0c0400c410c03d03000043c40300000300000000030c400310400000300001c0030040c010100101000031c00001c300001500000303c003000000033030003000000c0d0c33401301d0000101000000cc030000070001407100510500d3c4110030ffc1c00400c00c14000c3f04dc043001d000500034030440030003030d0f003000000000050030410000003c5004c030f140010001dc1c00030005c303000005c00000410004d0004003c03004310d0f4c000003301040000cc330300000004c004040300dc35c410301c34000c400c043430d400000033c1c0100c000100010c0d44f00c530400300c;
rom_uints[271] = 8192'h10c00003300d00001dc003c00310c00110330fff000000d003c7c0000001000f010140c0004700000103c10400d311c140d303c0c0c00100040014400c000000054000003500000d0000013140004004d5400051000c00c000004054300413033c10031000cf000000005cf00101c00c010c4f040300007d40c0003000000fc040001000c0001000c30100c0001100c000004453c4c000000404010000d734000313c400100040c0007400004030000000000130c000c0050403400c04010040400000017330c001400040010440c010f00001030040000440044000c1400000000100000000c343c7c130100300000007000000401140000010c00040400000000000c000057000000030000310f1003017c3000c0f00c044040c030000cc00004f1003000700c00300000000000f100043011000004003dc0140cc00431040000010404f73c3004004000004c0c000034c0010c500031000400100d003014003cc034044004f00d05300000000131004d0000f04030100000013d0c000010c04000000c000300000000300c3100301001000401c0003030330031c100d00000000010f100100040c00030400f00400d141404003c00004000400403d300003030101003301100101700001041031000040cf00100040000003004c03403c330004c003c3100400050000000f130000400001014c0000004000040cd500070003c37c000301004000444011010400c4c000403000000040003000c4001000000003c001000040014f0044000000c00000000031010000013000004003c0000000001000000340001c40f001000010c30040fc4304010007010003c0000403000cc5000713100003d00f00000000013004000c40f30d40000353030010c401340c000410000f140000c0404405c445030c43103ccc0300010f000400100140cc4d4d100001400100d30c00d040c0000001c00cc300c00ccc0330000c0031000000000004cc0113c34000f040430f40c3c3100000400400004f0000000000000035c10030004cc0010000000c00000c3700c010430300004001300c0001c003c7014300041044000cc00300000130000010100003c003c00000014d450000f004c40c03c000100043004000000043c70403c010000500000140c0300000040c340030c3001c01001305040c004010d000700070043044c01000030000000000c030010004c3014003c40000d003d100000104000001c1c000400140c0000103400c40000100c00004c5dd40404000000cc013c40000c400400400010010dc0000d001014d0000000100f0004330cc7c000770001000c03000040503c00c00344c1040d0c0300001000d000000000040c000c15001400340000100000530013100004c003400c0033000c003000100000010000070c30314cc000700004;
rom_uints[272] = 8192'h1f0000000c0030c00000400000c40100041000000f03000004400000c300040011005000040000c0c0000c00000c0040005004c000f00000c00c00300030400c0ccc4003001000000000313000301000000c0c1000000c53000030000010000430000f700c00400040000047f000000001440300047340000c3104000030010404f00000000100004c000c0004000ccc04000000001000c40000003000c00000df0f00030030c04030040300cc000010000f00004000cc0400040c701f000001c50c0c0000c4000d1d04300c040004043c0004000000044545000c04300000004c00303330c000300000043d000c0000104443400000004d01000400000040040c4c00000001000c0001050031011003c0300050100400000c0040fc00300340c0c0000071000000100c040c01c00c4c0000f000c00400053001040040f00000000100340c000030c00d30030004000c44c00003000c13ccc5344c1ccc010403f00c04044303100ccf0c4000010030300000300000000c054c3400000c00000f0c1c504c1c43044c0000003c400100f004000c0000040000c7c000000004cc015c0400103000040c40130400c03cc04304c10031131000400c000010c40000010003c000000c400c0c0400c40000c041c00c10110c340c00c03d40c30c00311000cc310000c0040301c03000310c104c0c001c000300040c0040443c040040c30000403c0f04c030003c07140c003404f7c44c0c01cc00000400000c040c00000c00000c44401000000500410cf0030000007404030400000400c0000001c000030504011f0000000c000000dc0c04003d00000030003400150001c4c00344003340100040003c000c40f034c11c0f100000fc003001000300c700300000400000003100c000c00c010404040001400010c10530700000004000000400010000cc004c040c000105070400054f400004c000c4040040c0f40c0400434000044c000c04c0000c00000000c0000000000c1c0c0300000500030000c00001410400004004c0c0c44c00cc4c1030cc00c00c00500c4000400043001c00040430007404000010440000100000cc000040101400370000010100000c00000000f1003c000107f0cc00c04010000000001c0000f0ccc0404004300130c011040000c004dc010310000c00400004300000001c0c40400c000000c410300030000400000000c0c00c0010cc00000400004001007005000104000c00cc40000404001c0001c04000400010000000000304014c000c0105000004c4004005c400f01000000400c1400c00d030000c0030c100c44000030001000c0400c1403f000d3704000000c10c304300c0030000005003000000033400004400040040c004c100030fc00100404c000010051f400c40043504350104000c000000000c0c01000c3000;
rom_uints[273] = 8192'h400400004400073300000c0f07001004000003d40301410c00050c00030c0300000d010000170303350000050f03340d03000305440c0000100100000d000d000c011f0f00000040000003050d00c403040f0000010c33010303010300340c4303d1330300000f33030c1c000c3c0f033003000703030c1c000c0300011f0c0c000c0c01000d0010010001004400043c41050000000c0010110c00010d00001c0c400004000005000300000004010004030304030010000301000007730d003004040300000010000001000110103c0c330000003044030c30000704003c300000000000343004000000010d070f0c0d410c043330000001030000000003000c01044f030c0f0005c300011300010304000000000f00040d1c0c0d010003001000030c00000047040c400c003004cd03000403043301cc00000003030f04000c01000100010044040c0d000c0404010003010007031f400700010101100c000c0c000500010004000f0011000c33040f01000d04010c430c01730000000000003707c007011103310c0000400000c30c110100010000030c01013c0c04001100000f000c0330330d0c040000000405010310043d0400000f03000c3c0f4101000503000c00000100010503000300000105010001070c030401070400000041c01c0104f0004f330304030100430f030c03030114c7040400000434000400030301017303000000040030000f044004000500030000030001030001d503000700040410030f0c1001000100010000000f34000f03040c0c03030c00000d000c000c000c0c030000010f040c000013000100301d03010405000d04070100000d010d0104000f0000030507000c0100030c0303001000010300000c030011000d0d000f1c030c05030c0f0c010c4304000c3c000103cc01470300134c00033f3013000033030110100003310cc4000003030150000c00300300000003030c00000003040d000c0040003003000400100305001001010033000c3300100c03030100000000053100000703003c000f04070003000c1d033c00030004040400030c00040c030010030401010411c0000c0c040004034103100d0301000d000d04000f010100003000000401030c03000403350000000110c001000f04100d01030000c110010300040500004c000400010c040c000d0001010c0503000c00000000040007070f000c0001000005100d000140034000000005c10300000001034000000d00000100041400030c000c00004c0c0300010f030c310300000301400c03000001040c00000d140000010d000c000000003c0300050403000c00000000101c0c0c300700000c01000004050001000000050c000c0304040001401000011130040c00000334130c11003300100000000100000c0004300000010001010c0100;
rom_uints[274] = 8192'h40000030301c000c3100c33d003001000cc410703c30040f0c700004033c0030301cc00310000110100000010f404430031413503400c033040000100103000007000100000c010000040c0000030c4c000c15c010030f0010001004c0440730750d14f131fd000c37000130100400030341000c7f0f0000c0000000cc07040441100533300c00140000300001030000000300000073000000330401000c000000301004003430030100014300070014040100003cc5000d004017000300000001040104040000350c110000000c003000cdc01410010c3000005400500301103004010010001001d003c41c3130003f0300030100010030000010000004d430300c0f1014c101000c0f0007000103003507103400010c41000707010010030c1c0000330073030c100c015c10c050043000003011c00401050000370030cc300300300d03f00000003df5300000043f34013c0441003030311c00000740cc13040000033100003104033c300100031003130fc00030003470003d3030040c44050003000c30050410000400040411030d050c0000100000c000c5003700000500030f03300d000030030c001030003c1034044010030030105000100304033c000f103713cc0030400300000001040104037f100011d30011040000010301103c073001fd10d3040030001010000010007104400300000f100300010c333440030310301004103c13011310140c00103d043d0400031000000001030f310004110f30473003001001001d00000000100d1000000030340341300001040011340001f4100c003104000000004c0c0004010000013c0030474d040000440300440004010410c10c01030300303001001000000f001004031007c0013d00000000cc04030000300c300c3501050d0300105007100f0300100c700003400413130c3700000000000000043f010c350040040c01000000000410030f3040300c0f34000f0030073c03007330000c00370001033c100100100003134c0cc313000c00000103030040000030d4f0300c00040005001f00030001013c4d0d14030c00000013410000014d4001401000300410100001350c000d0303303404401403000050000100110000cdc010030f0f340000551000000000050c000734043011030d040c30000300031041300144f0110304010000000c13130300540030331430040500040000000130003103030303000c0710000c0000000f40000334100001000413000003c03cc0000307070d3c11414c0c040331003f000010040d0301000013410c000100300034030c300000000c00000300000010404100001410003000f15033003c30400100c73011c40000001130100c000f07570c04004c0000040c300c04000040c43401c50dc311100414033c3c00300411000034000530f40;
rom_uints[275] = 8192'h4703000500030fc010cc00c0d003f4c3340000c10c0f730003d4000c300340c0440ccc03010004000cc10001000c7030c3f1015f04340cc400000000cc000c0040014030501004400004000cf00c100cc000000334444030044040c001000001001c41c00000c0ccc3004c0cf000c0f00000c014113030cc0030004cd0d00400000430040cf4040000c03000c010c00c0400010000004400000c4000001010040c30440d000001d010740c0044c400504cdc3400000341153c00cc4c03c00030c410010c000cd1440450400f0440303030d014004000340f400c01c007330c000c10030c000003000c000c00004c0400f4404cf303004030000000c00700000cf00030dd4c741cc01000004053040040434c41c0014c014c1cf0010f00d33d00c3370004430000300c30043000c03cc000000c0c0403000d000c3000f440150340314510c010400300000540134074000f07040300003000050540400400000c430c0400303f050011c11330304001003003c003cc00003400c01d0c4000404c30c73403c300040c000000c01000003000c0404000010004030c0001cc040000007010000310c400000c000044000000d0000345103474000000000cc0400c50c0130030104100000013000c000013c05c0000000ccc0c4000301470000000050c0005015c30c440c03000c00470000000004c1cc0741000d03c0100ccc34f3000000000030140cc04104cc5c005c000d044cf440007043000035400d13ff0100140400d40c5303001c000000101013c0f00004004f515c00c44700c0000dc003014400430c000000000007000d4c44000d10c0000404040004013041cc440fcf440150400470f01f0100000000100cc040000c4004103004501c0cc0c10003000500000300c0c10c0f043cf0004c40f04c71000070333000074c00c00053500c04fc030101400c030300f00000010100d030404000f0004400f0350404c000c401001003000340000400040c7040000000c30003c03007f1c003150000000000000f000f400001044d000001c001c00000133f030000c40c0100004410d0007700043305400434c40100c1c30f0405000c04004d000000c4c34740cd4050140d030005000430310c00040d100050400003cdc70c0000005105c0470c00c0cc004c4000000c07300043501040000c03c3c004040030007c00104000f3000f0400100c04045400011300000000504c000000000c100c330500c0c010374433440c0c000c0000100c00140004004300c401fc4730cc401000130310c4000400075004c01000001000000004031133000000c30440300310c4400401004000c000003ccc1c00c0001d00043d0133000401040c40c00003001f0000cc0000040c0c0c00c00c04310413403037cd00047000d70c0c000c3110347f0c0043400d0003;
rom_uints[276] = 8192'hd0c03000040000d003000c0133331000030307000c0000001c4331100030004030f100001004000cc00000004c0c00c00003000c07003400400040004300310fc000000000000411740000003000c00c0c0110000000451f0001f400c05c3303000000cc001c00330f000c101c044070010444c000c101f4010c0d0003f33000040331f0040304000c00010c4354033d00c034c0c41040430c300c3103000d000c0401cc300c0000100000540400d301000cf000c00010354000030404300330400305c43c04003703c0031003040c400000c0c7300304000010c031f0f00000ff0c0101007400100cc30500043033c713000000c000310cc0000000000010000400c00c000000000511010330501d0001530000c17400000701000010f40000300003d43c130c0400000100001430c030000000010c30c0000101c1014100040c4f0c00130031cc4000004140040f0c03013003310c1054f000050101447730370310303d003040070000700034030c0c34101c350cd0100000f4cf0033040050010f0300140000303c0330c0013000c000d5030100100040143c33f03030003f003c000401100c101c305403c4c000010535c00404004010003000017003117cc0114300304030000000000400304f000030f000c00d0030311001040010403401510300015004000c0303c400044c04000000d301000100c00007003003c0044404c000d0031c3003f040003d0440ff3000000c00f707d00c04f735103c00c531f004400110110000004403033c000030000c3440001c1c00301004130000000040c500f30c34543ff0c00040010004000310003c450400304340000403001c00034153004000000c300c50330400100cc14010c01c01c0440310043034105000040103330000041c0000140c0cc004d0c3f300013000110041003040040004004310300030f501000c35004c103d1d1304d01c030000040000000000cf0100000c30c30040000003c30c0c00731c30c0013c1300030d130c0cd0f000030403f107000d1c0050000100040c04c30010300000000030033f400400c300df44f0100030c4000004030f0000f0d3000473300ccf000c1000001001f1000c3004000000000c00000430d0f04c100403040300300c00000400441c0010370f540313005000000000304c0340c010130c0c03d0000000cc00000f700001c4004c15001c0000001000f4041300d0c433000fc4414405040400004330440440310c0c13040131010043d050013100003000c0000014000303c1000c00503000040130001000c034000070000000c003c3045000000f0000000000330000c1c41cc03300101c3003041000004300000000300000f4cfc5c033c0f0f100001c00cc0d003003c0000003004c31000c00150000010c34cf105c30000c0c0c1c70;
rom_uints[277] = 8192'hc0700c00ccc400700330c0000300011c3000000040110430007c00004c153c0443c047401007000030c4001000100c004410033304703010c00300004d0031000c001c1c0000c033d00000c030004300c044c1003000300011705f07031314c500401504000104041400005004100000000000043c01007c0040030330010310fc000404c100c0000010004011007030003c100000f0000c03c010004031005000100100101c0500001c00c000c0033d00031403000c00c1c0cc00000110000f003344c000040300433c00004400c03c000030300300001401c30013000c0000140700cc03103000001040000400c0410d030350c0c000010001010040030000f03004000f310fc0470c30430070000000030003101010003110000c0103004f005c0000001315311c35000040c0c3554001d0c30100000004400000000c4000c400c03000c0f100530430041301033c00d005f3404cd404c303033010100300000c540035140040c404030000c3c3504000104300000003c0150c000040d4040000d003041000000f01400004043000030005030000100030c0301000c0c000fc14c010070300330000c04037303504c03000470400c00c100100173001300301040c0303001030000c0400330000140300004c4000404000c310000003f00301c0003000c10c3000303000f13040cc1c0000c304004300000c000100c00305c0000530c03400001030030103010005040434000000c10004f07043f00c01004c001010413130500100300c000000040000000000140000410000000300400300c0f5000000c40000c05c500cf0400f0003c00030140100500300100000041c00000400431030010000115014301000000300401010c3c00333f00044004400d04c0040400000c14c00300001c400304100c0000003c33000c40000770c111000000c43000000c0000010431030107c0c40c3d0f00000f000401f70004c0c4f0c00c030000011434010000300300000c00410015000c3c047001cc7d30c4c04400010c01453007000ff0033300000050004104000d010000000c000350500304000300d004c00050404f0100c004000001017053000f00000040f0003003010003d00c0040341f010000000000310000004004d400c0c00130c03d1c04040c0730030001100000000110c41000070311310043d040d0d301031c100003003c03c040000101000731000c0c35100400100040300033010100050000f0c4441003c005343030000004f00c03c000c010010040c001470714000030c040510504070000311400004030040000c0303000140401f4c4c0000000031000030413000c000c000000000c4c000cc00000f004000c4310000c030510300c004301404c404c000034c13300d3d3314033001000000000000c0700700004cc4c053000c31;
rom_uints[278] = 8192'hc0000000c00000000c000d404000c000c000cc000000033000fcc00003f500040000c400000100c0400404000000c0000003c0300400000300000004430000c000000014400100c00000003c3000000000440000400c01043143c0030001300400000400d340004cd40fcc001c0000004010004c0000100000300100401c0c0000f000000000000000000000000000cc00000410000010000000040030cc40400004400c0000c04c000000000404c0d00c0000000000c00000c30030c000004000fc0010030000050040000c00004050c0004040000004c0000c0400f10000000c010030001430004010400040cc00c0010014400000000000000000c00000000000c000c00c300c5304ccc1f43000c0c00410000030c0004c00030d0000000cc040010000c000c0005000c071c04004000c000000c40000040c01c000400000c040c031c007c10000c000f00d000011000c7050cc0030000330f4c00010ccc0000000c0f0d44c000003c114d0c000000000040c4410f0030001c000000000c0000140c100c00000400000c0c01000040c000000500004003f01000000000100c01400c0000f007c00001000007030000004000030400000340000c000054170304c04001000041040303c00000040040ccc0000c03000000000c0003c4400000100c00000000003c00f101304c000000000c0c000c00000c0f0004000000c0030000400c004c00004400040c00100d00cc00000c01004c00000c50000c0d000400400c010000c04000000000c00030044300300000c004000500400300030031c000400c4400000000000000040000000000c000000000000c00000000000040300000000c0cd00000c0054c03000000031d05000fc1007400c000000000400c00000301000000000104ff00400400043000000000ccc740000004400040004c000000c0310c0043000c00030100010c30c4c00004010f300000400030000000001105c000004000c00c0300cc00000000003000040000c3000d0f000c400f000004000000000010030401c4c40000c000000c103c401004c300c010310004000c04f040000c0c0000000000000f100000000005000c00000001000005000c0f1000000400011004040f0c000000400040330000004000c0000c0c40003000000000c000000c00000340cc030000c410000503400040000000001000000000000c4000040c0000cf040000c0400000040fc30000104c40030040300300100004000000000004400000007000030c05c04c0000cc00014c0000140001400101000f000004003040c10c000103004c5000004c01040000c0000cc0000100c300c4c04c01c04f00300c04c0010004100404000004000110c00000107000c00000700c00300003c00050c0000000c40cd0000003040100000400001000000000000;
rom_uints[279] = 8192'hc0c0000000c10000c100c040000000000300c3400c0c000000001000d00000000001401001500000034001407000c001030001400000c3070c00000150400001c030000000000000000000dc0000fc00000003004000400400404c40000c400337c1004000c00040ccdc000c00010000c0000000c000430001000c0003c0400173c000000cc00110010000000004030000004100001000400000000000c001400c01d000000030000343000043000000c00000000410000010400c3f30030140010040000001000000300000000000000000030003010000cc3000410310000040000040700040000000000300d0070300f301401000000000c00000030000c0030000434000c0c000040000011000430030400003000000004000c0000004c043330003000040c0000401c040000c000001000000040000010000010cc00f0c3000c0400000c00040c00011400070c1c001c00003400000c00c4053000000400043400001500000cc050003000333000c0753000003c00341c04c013003000004010010004050000000000f0000f0400003000003034000000000c00000000004700000010000000000400000000000c00140c0004000d30000000001007000d0c0001110404c100040000000000000304000040041004300c00000000000c300000400000004001011000000110103000000000400100010000000010000c130004000c0003f010001c00000c05100c0c0000010034000000000040401400400d00000d0100000000043004343400000000000000000c000030000c000f04000c40c0013003000001000010001000400003000000303003f0110000000c100cc30040343000000300010c3c00000c0d4000c000000c1030700400000001000000041510000000000133303c1c003c0400000000300c1400010000000301040c0000400030030000cf03340300000c3000000040130d00300c03000000000000003c1000001104340000000c4c40000c043301011400030c000d0c00000c140000000003010000000000000c030000000307f00400000014000740001dc0004500300c00700000000301040000000c000f04000c000d000c000c00030c01c0070000030c004000000cc00000340000000434010040000033000010000004000c000c000000cf00000330101c30000017c03000000c0c3007000000003c010007101447c034000310000130040040003000000c0000000400300000000030000300300c100010044000103300100c00000000c00000000010000c00000c000003000030400403010000000004000c0000030f100100303000013c000c000d0000000030013000401000030c004c000c0c000c00000100040415400000010000000100041d3c01003000100000000100000000c0000c0000000c001130010000;
rom_uints[280] = 8192'h1300070103f30105c10010c11035300c331c000130300300001134000370030300040135013d00000000003111003030031c10100041c701c0000033330043403003014010040000010030373c1013410040003001030c000000d140040c45c00403c10d034001000030040031c01140000300044030101000030330001113305003400030c30001004000003000c511d01f00c1000c300100000c3343041300000000100f3000031040013043f0c00c000030000000cc003043000c00011000330001c00100c11f70400044c03301c00000000300030c40000c0c30151000004000001001c00010003300300000331300c10c0f0d0300101000000100001000303300000310ccd400305004003000401334c01030303000000101c0313300f14000cc00003000700000000340000040110440c30010010000103c0c3f0f0000c333030003300000730103000004c0c3430100c1000f00f005303f000010030110c300300730000340130100c0341043033030c00000c33000703330000000c30500000000000111013000004f03443c100000001000030000d10130330300004140f000d13010c0300c1405000300000000140314130500c303031000030113130c0cc0c0000d0400431140c10004c0043100001040100c00c1034013310c110040045300c10300005f05000310001140004310d0010f10030000000730007303103300ff40c0034003400000000cc307c3d003011030004100030f3f40010000000d00030400400c00c30135300000030000004001013014003001430003143700c0c04000010000010050300040030000c000c01000003004343303003330c4c0331030010003030030300c00050000f010cc00030030000301000fd0130300f104000300c01300c1f300c010100003001000003f0000000f1c0013010040301333100303c00004c001433003c1007300100330030f0000c00130fc00013311000300000004003340c00c00000300731570010043c103003c10d0307014110c0000030100444c00f010014f47000000070173310100004004c00000100000100010001c001003000cc700000d130c03331c004001030000c30c0003300000510f0003f01000300401100f070001c4000000314103003000000011c100001000010c0f0004fc0c003043c3c00443007000130000010c00403300000cc01c00000054000c0f01010c100000f000c000000400000300c0d3003000000043000011000c0000000043d000440000000300c000c30703000300001040000f000000c0000000104300c3100000101c001f030010000fc000340c0400030010d00400500047730c1333d04c10000300300000c001000040030073003000000403400013031c00040003310010c100400c01000000000f00010000c0030347530c3401;
rom_uints[281] = 8192'h40003000010331750100c03c4d010cc40f700c0000c14c4000030301040340c1400c3000030c0c01500103d1c0004443f00f300301030c01cc01d0403100410004c00013c73100570100040d4100444440004cc51404041004c3f00400c0130300410000cc44c10d010cc0410003433040000c00000000c4000000c1c100100f404370005000c0c410000003000001400050000000c100c0c3f00f030030cd033c0d04100003001c00430140000c00c0c001030000030101000c3cd4c04000c10c4303cc4000c1035070c000001070050044ff4cc01050430434410d4c7dc0cc040030304c04c300000c00c31544400c00010004c0400010d3d0100c4300041000100301c005040c03014444304d0c4503f00001c30d3003c073005f10c10044c00700000043000003340c0044c104300c1000c00440cd00000300c074131404503ddccf300fc0004000004cf007dd433c333c00040310c0000dc4030c404000040014010700700044110ccc1f000c000300334300c04d570c4034c045344000500cc100d043001301f04000340003100000431010004c007033c474030c00000c4c11c0000304010310cc0c0030c00ccc0400300c70d44000c74011c0043500cc5144010003c01000000300dc00400c01441c03040033430305c000000c401d4c1c014d40c0f10300c0400dc4010374330040c0dd0040c0705030000001010d000004c00cc00c00110003010c37dc1000c3cc53c000300000300c4c0c404000040f001003300053100004443400c1c7003700c0001c44000fc0cd30400000cc01000000403000000c1f000001cf0040c0011c00c040000c001531004700004d001000001c1000d500d07f0340004700c5c0d0000054103140100000cfc00f44000140010000000104d043003d1d0000c1004300430401400013c7c4d00c4c010010cc044117300040c000100c0d0c0fc0010dc0c030314c4100310c001fc13c400c00050c00330373c1734001070000300f130000700d140d0003d4004000100000000140404353103c0451d04c011003304c440c3cc3003c0cc7004710cf414330000753400433040013f03300100d07014000000cc1cd0000000cf0044300fc0500000c00000000f10330c1c00000000330c003cc00400400314c3000340540044c0000c040c0007401041400d103003c140cc44304c11003c1c0d00c0010000c00004740000003010000400c40c40c44030010014300007300000003c043450043530001000000000001d00704047c7301000c0040000f30c1c005410004100c430303001010433c4014c0000503c01700014100004401011f00c400034301c0011c03004fd37044c10c34440010c000d040040c440340c0c1cfcc0000c00000d0000c1c0000c04c40f11d01300000037000004340001dc00c4340ff0003;
rom_uints[282] = 8192'hc000f0041500100400f000040c5cc0dc1030c050004301c000c100705c7333000ccccf01005030c005400340fc301c100130000331dc0c4030000c10000c00000400010d0000040300041007400410300040000050c000000c01d010044034f0431c0040c00130c00d00103cd7d1304000dc0c030001c0105c4404105004040000c110000030070300100010400010000030333000034c3300d030001040c00c000030c401000430c00001004030c440cc0030c000000440000003134d0000030c000030301030405c0c004034001010c0c0010014c03010700003410000c0301000040300003040104017017d0031000c7043100d000050c1d0c300c0000c400044000441d4c000145001c030500c13c3c43001010c3130cc3011331c00000000100000000007103c0050c313001c000000040010001000400c0000d410000cc00045c00013040c1c3030401000c00df1303cccc101043000300130c0cd003000c00000cc3c0000d40440c0c400c040000c1430330dc0500f0404300303000003100c01c0c00c00d040100c10001000300c100030000c30fc304c0050c0300040104171c000000001000110300400004c00f440003103d00450430003100041300050d0004700513c0110000000c30070310c00041000001400504d400dc410c000c110c00403d5c103c00001d40d00000330f00130010cc7003040c00d04d0010004000cc0000050c1c300c130704001340001403c00101dc01f00cc01c300004000c404f100c004f0101c134040034500f00c1140000170c4c0c10000070010c101001c0040004707c0f0c31c000304400c0040f00100010f0100c0300c0000410005cc4113c0f0c04040f040000040ccff013041d010040c10141dc1c0c00040041c10c40001c0c3004410171d34104c10001d040d0001410050c0c034c00c051000313c00403300c300007000000040c04d3300d4534000f1d1f0c00cc0c004001000004010000000010110c5000000003c0343d4c0cd4004041010044030001000c0401010003010440003f0000c0d131040100000100104cc01303cc430c4c01100c34d30400d40d00c01004c000300001c1ddc000010000400400004315400030d000000304070c0304300700ccc7001100d10d0500101c0c00304000010003cfc70d0c0c0c0000004110100100145000110000100100001c0c00007104004f000300000f040f00c40c3c500c0f0300410000c00400000000c1050c0c4100344c00c0003d00001040005300c3c0040040033401000000003503400d001004104c004c13c000000c0730005000114401c10010010010c000c000d00000413c434c00330000007000010400140000040000400434001d000c0c0c044701d040000000100000c01004c101110030c10c01000c141705400315001040c1;
rom_uints[283] = 8192'h4c00000007104000040000300040100500040000340c0c000010c0000003c00000300000005001c003300070300000cc3000000c00111004410000000c010000000011c10000003000004003f0100040000f34133000400000c010cc00101100000040000000fc0000001000000c0c340000000c041000c01010000000000404001040003000000000000000030c0303000100000000100400304010d0010010153330d00010c1d0040000300c07300100c0f000001000000300004030001000000300030010500013010c10cc100101100010c000d033001c0030300005000c00cc0010f0001000005000cc104100d300400000000000000013100010000010130000000c000000c13000000000000100130004d0100030003c00040000003400003000001000430df110000000000c040140000000000010303110300130000c005003003f01000033041c310000c1000000003010c00003030030000004003c000003000000c010001010c003000000cd00001c1100000043001c10000c0000043040004000401c0010031000100000001000010000001000000c5011c0c010010c0c000000000000001130c00010400000c0073000531000d0000100004010004c0c030070100040cc001000000c0040c0c010000000100000400000103c00004000c1c0005000000000cdcc00110000d000000040100000c00010300000c000c0f31010000110c07030300d10dc001d00c00014300004cc4370004000013440031c000d10c0000011000000000000f00000400000041001003310000c0004000000431ccc00030010c00010101000100110000010300c1000100003071cc00300043001100cc004441cc0174000c01001c10c030140340001101300001030333340c010300010001c3100000c000c0110d000000000000000010000035010100c000000000040140007000000001c10440000010c0c01004000001000004405000100007400030000341000003000000c010471cdc03000c0000044000310000000134010000030004300400000441011c0400100003003c130cf0010004000070030140003c000000000fc1040ccc000001100100300500c1400300010f000000c330000c0000401001000000000030344001330100057100d30003000d00000030c0000c1000cd30300c0cc010000143400400000110410003010000130430c01040000dc00000c00f0000400141c0300000c300051010000000000001000c00c00100c300000001000500c00031c40c00000101000c0011000010010d03300104000410010140000030c0000000000307000d00010c00c000000d000003013c030c0001030003d030031000001f010000010003c1c4403101000000300000000000310000431000010c01010fc003000dc0010101430105000000030;
rom_uints[284] = 8192'h4001330314c001310001c030c00000cc0000100030c0000c0001c300c330310330c10d33d000000107040cc1500c0303c101c000c0403c033000f0034d0003100f040fcc0001000044000cc0000000c303f00c4107404301014300c7040c070400c00031d00000130000030c0c1001410003034110030340000c04c310000400000100010031000000c003000300400400310000000134f1400010417000031f3c37cc00014fd00000430d01400000004c4000010000010000100003300000303000c000c0003000c03d40340000fc0f0001001000140c00000700f0f0001c13003d0000005000003c000007001f7d10050100031c00010050100c000000000c0c010c070017cc04130c74100cd00430000707300c34300000c30d004f010c000c43c000044000100050100004004fc3030350000c03100013c0003c7000cf000440010101114d00400c341031400300404c0010340300f7030301400400400cc0000c00040003010307c003000030000440700131030400051073c00041c00d1304074d130300014c0000c03f1003004d000000000c1070053c0030303c00004dd000100f30c70d000c43030504001004143414f4c31740100c0004400c30c0c100000304000c030033c0013300000040000100310000c00003000cf70303030400000d0100014c0440c00c0000003c3c4000c0c7000c0c304103000403035c0700d004010000c700010f04c41500d4000cc1000c00100fdc43c100f03c130130001c0300440c0300c4710000c00110050000c01110010014000000340031c411c004000c0c040000003d0c317c0c4c410100003001001003400000c0100000070c0d0011030c013400ccc000010300c031300040044300003153000400004000c10100c000c0c30c00400400404d00030500430c300000000f0100530d01134c0300003340040107c70c1f00c71c10c300c000000c0f00107d1000030000004300140300001c3171f30100030c3d0500c0c4100c1f0404d04000c33400001000000c3013cc030d00f033010c10141000300343cc1000300c0407010c134000013004410dc1000040000300000c030c040400140c0000c00c03003300c3c01f351c010004c01c31003d0130040100c500003400403101000c110300cc0000030000cd00030034c3c000c1c1000710070f300000005000050300000000434000411004011f0000400130004400000110100400c400d030c30c5f00004040113100000c0cf0301c0001010004133c101304100114010c040010000304df0c00000130301000501734000000003103000100c30c0d4c00c700000f10000044300001c07704f00430cd0cc304d0003c1000300010000cc010330c4c0000d3003c0400000330c000033c01450000000c0c0340000003030050030001c30c110c0000;
rom_uints[285] = 8192'h3440000040304010000000000c1114c110000035000c300c0330cc5d3000004c1f101df03070000400d000300c1c00101410004004fc0004004700001040c00c000c0070000000307000000c000010300004000040003003330c0040001c033034001c0000000400100c00000c000c0030f00000000000c04103001110000c0f00003000010000700040100000404030f53030300000333400103f000c401004000010033d1c00c0340010011410015000040000001010000010003004300c10003004c01000003c300000400030c00c00030c100040000030301000131c01d00000003000001000400004303c30310030040c00103000003000c00000000050003000130010c404c044300f0c00040000000000071000000c001003401c0010000010000c0c3c300400407c100c1c100030400030300400103c0300000030101c0040100304300010000000000004d00c0c44c000cc0010f11004f4c0c000010c10000c301001000400001000300000c0353330003c4030c000f070000c304c1003141c3100000c000c0c4410300c00d0000c0400003300100000400400c401031000000c0000100000443000100003540510530030003c0c005010000cd1400c0c50000c0400000f30303030013010300001c0c00130100f0000000cc4c0f4000c30c410001ccc0000c01010c03000cc30c500000c00000400000310000000500c4c1011500400041c401034d0f010031400010004301034c00400000cc400d0001c0c40c01c0004c000f0000330334f0c000000fc001000300003000f700033140c1000000030000c040040700c0400001f00100c0c0000700030703000300010300030110c10030030c000030000001000c000340c50cc44100330c01000c3500300000030c03031004f1010010c7000000000003c000c10304000000cc000003000110500503003403c4010000030471000000070340000030000cc0000000030100000000c000c04000000003c30dc05c00000c000000014d0f014000000005401000c3000301300300c30000f100000f03010000000001c03300041001017003050c404303001000011100003000410103001c0000c00304004000001301c0c0000000000000004041030100000c00050c30000001041000404000411f00004000c1000c0101004001400140c04c054110400000c0f105000040c00030000300000100110c000040000000400100c0010003031c000300000000004000010c00c100000071400300c3c0000001f0c0c40000010000004740001c0001000fc301d000000000c300000404050c0004c30003030010001cc00000005c0300000c414340c00007014000040107070c41000003030000000c07410000040400104000c30000000133000003011d0003c003000d5f40010d00000300000130;
rom_uints[286] = 8192'hd0c007001440030100c04c000303000001030040cf41030000000304010c030003cdd47470110000c011004703000cc14114000d03040000000c00013040001000000300000c00004000010110000010000400700007000001c03cc30001d0003140000c04000003d40400033000030000f003000000070301c100c00000c000c1030310300c0000000301000100000d103001000004004340000c00c000010003000f00004c0370c0c00000410c00000000000400000d300144000cc0cc00040003030000003000c341001340413030c000341004c0000000c004000003000030130000430000004000000c10d1430103000f034110000100050000410000c1c30c504040000000c10700cd0130004001300010000000c04f1003013005000000004000c740c300014c000cc4100d1c000003013001040000003001340103cc00004040000140000000000100410000004c033000c010c0070000040101010300040000c3040c00000040040000005000000d10300050c10400740d000003c10c40040cd4050f3100330400000004c34000100001000344c00f04003400cc003003c03c00070000430300010000000cc1c000137100c0030d40c0c1040103047c50010d0044030433440100300031c1400c4003014043cfc0010104000c004140cf000000c00000047c034703010400030001c10cc0000c11c00300c00131000000c00000c01000003041c0c3c033c011010400000000000c0041303435c340304c00000733000040c331040400000000c00000c0c00f0000300003000000030400000c00000030017d010004030144040100003000cc0000030740000040333100000300cf0105003133000001100001044000100cc0040141cf0110c34144c00103c1c00000030000001103c14dc00740c3004010030400543000cd00c310113044d0cf00c00000cfc044c003000d04500303000300310004d3000733c00307000c30030043d0040004c00401050c05d0100d10000c0001000000000d010003000000c0000404c10401cc500403c301c300c0c0dc000000040370c00c4303c00011003c400c433c103031c30f000c0cc1544034000400010d30c34400301000c100400c01000000010030c0400301000c10010034c001440d0100000000010c100000cf000000100001c0fc00c000c411400003c000c1c4410040000ccfc043c003030f00000010d10c400000400040d30c00043000c1c013000100c10040f000c3030400cd040c0400c100001c4154100d44040c00001304c10040033000c14040cf4100c00000430440f103010300f107cc0d000101000700004530c100100005000011043107040040040d01000400000100c000010000000130110cc1010400400300040f0000c343000001053f0000004430c001c040004400000000;
rom_uints[287] = 8192'h140c100074040000cc00300010000013c0301004c000d00400334000d4cc0c10004000ff70740000c444c00105fc003cf07c340410c33034313000004f000400000400004110000410000c10c300000400333c3c003fc00000010c3444033011003cc0c03400c0c4100cc030f00c30130440fc003010f407000c74c04045030cc0000400040c003100000000130000300c007000000000043f00300c3400540404030000000c00040400001000000d14000000000000340004040001000c00004c40004000003004300000c0c03cc0c010003000000000000004003043d0003c3c7004000c740004030c10d30010cc041003f0d000300035003430040c000045137c0004300504503c0034000003030c30540c030c00d00044d03400c07cf03c003004000000100c0c100300300030103040000d1040300c0000c4f0cc140c003403000000004000f0c07c04d000c03c100c1c440005710d400f3c040c30403c000c3c0004000c0c040400d000044c33000c0440403004003cc4001000007c41100300070c0004403100003c7000003cf000000005001004340000001710c0047c000104343c50cc0000c000541314004c414000403000100f3500000030030040000000c0001304c00c0030000c0cdc443040000400503000700034d0000401051c10003001001054f050f044043030003c3000500004044433000000030030103010037c144000304000000014000ccc0c3d0033000004040434001000144c0c0003000110000304004100f5304ff04c003400c0f000004c03c0007404005404445044030000000c403c3010c104000c0001c03c00f404c04c004000c03000000040013030340010000403310c000c00f000c0103030000c0c000000300000000030c0d43c0014000d340304104400000000c3fc0414300000043144310000300cc0c04411301010d0300c00143041003c043030c1c0143000c000c0c0043010041410c00000300f000c1300c740000003c105001d00044c400300000f10440300c0000030000310c3343c001c00001c000000f0010000c04031403414330003304413000c0001003000310003c1403000f0d0003d04050030000377043000000430000c040000c0701c0c7030007003305c0c00014c004f3340000c0000003040000110001004c0d040c0dc004505c03001d703140040300cc000d414301000340f00c03000303c10003c040010103f0003400c40fc303014003000cc340c00000c00d00c00003030c004040c05151c00000cc1000130d43000010030103030004c340404c100000000030c30000100c4300113000c330c04f0000410300c001030000010cc3500001044000cd00000c00c003000030000d40000400c005400004430170304cc004001400004370010700000003c0400c03530c4004c0000;
rom_uints[288] = 8192'hc000000000010c01000700000000c411070401000000030300c30000c441040000cc00410f300000000500414400000c440303010304004300000003070000400003000307000300010000010303c0400f4070031314000000070040c00033c10000c101000100000500000003000f0c010c0c0000fc04c30007410c4700000100c3000001cc000000000300400000000d00000100000d03330000000000c10c000001000000004d0000030000000003000354300000c0300100000474330000000c40000400000444c300004040c3400100030000444400030c0c40cc0f00000000000c000704000000004f044000000c00c3000003000300c0c00d400000c40f0000010003c100c0000d01c0440c000004000431010000c404c3005100030001400300cc034140004100c10100c741c00f0304300003000000010030c00003c000cc000c0101000703c001c001c3c041000c000004040001004000040c000c03030cc0c0070f140400040007010003000c040044033700c04000010000400000000000c144700c0000c040000303130300030f00000cc0010f00000000000000430c00c00000c3c0000000000004400000010304030000030c4004c0000000c1c300c0000c0003004c0003c00004000033040003010707000c40000043050004010c01044c0d0000400c0000c004c004404400010303c304030000c0300000000340c7c0c7c00100cc00000040040300c0c000c00447000001c704010140000040043f400c004100030003c04001030000cd03c003000cc03c00000d0033053403000001030c0cc0040303c30000000500030c0000030051c001030c000440000400000700030041010304030000001c0300d40133cf0000c0000040000400400400010004000c00cf0f0c0000c403410c0dc10f000447000703c0d0030000070300c001c5c0400c010c000303000740c1c103c400c00300030000000400003000030000007000400000000003c00c00c14304047000c300044404010004070c0040cd004000c0000cc701c04c000000000c0043000001000003040c00000040000701000000c00000c0040305c30003000443c000c000000400c003000c0000430000011040000003000c004340000000c044000c000c0040000cc0004001000fcf0c0000000000400000cc0014000100c004400c041730000300310003000c0100000004000300400000c000c00007010f000000c30c3c3c0100010040c0c0000000c000070003000444010001040700000300000300100301004307010000000100c040c000c00100c00043c000000003c45100000c010000000c00c000c0010000000300c443000c40010c000303000050003c404c0f000000010040070300c300000000030003000303c0c1c303030d0000fc0004000c040043000400;
rom_uints[289] = 8192'h40c304040010000005100304c0001c0c40000000c00030000c1000010000010000004fcc0414000000c000c40c030c000430040103130034c0c03c0c700003101400cc113001000000000100000f3000040c00c0003c40c0000001f000f10400044440000403000000050000007ccc1c0c30c004d00000c000c4300cc410c00cc400003030f00010000040003000103c030000c0000000000c00700d0c0003030000c40c333400000c0000041f343c0c300000c000004cc04410000330c0c0003710c400000400c4d0c004103000f0000413c04411010c40000440c40c40000034100030c0003404c0004c313c0f3040300ccc41c00004040010500030000110c40000c03c4c004c3000000000003c003cd030c00000004400fc001040c04000007400000c000c7c0011c410100c00000000007c40000c0c040d0c44d50c0c3010c4001c3340000c03400000d0040c330031c0040035004cc0444000c300000c0100fc40d01041c0c073dc0007100c044cc000300c04d030c35300010000c003100010d0f43000100030000c000cc0c040000004000040001000c130000cc04f0030c04100f00c000c0400004044c30000007c0400000000001c344c0774c00000100040d030c0f400c00000d000c00c003000c0c00c00c00474fc00400044040001c00c0f00007404dc40c1d0010000000f0034000c10140c30000500403011100040000007c13c0c0000041470300001040000c000000c1f010cf000004000c00400005c001c004400003c0030f4c41000000c00c110100004d4000000c00000000000c0c00000000000c00d00000000000000d03c00004100cc00c0c000003000100c300c0c04c03cc000440000c0003c4034003030000410300030c4400c00d4000cc000000c04c00cc1c00410310c1c000f403400cc0700713030140030ccc0701001c0000410504cc04400c01330c051000000000000001000030010000cc0c004100c10000400000c0000003040407070404c00140c00040070100400400010001000001000000504117000000300000c00000300140100000c00c001040cf00000d004031440000000c0050000c00070d0c00000c00c4404004001cc3c400010304c000000003000c03000300044004cc041003c00070c0000007000c00c00704410003000300f40400404004305d000405c003c30301000001000003700c0000040000740c00004f4040040c40040c01c030f0000300044d5000000000d30c0100c00004c300c300c141000000000d100c040005000c00ccc300040070cc0100101400c0000041400000100000030401007f000d030c00f3003000010c444c300300000030c70011c040001c07c0c300000303037044c0004c0050000000000100000c004c4c0000003c00300030c0c0c1c30ccf000f0043000400;
rom_uints[290] = 8192'h10040c33f0f00003c01300000077000400000001041040c101000050400f007040333dcd010403000f030c130540c0c00004033001030cc4000003000013000031001030cf0000000000f7000c3cc0000c300ff10300100140000000013d301311f0003013533001cd3400000307103003f04c7c00c00000310110003c03c10030014030000c0040003000000000000000000030031301d0040030100d10000040000013315000301000000700f50430003300110040000c0003330000d003cd001000000003c30410f07030c00103014c00407100000403003f310030400c000000c00c01000c071000703c00c000d007003d10c00000003000031300013000000030014c107500c10c0010433010005cc000304300034400740c0001010c0000000000301300003430c030103003001010300303033000071400510040004003c000000c0000143310351c01340130c00cc14d41003c00003c00400010001030f03003000470000004100cf00400300c0014f5f01030300c0000043003300c0c0031010c31140000f07100300c140000003000000100dc0307010000103140000c01330c000003140cd4000344c40c0d04303101103730101c0131350c31001000311003304033000033000103133c4000103c000011014000000100103c000047003103110cf10500030f00010000c31f01c01003f0300c00000040004c00010011010000030f100f1001003d01110003313001000f00d3100dcc0d00000c10031f00004410c0d11007030000000030c0f433c13030c403040400703000103000000400000ccc1000c033001313500000300000100130f0300f04c4303c500000300001700103030400003000101004030c0f000310330000000010d3000c010c3330000000030000000c00030cfc40031304013c000111003000703000300031303cc00030000317130141117000d0070c0000d10000c0003134f00000cc0000000000000000040330000100cc000f10c00000000030101f1033000110001000030301030010d0040c1000010001304410131000c00101c01d0d04301c0000034300003cc01031100030001330001c1100000103001110300c1c4c0c0001000100001f3010033430340c4111001c4c0c0313040c30c0007400c003000030001c3004040c1040301010000d000100300c00140c0001c001000000044000017034470000101000d4303000000000340033003c07300410001004041330003070070c30000011010031003040300030003c001c0000043377003c000030003d30010c004c3c00001034101003c000011371100000003f0d0100103c0030000c01330004304000001100c0001300001000100000003001f1004c0310011c00014c030000010c03073f73c0003c0030410003000300010014003000001470;
rom_uints[291] = 8192'h13f00100414000000000000c00c00c00c00000330000000003144000030403000000c1010cc0000f00f0010070001fc013000000c3000c000c00000000040001000440070000010000001c007010000000000000c0400cc000d043004005030c010401034000104f000040c0000030c0037000c00400040001544403004141000040c30c100044000000030000140c400c10000000000100007c300314330000300040001f0030440300000c000005d000c334000003107011000704100000400c00c000f000101005000007071000030000700043d0300100001300c000c034000040144f000000400c00030cc00007c1d110000000000c01000000400000c401d00400004c0007c0c041c301004003c00300000303f0001f04001dc1000f00000040031000c0000000000300000300000cc0000c000003c00000d000d00400c00c0d401030000000000343c001401c704000000c1003c000301030130d00001000000300003000300101000000c00310c0c0100300000001c14004000343c00c0d4010d050000000100003000301c30000100000000000140000001300000000f43040c0000500000300000013403007d00300000400c004000000000140ccc0c0000c3311000503000000300004c0c00f0300d0034300c00001000f0ccd7041000c0304c300304f00000000100430000f10c040f000c340000000104300ccd00fc311030003010000000000100301c4c41334c0000000341551100000f40004003003300000c000000004030001004040000004c00c000000400040001303cc301001000400000c71043c04000004004005000c4000400100f000000000c00f1100454314000050403010004c050000100300005000014c43c010040000400130000000000c370040004000cd0011440700100010004000041313413000000c00400c00c700300010f04f104000fd4f0433000040030000013000710c0001f00300000001000f000030000000004000030003004000c0c00310004000044300000c000c000000000301c00030070000000cc030c010000043c0430000310010000300040004100000000003c00003000003000400000300000c040300000330004c00c304000070000010f010000000031000003000430c110c0010030c00000c00030000000000c100000303000343330040f0000000000000000c0c000401c075400c0000100c000030c100000000004001003cc000f000000000d0c00cc00001103000000000103303300c141c03c10403004300000000c003c40000000100f1004000000000001d5c000000300010000c00001050000400000000100010040000030c331000003d0300d0000400c4030007000010054d03000300c70c50c30000103014100cc0030100c4000000004003000c03304d000003d000000;
rom_uints[292] = 8192'h4034000400000000c00c03c4c00001030030000133001100c03100000003f4000030c0300c0000010140000000100100103c1004031c04403001001300000400400000040c040c000000010c000010070300310141410c30103030000430310034c703001000001001100000100c3100000000000004100000000c0300110c00000c00011400003000c00c000c0c403030300300011d7c044000143d000000101044000100011030001003001cc4c3034037010000040c3010000c00c00c000430000334010030c40c30144030040c00000000110004f705010000034000003033340000c40000040000030c1d11331033c030000000000001030000000000140c03003003100000000130c0f00d040031744c300030301430300d014054300000330005011040000c33100070000c0c0000110c400000003400000c000c3c0000040040001430003cc33013000c31f04f0000030c001f3145031003000c003c1000311017030c000103cc10300004340c001004303014110f03000c0031070434c440c1d3c0010343100000301c4c0c300001010000000134f410403000c300301d00001000330000100100043c30c344000c04000c3007c300040010300015040013100100f41400000004000333c300311004c003f3c010c010100cc410d00f0100c00c0403440cc00c300010001700340000c00010d304343010040000140c70140c034000400470000003100c1c100c000c00304c04c1030004011003300cc003003070d1000030000c000c00033074101001000030700c0300700c3d70074300100c013000403d00330000140d30011cc03433c0114d4030400030110143d0000d10d0d1403c00000100000cc100140d401c0010033f1430070c04c0100333014c000000013170100d000fc1d000700c01410703c00111000c1401301c3c101410001d143500c0303c04001cfc1c430100013c10003000000c3003000000043030300c0000040003011f1001c010010001003c00001704f1010303000000030034003141010300004000003001100031cc0c04d00c1401170000040c000010004c030c347004000c00003013013404100c000010043c040070040130043cd100107304403c0f0304000404d00410143c000010010000300d003034003000003007c0303000100414040000003004c40304101303410410000c004030100010303003c0000f0000003017000c0704300000001c40100c1010130400040050000033000c3407c010000310303010010005411cc7000cd000003f0400001000107c1f0400011004040c30340c04000713d00f400f00107010000c00010c000001003ff0c001340004031504c0105004000000004001010014103134130000041400013f0510f03334300c100cd41c301400100d34004c030001110300000;
rom_uints[293] = 8192'h103300001c300fc004001000000000000040014100401000001011000000000010000300f00f001000c00300c030000000d0440c403340c00c030030010000c00100340000030000100040104030003000c0330000101100000000000033c010000130003000000000c0d000c0011330010000c33000007300000cc00000000000030000c000403000c000c000300400c00000000000100000000000000000c00000300000f43000000000ccd0040033007030000000000000c000737f30100000dc000030000004000300003000c050100010c0103d00400053000000100004c3000000c4001000000001501010100000404003304000000001f400000030c0400c30f047410001000300000301000300100c03700040c0307000001c40c4005075000000c3004d40c040d003f00030300c0000c0344100000440003cc31c00000000c000cc3000000000510000c000d31010003001c0c0305013c00000c0000000cf000330005030c0c0001050030010305c0000340141100c00030110500c03ccc070010c000000c0c0303300001c040003d0000010034010f040f000000000c30010f0c00c00000000dc000040d170400030c30040400030d00dc0000700c0044041000000c0c003000000000430f044c00c0003003300300c0000470c1100101dc47000101400d04000030001c0050000cf0000300000000030100030cc00c04c7c307100000110c000c4fcc001000003c00fc030c000005500000c000037304000c5004030000010111013c30010301000004040c00300100410000f1c0003100000000c00000000000001f00000c000000000330000c000c00000001cc07000f0410000000c00004000107030310010010c3010000100c000c00000003073100cc10030d01010000000d000701040300000405d00003010001dc0130334c4c00000003c04100040c40000400001d3041000c1c1010d0000000000c01031000c0000003003400000000030000030000011100004030100001011f00000c0000000310c013400000001001000c00000070300300000031f3c00f0d1000010500c03f3000003043000000070c03313030011c003c0000c00d10003011c00000440400c000000c14000000000000000010c0000154010000100030000c3c000f3c0c0000030f0030cc000300003000c0303c00c01000000004030c000c00007c0500000000000c0070000000030000010001000307000f1c00000003300030100f000000000000c00c00030033000c01000d1c0001100000040000000000010000010c01000c30000004010001000000000c10000000000f00000c000000000111cc30c3f00c0f50051c000f0c0004330100100000030d40000003000303c0000c000d00c30005043700310403300300000300000c1c0500030c030101130;
rom_uints[294] = 8192'h13400c3001030140103500c0414c053143050303010050f000430100400431300000f30c0047000000c3000cc007330143d013f0003140c000031000101000c00100d10000c00001d300000430000000070101103444d0000c010f31c005151010001303c111130d1c4300000011041000d0003f0411430000053d035500330041c434c0f41400310440001000004f041330d0c0000cc10003010c0400003300030001c00000dc144044030300c000c30030c1000001000104f0303cdc0000040c010d30000010000d0030011004d00100c030cc30f001d100f0c01400000c00c13500341015300c101c00f403000003c47144314f00000000000c030400c10003003c3034f4043041c0f1341074000310000003dccc4013f04013d5347030107005000000400030100003c0c00c43400c1040c000c30440030000140d030000c000003110503c004000c005c04101055d1704300000c00003304430030000d000040404304c0f404033014c5700001075000300d0004040c33071030110000030340040343044304000000030401103d00000040cc000f1f4c441130c000000cf0c3010d00341c010004010030401000f0c00c000f00170000411f1c0c1010c030c41034c41000d040003001c0043105c00000000c03000300000000030cc34f1c0403c000f00000350f000cc4340c0470004033c00700f001c310000c1c140301030c0d373c0c0500d4011330000d0031c10004f0000004c00700030410030dd40010000c00105c001dc01000000403000c50000c00c30c0100100030004000010000043133003004041c5c431010500300c00103010030013004734f03004031c3000c41c13dc30104c01c40540c300001000000700403001c50f14000000000cc13400400c0001d5001010033cc0300030303004314d10310400404cc113100100010413d00030c0f13044310143710074100c0140f304014353010010004f0010010000433005c0000350000031400f10131741c3f00344413144017c0501005400300300710010000cdcc000c000c000044f1c003040011100310041005500070300100c35043003c0310ffc0371f000c0403000133040015101000100f0c00003000f4cc00113003404310100000000000000c3170d410304c0fcc1003c0c00304000000001c0010101300f11c5d04cc0301f00dc500001003c051f00cf7340c0c000000cdc0043301f40010030300430010c0000cc44003300c3030f10f0f10010005300000c50f10c45010c0010701501c0c140f0c01dc04cc4000500300f10034311140c700141104500c0001dcc0143041000c10000000c000710c04007110cd041d00010307000003030010310030040050104353743c00040fc33010001740f30443040cd00003c4301cf00444000003100000500440500031f;
rom_uints[295] = 8192'h310c00001505000400150404c100003fc30000001001c00000100410c0c0000c000000ff00410040404400c300c3cc00cc47000d000d300700400cc00c0000000001c00c00400c45000000030000cd00000c1f05cc300000d04433c0003c4001400c000030f5c0300100400ccc403c100fcc0c3c0031000d00cc04010004000004303f00000c0001000000001cc010c00440040000300000ccccc300f443000300033304400c04043c0c030c000fc0010cff110700c30044030100c0c000000440cc04c103003400c13004041f400c40001c0434010d0100010c0c40c04000043000000403cc1004304300f0040c0034004330410c00000cc000040700000004c00c00000000f000400005004300000001010fc140500f03040400f400c0004c0010c0000077001f0c4000000300040000400dc00d0000004400003301010407cc0040140fc0fc0100c004000101040300100000c0f003040040010f000c0003c033340003cc000c3000d00147010f0000440004000cdd0340c00010c000010000140c0704000000000c00100c3041f3c300074040000500130003301404040c577c430000000c3000000444005c05000c00101010000430f445000c00c104000003330c10000c0300c00c00440000c07c00000000cc10000440c1340007d00410c000300cd3000041000000000300c000000004110c0434034001044000ccc11d0400cd3cc0010000000c040100041c1c07400c07010c00c00305301c0c00000050000010cc00000000043007000001057c040000400001450c00003000050100000004330004000c0c0001cc033c000005040000000030007004000f04000000003000c000000510053000300400f007cc110c000000040c054330003000d0000300043000500f4000c4405000c500014c43443dc0100400c430400100700000c000c0d10003100103030100d1341400001433034030014fc0130500000500330000410000cc000c0c00000000c0c10000404303714337c100c3000003c0130000010003440030040c0030000c0050000c30700030000030d1400303440000040c050000c0400fc000040000c0003007dc00cc40c0030400040c04c00f4500c40404c0050300100c0400000305300c000c00010cc00044cc04000c03000000000173c0000000000000d4000000d040000100101000000f404003000000c4003cc04443301c0000300303003f10c4001104000031cc01c3544d0000010030000000300000004000000300000004c400dc70043cc0041000013034004003010c07104000c000000443c140000000000000000044310000300000c00000000340000045c4d04cdc000f0003c0304300cf004c0043000000410001c144000000110010040400cc0cc4000c0c0000000304c30401003cf003c437c0c000000c0100;
rom_uints[296] = 8192'h33000004004003000004000c4000004c0000030000030f00030004010401c0003001c00cc100000040440000110033000300cc001103043011000c0000004000000300400000000c00000005c3000000000c000300000d30400d0c0004000c0101330c0c0470000d040000030404c003000130030300040c004c3100010401000134d00c00000007000000000f00100c03010000000010c4ccc00000000030000000c70000331305000cc0000001007c00304400001000000510003000c40300001000000100000100040050003400000000c000010000010fd03401140000040c0000003001300030040000044000000c0c000c0104000003410101000000040000000c0f40411003000010c1400000001c00010000400003cc000000c000000003c10010011040004400000001c1400001000400000c0001f010c003000c300004001000030c0403c00040c000c00c470c40001f3531030c14c1110000000100c11f000000033000000000c100000c3004000c0000133f3044cc00030000005700014003443000c40c000000001000c00007100000c33001c0000040030100003f0001000c00c40000c0c0100000010751403001000000000000000c0000d005000000c000000400010c00d0100000001030c00f10130003c03000cccc400c040300740c13010c3000dc00400400040f041010001c0001cc00000cc34010071000700c30500000004400400000300413c0c400040054000040303101045100c403000010040030300000000400030000100c0000c10c43003000c0c00000010300010071031000034c033004dc00000c031103000c400114c0000410c300c4110100030000000040011100301c0000000440401001cc00000000000d0c0400010001004100000400cc0000f00000001010c000003000010000300141c0143010000400040c0005140000000140000104c30100010c30405000d10c000004c30c00030010001000c007c0c0c000003000300340fd00110403401c010f0030000000300044c4003000000430001004c00c0000c030c030000004f3030004c300000010300cc001100000c0c3040000303413004c300c000030300300c000c00140450c0003005000030ccc01044000000041531c0c71c000300100f0410c1400003c0000000300030c44040017400030303030000003005000c0000000400c00030400000c0500c1c1011000c000c10303101010c3440000000f40c0000000003404030004034000c300c44334004000c40400100044700000c0c00011010000f000000430000000040f01000100003c0041c300c3000301100400000510100c0000400000cfc00000001030000000000cc00000000c00400ccc1c0004cc0000f0140000c703043000000000c40001000c00003c400001c3003c004000001030;
rom_uints[297] = 8192'h400d0400004500c40c340070f40c30c14400000371144c0c00c0740f10cc03000044001c0c15000c04cc01314040400004070c0c001430c04c0c0c404c013140d003004d1014c400000001d30f00c0c400003d0c4c000cc000cf3c0340d05341cc00403340414d0400107d000043003000000c1c04040400530c0413334300004000001041000000013c000000000700040000c0001400700c400c00044c0004c4c301c00c0c07001100f00000cd011f00c3053000000c0f1070144003c00c03000cc001010c40000010100300400017040001000c01010c5410103000cf03000c31014c015c0010030c000fc0414d4044cc00701c3000011000dcc0400000500040343440005114040c10044d0f00011c000fc34110000c30440000000400000044010053cc000f00041000d3005031000300001c1000000c003c000050f7035400101cc0143d0000cd31040001000d4070140500004c0403cc000101010000000c0103400d0f0c40001d4c3c30040c0c4340004c0004140c550000540d00cc110440000701040c430fc0c0440003700c0000000403074070c0dc1013c411003f007001000007000c0c400000d1000c000000071cc40014044030300c0d001cc30c00dfc400fd003cd100c0c30000041000010c0300f00010c700400c0341400003300f0004f0c3c00c14700100000000001d45f4000001000c4413000c00701c004c404004401400040000d3413d10d7004c00fcc000f30c0cc0300000413c30003c003013003001c41d000c0c0ccc05017100cc4c03040400401300000cc00100c0033000000c703100000c040d00103030000c100110c043c000300c103ccc10533040030c47c0010c01ccc044001c0030403110000013c4070301013c4031cc31030010300c400013303003001000c034c0003034400c003c10fc0dd00000300104400100cd040701000010300f0dc004001000c0170c10cf40401000c3000004100400000d030000cc0c0c00001000004c0cc00f1000013c3d0300c3cc100040003c0304011051130cc01000c300f00ccc3001100c40041731040cc0043c341440004d0c7140000000000001000000cc401400000003001103000d70400c4c0000334570455000100cc4003d00c371343d0c4100000c300c00010c01300c300c4434300071000c10014c0001040f0015043cc0000000030f00103007000030073f10010000000000cc0014100000041005d7300400c33110d30c1100100000010010003031c30c0004400040040030d00cc0400000030044c0000c04000000f3070004100c00341c000000015430c00c030000c700c00003000c004100c3c00054c110404d0d01030110f0011010000400004403070117044307c03014c40000400400c00c00c0000c0ccc00130c10344c400cd0c3334d4410c0400003;
rom_uints[298] = 8192'h4c0cc000300003003300400000440010c0104033c0031700004c0f01000100000000001c40040c00f114001000130fc01c00000100c00000d0400404f130340cfc4c001400c0004004000c04100000400403cc00000100001cc0403040c0c300c1300cc0100d0c1000d004001004143000c700c0003f14000f014403010001001fdc10003530000d0c000003c000444c0c05040000cc400001111300300004d0c0170c00d0cc3c00030010340c1100030c4c11000010401401c000001c00c00c041407d0d0000f050d01033000c7103f4300000300450c005f44f0c434330c000010000003111000cc13001f00300c00400040c3034100050001000304000000040000000000cd07c7400c00000c00000c7cc0451c0401104403003d0714000f0c00000013400003400000013c04f104010700103cc000000000000cc3044040031004cc00cf0c0000cc7cd03000c000d000ccc000001003700dddd40003f10c400c0000070c03c004d41d71430007001143100ccc4c50c00500c3000f0c0c00331711401401c30d001500000000cf1731014c0404c030cc41000c00303c000040c4000413030400013103050cf054004014f340c50447000c040c00fcc0400c00400c0430100014000700037334c0503c3f014300c0140040f03d00350cc511d54033c10140300330003001040010c3070c7c3f04300004070c000003d0d0330500c071d301c0c300000c0404d41d10040c000c4f00c005000411c0c000c4000004014c003301430104c4000f14000c0cc4440000d44c30073c0000700040d30c001110000c0000330400cc000f10000c00040300cc00c03040030000030d10d00c0004035010c4c5071710000c0403001100340010013dc00d0300000301010040c4f4000003c4000f0c0473040110f7340740c400010300d41000c50d0004400cd0040400143d0f000c11041500c4d0070300010c0f04000003730cc00c00730040033000000cfc00000c1000d0041f170c07000c30100c007cd11f00011c100010c000000c3103c1003c00c310c000c3000700001d4c33d4c7c00fc01d0007004000300003c0300c00c0003f001004011cd0100010700c04cc0000003400d4c100001005c100c00c4f31cc0c10103000044c40c00003417030043d01c074045331001040300000000100344414c4f010000c103c000003000cc0330404350f100cc303c10000dc05030c000000000040000cc040fc0f3c000c000f301c003000100dc000000030d00c0000011007c01031170c000000fc000000073300004c053c1004000417003300300100000300c01c00f0000f0f00050f000033001000003c0004c000c10c1004c00d0001cd0c30010000430304000030007f0c041001c400033c10140c00400c0540000000040f0010404c011c070c1c0100cc3000;
rom_uints[299] = 8192'h4431000300304043000040c0c344c00030000400c1004100007044114010100000000011c0c10000003300d40000c4104501000dc00030cc11000cc11d00c0400003d000400d0043000000c0000031c300000040cc40d0030c07c00c001040c0c00c00c00001310140400300710000f000fcc04000c140f3403000130100000310c0700cc10c000500c0010004c0d0f0303301000000c03030cc00000040cd4500dcc0000000100000f0400000f000300300400000003000000000011004001000c00001400010c317034013004031dc1000004000c0330003cd14100c0f000003010000400c0000000430010c344c0f000010d0433000c1000040000430000000c1400ccc11c40f1700ccc1f30470000cd3c30430130000f154400c00000033f0100000c047010011100ccc504140c04403040cd13000001000dc0001401411c00000013001f4000000c0cc000400f15c05101103c500d1cf1310000040333000030040cc55040001c0340000000c00f0003030400c00300304c001400007301000dc043310000044010404f000cc70fc00700004000000c00c0300c101cd00c05100040037c04c000010440c11330000000103c10013000000100000c05cc0c40014001003c00000c00400d000044047c0c10040c00004300c300000c1c1400d04313cd0500100c0440f00cc404040f000c03000c000330000001c00003073c10100cd430103100403400003cd0541037011f000000400f43043010000114031007034000d01d300d010430f00040000330100000000f01300000003000300000c0d00041041000004440400cc0103000054040000c1c310034000f00000444000000047003050cc400503c003044c417c101d000000100300010400000540c3404007000000c3c004400c0c00cc00c0130c0041c10040000c401030501000003070c0003130000310010010cf00c000030c00001140cc010c13330030110401c0f01c0d003403004000c00001300000145700c4130ccf4000003001c40003010010000004030000000c43030c3000000c14730044000040005100310c404047000000010311c0000300c0000d00c003cc41dd1c437c000010c3000f000001cc00000043014000004100c10304053c00040054031000043300001c030301c030010401f0140001030000c1dc400011113103d00c000c3003001100f000000c4431400301040030003010004100c03040003c01d0fd01001c370000000344000300f0c0cc0005030040401f31c100011000004c30c0dc0000000c00001c14077300434730c31130133310000001000040c1f0c043000040c000000001010c3000c00305f00000133000cc0103030000100c0003000000d000c0040000c40c4f400c0300077343c00033030000c07003014033007130c00fc00003c000000000;
rom_uints[300] = 8192'hd0000030074404c0430404400441c0000c0ccc0000000044100d0c0c00c00f003f4331c0040130000c030003430cc31c030cc1100100c70000c0c70100000003404000030000000000f0c0033dc34077074f011d00005000cd040fdcd00c01000034c0000004d10c30005000c1014c1000311ddc33300d000c3010330f0040cd3004030400d000100303c303703401c0c00005c300030003c401304031c4cc07400000c030c44d04040cc70003400c43c00000004000c3c0007c00000000030c30c43cc0c1c001c0413010c01c4d0004c000c03004c00d101004400c000010300037435cc01c00011c300d33000000400d130100010000054004044000004000033c1c07000100403d3001100534c3d00c03c1ccc4004004000c0407040c01c30000011c3000c011700c3330ccd01004000d0000000f7c0310d0c40d113f0001c4030000000cc00004d0000c10000710011c310331fc730411010001ccc403030033f0044470403401c01c100c00034c33041000c100c3f11301401c3403000f003c41d0c0050c000cc3004cd030d00500c0c005c001c450700031110c03304030c3f3104540d00c000404d3000040c00030311c010000004c4c00107d00c041400d3c030107c03000fc00300004c0100f005cff043103130c010f41cf0100334401c07101c00f0070d4304004311003337f00040403003cc104130c1050000cfc73000011013400cc003077c1013314c3073c00c04f004d01d0cd0df0147c000f031c3550000104100040000cc10330500043044130cc5100010004cf00c010140d3403300743c4400303300400007440004400010c0c5030cc0030f0f00400133dd0400043c30400d3111d0000430c00c100040004151c0004c037c003d040000d0cfc40ff41c5100410000c0f0f0c4c04c100303000000c010403fd300c70c1100033340d3c43740003c343100c031000000c0110111c0040c404040d13040010000d00010c00000c0f00f0410530cc0cc1100c3340030030030d0c00000014c070f0001004c1c10104340c0c00c1043003010040003030434cc0013410040000044040c00005c4c003313303f001100d00400c740c0010c0004100007000400304000400174044f00030070d00cf700004000410004000000030c30033470ccc0040100d00c40504107c31cc00c700007500000c4000400c3041c003300cc370401040400c40050001c4c105c1333401cc01ccc4f0c40001000015010000400c100000c710010d0000c00100d0f10f0300c01001100d00df1f0c04040d4c4040100c40c03030000700c0700000443c41c000c050cd04400700000010010c01cc1410c7000d00040d0740010f0410004001000d14300003dc4415043000c030004000010703003c010000700f0ccfc00000403cf140000cf004c0000;
rom_uints[301] = 8192'h400140004c4040400cc040401000c00c00000040c000000001d00004d4cc000c0c40005074fc000034400300400c004c0000004400c004400010000c104c0c000c0000c040300c000000c44c10040004401000040000000c004c400c003000000004c0c000004000010c400c0000100c0030c04c00c0c03100c0c0400c0c400c0c01c004000000000000c0443000500004c00000000040400000c0c00040000000000044c0c100000000c000000000000040c0000000c0000c0003000c40000700000000000000000010000004004004c00c4c040000dc003004000cc03100c0300000f300f00000000000c0c100000000c0c40000c0000000000004000000f070c440400cc00040004000c0040700c4cc0040100000000c0000003010c4300c000c30000030000000c001000030000000c004c0000400001000c00c0000000000700040040400040000c1c45000400c3040cc0140c0c00d0003000c0000c0005004003c00004c000000000010c001000000003c300c070c00f0000c10000000404000000000000404c0c030c00c000000004700000000000cd0400400400cc11400000040300040000404cc0300d0000c000c04000000c0c0c0000c000c04000c04c400140741430000c0c0000000007c040c0c000010c004007400c00c040c00000030000700040410400c0000c0400000c0700000c0003000010c000c00000400c0000c1000040c10c00100c40cd04400300c400000c0c0000000000c400004000000c00c40040000400050000000000cc00000000c000104000000000040000c0c040000400c040000c00c000000104043004000c0c040404030304000300000030c100c4040000004c000010c444c00000103c0000000c040040000000030001400c000000c304c4400470c00004000c040400ccf1000001000c00434000004c1000000004000f4f1c0cd40000c300010c0400104c300400c5000004c000000c000400400c00000030c0c00c4000011000400000c00c000c44400c0000000000000f4cd00d000440000004c00040c000004007000004040400cc0000c040cc0c00000000cc0404c0000004000007000000c0c003000040400404044000050c44c43404cc0004010c30cc0c00000000c0000c03cc400000040c0c0043030c0404030c0000000404c00c30000c0000000340000cc0c0044c00000cc00f70c7430000000c0400000000000100000400c00c304cc100000c1700030dc014c410000c000000c10c030400000000c0c0040cc0144c00000000000f000dc40000c00014040040440000c040000400000000000004010040000c0000000c400c0cc000040c7f0c000c00000400004c00000000cc4000004003004c4c40000004010c0f00c01c0000c00cc00000140c000040c0000400010f040440004040000000;
rom_uints[302] = 8192'hc00000413dc00000cd0000300c0040c30104000f00c00400040001034d000000300013411000000c0000100007f0107000040551307c00001000100f010000000000c504000000000041003000010c000400110100403403010000404100c0410007d0300000040030c0c30300010c034103c00cc0c00100c0410000404001303000030d03400c00c000004000cfccc040000000c30030d0c0400040ff4044c0cc0cc04000334000000300c3004000003004000000011d001410404c0300c00100110000c00001403000c510003000d301303300010303000f0010f0310cc015000041c041500000d1001d03c0c00000000c00440000000000030000000040000104d0030000410401003070000100404c1d010300100001f30000c003100000330000d100c10100f040c44c1000000000c0400c510000000c3044cc03004303c040004c030000003000000cc000004ff00140c04404c34d00030000010100c00004f00300c3034301510004400000000340310410000100030404c0000030c000d1000300000017410003f000000310000000000004001033310301c0000010050c300104000000c00500000040404003003c410440c000003000000331004000000133050140300c0000000003c1503300303401400000114000f050c350000000100000400001000011000c013004040003400000c700400003c00000f43100000300030001000000ccf0035030f00043000000030004100103c00103040c5000100010071440000000000011f0003303000344000000c41400000c010d030000035cc3f000c010000701dc00400f0100c00000100010f10301cc0c0410010041c14c00001000000010c00040f00000c003010140000c00c40014007014403004100f003000c003040034c00000013000000000403c004400040c0000c010000400011003403f0c000003f000004100004040cf03004cc00100c0c00000cc003000c0000c0000050000c0400001000c031300ff4c30c0000041c4014d710300c040d040010000400400c10c00007c00000000000000000107100300c4c0040041c4f10100c00c04030000c0c1c73f000300c3000000003301c0c0000d004140000041000000004c000003110c70c00000c000c33004000140f1000400110101000303007000c000044cc00d0100c0070040c0c0c3000400c0000fc00000c00000000000000003000310040000c00033300c0000c003d3070000d4030300c340c0310000c000300000501001000c033300f00000000004001f0073c0000fc00500000100f00130c3000c40c040040014400d00003000014000004000c301040d017100310001c0c010400040004000100c00005f0d4104c4c040003400750100400000c1000301700300c44040103030d0030030c0411040035101030000;
rom_uints[303] = 8192'hd000000004c10c0400000300c00c010c00000000004f00000001000003000000000000500000000f004c00500c00cc00004004f000000cc0100c1000000004010400010431f3000400010d00f001c0030000403cc10f01004400fcc000f0000000100c0140000004000140000000001c0100004100000d000000fc7040103001c43300000c30000000000c7cc00403c000d000000040030d014300c170000000000330c000043000cdc300000c0400f5413400000cf50c30c010cc0d000000c000d4000000010c304c00000f3c3cc100100003000500c000000000c00011400c34000003f130c00000cc1ff3cd04000001d01f0140c000000000004000000000c004007f3000030510400300cc1c0c000100040d00000c33000000c00000000c0c51c0000cc00000000000c0703c00004050500c000010c040c000c030300c0400010401041cc000cc00005000004100330c00100044301100030cc00000d00000300100344000000047405040d040003000c3f0c4074fd0400000001103000340000004000cc0000300030000410110f0003000000c00000f000100c14000040cc04000f0000300314400c40033f0c400004140f00003030001001f0004cd0100000004000040c00c30000100000000c0000004c130c00003000013303000d3001d10f00c4100443400d5000030000000c030440100400fcd000c0003050400000030f1010050001105004407c001100400000034000000c0311010400c0003300000c00134000000cc00000c0034f01030c004c00000100000030fc00000000101000c1140010043c00000c01000000000430100100000051140003000031c0004030c000130003003c000003000000030400c00c0001c14c0000c0000c0cc0f040c10c0000c0100000c1051c00c0c303c0cf1cc040c0004003035131cf004000000c001013070c4c401000444000c0c00f10100144010000014004004000c04344003100001c034000d0001cc3000000c4050400cc70700003cf01cc100010000c00cc0110100000307100310000000c000330040000004043004c0030000000000c0c1341300c40000000c34c40030f11051500000000010d000000c044030c00400000c030003000000000c00cc00000f40301000000f4030c0000c0000004001000000000000344cc00007f0400704000000100c000cc0000c10000000431f0300c30005030f0100400040004c430134040130c14050100000003000405100cc15f000000000000000c0044c0040000040407010c0000000400030030000f0044000055cc40000310000c000000cc0c003d00070f000375001c00c30c00c010073c14000c0100054d00c0000c4400100000c400dc044f4100105030430000403c00000f040c0c4003050c0f00ff0040000000000010400500140001c0;
rom_uints[304] = 8192'h30000013000004000000f0044311c0c0013c100071430010004c004c400000030000000cc03c01f50104f0c047cc170c000cc17c130fc4004cf001c03000004003000c50c00000000015dd000400c0f00c0c0c044500000000000c0cd00c00005c40c31400c400004300404d3001c00043c4c0c000000001c000000004001c70034010c0c04000c400000330000000011000000000c03c10c000c004001300cc30000001c000c000003030114c0010005440000100000110300c30000000000c70003c001f01001000000c010000000c44c000041000004000c0c35d00000c0000c0cc0400000005400c14740030c00040300000000000000004000000001d101c003004000c000d30003cc50010000d000cc05c0030003000030040c00004d000300040004c000cf4500c01030004044c017c004400040c300000c000000070400001030500041040005000000100007010c0000c7300c003c0cc101000c00310c000040044f400300440c000000000001100f070010c03c0c3004000ccc01400110005c000074300c000000010050000000000000c00c03004000400df3ddc0740f3300003400000f00c00cc044040000c40100040000c10f03c00cc4010304105040c30f0403c00d0004000c0c143003004c00030000134c400c00cc0c0c0450500010500c00400d00c01400c70c0400003030104040104000d4000404c0030cc1034c0000100c030000c04074c0c3101000300c40401cfd4000000c00005003070330010300c001100100004c3c40cc0400c0100cc0030d004c000000000000030d0c000001000400044545001c001400000100c1000040000404010704d0000170000004033010c1300000f017c1034043400c3c0100000c3c0000700337001140000030000f007303010c01010170114000003000050304403c1c001400470030400007c030f700003404103300330c01003710401cc50005c40040c1c0f103c0000000cc040010340c01000430c351000c10c40005003740d1f00330000001340c0c01500f000000cf00c3f300c100400010040000030c040304045400c004000103000000000000c004030031c0c000000100004040300c140004f01c000000004c0001c0c30c041003001000000c007c0f000040000f1d010c0c00c000004000400000c0f1000d0030cc00400d0100100d01030104000044104cd00451000000000c07000c0d0040c00001000d00c04000030070000000cc4001000c0500f00400c0dc10030004f00100c00300c7000003000004041000c34040014004c4404cf710c00000400040c00000040000400030c00014400000011c040000000ccc00c00f0300c0000dcc0100c400c0100000300c00c4cd00000c0031110000030404100c000000000100140413040000300010030003001c0000000c;
rom_uints[305] = 8192'hf0400300001c000100cc0c0100c103003f0030000000c000000d300433010000030300c00c0d000010400001100030000f0003000d0030010000000c071000000000c10010c400c004000c0400004c000f001cc0000f011c000cc00c030d0c0103043450430313400403c1000c0000c00010000303001000f0c04d0040c040001c030c40000000100003001000010103000100000000400c3503000100007030100440100000003003010000c1000031000013c000c300c134030101404d0000311000000c00000cc00c0010070110c00030c0c70000000101073103d300000000c0000010000000030100fd0000d133300311c000300105004c00400000000fc00c3100f5000c000005000d0100000000547440330404c00c00d0070100100000000c00100c013000300743000000004dc000100d450001340c00000f000000c3c0c000103031000013000301c01000503300011341040000004400700010000c030000c7300c03400001c0003313003000400000c00307000c10000000c0000031073d00317100c00100c000001004000000000000c00000100000c000000cc14330740c0c00000010033003000c0140000034000100f00000030000000101041400430000000003000c001000d307c4000003034c001030000001004c000000003c43031004010403700400000000140000c34000010000110001c0c000c0c43031c30030005401034c1013f1013f00304000000c001c0003011000003100433c0003000310030100c000000044034013f0000dc0000c050c40047f00c30000450134010301030430100cc0000300500000000044000000fc00000f0000010440000ccc100c10030001330700000003000040340040c043d30000440c00000c4105010f003000c303031407c4cd0000c700cc0030000100001c0000100414500c00000000301cc400005f00100030000c000004101034030001000300c003010000000400000000130040003010330300f00000c000034c40000403004000cc000301c0c1000d0000430000074c0043000004000000100010000003030000000007001c4f01c010000c3000000c03001003300f1300400030000c0000000040c000000cc000000f4c00000001143c013010010000c030c00c03040c00c404410000c004017300c3001f0000000000030010400c3000301104000000100004f50d040001000000034014007000c30100c1c0000110030f10000000000f110dc3030d30000010140000c034c031010310c00017100c0300330035443c03001000c00030330000140c00010c450c00c0004c300c34001000040000004cc0000013000033301cc30000c047403701000003000007003100310001c03010040d00410440cf000000000100034010000c0001000000030c1001113040c003000030;
rom_uints[306] = 8192'hc0dc0110c101100010031000c001c110000430d400000000c014101031100103004f01510c47c00000000110c004cc0c03000004300000530000140c000030030c00000041003003100040fc1df004030000001dcf0110330013003000010004000004004000100001cc00010c134f0c00c3004040704c00030fd3010100300c10c0d0031040000f10300030000010033000000100c03000010c04700300000301031300c004143700001100c10100314010000d000003cdc00010d1005c0100003300040000043000001000030100000000503000000000c000010331c0c00c40f3000ff0c003c000000000033300307301003000c40100f400c00100000030c0c0c301000043c4130c0003010c00004103000014000000335000030c5d101040100000043f0000000003c003030333040301d07f000000f000000003043c10c000000003000000ccc000340d000103000c33730103c7330301c04d0400c003000000033305000003c05001f04c0c0c0410003000010d4311510dc1c000c1c030033f0100000010000000003000ccdf0000000300004100f05410310c0d00000c13d4000030300100cfc3143041cc01310c030c43401f00f50000000f0000303c0c004401330d03c0cc070350000000314f0043f40301100010c30c00030110400001004100010300ccc30144100d00400300040301f004c01100403100c0c0c0003040000c1103403c0c0113170cc0c00003f3cc00cdd0c0000400000003300005c5c030cf010000c10c00c00001003003000001d33033c3310040c00000cc300003c00000d00c00000004010000f0f00411000034000003c0700c3003c50c000c001000000010c1c04c00c000115d000400000000413c40f00010700304f00000001c3c000000330440c001000300300307000df000110014070330001c005c0f00f40030000dc1004343034c007c0c130303c040000c01c005330cc001014c34cf3c0100cdf3c0c00000100f00000c000003333cc0c0003003101011c000c3003000010003040301334000000104c000011000000000c0005330d3004d40030100040f0114c3c104014c000030041c00140300103100c013030300030040c3cc100400c40304c000410430000c004034c4d0334f0000f301011315050c00401001c7011c010000003c00040ccf401300c030304f000000c3c010f307f00003040010000111c4070000c01000003000003371330000c040700033c1c0c10033cc143000300300c4100000c00c300dccc043d303033c0037004501000000400100001040c00300c0000c0170000033007003403000704000000300ccc00100000fd00007000c130c400300304c0043c10000030073000c00003f0743050033000f0000000100c0000d000c300001000000000000030f000c07303f00000003;
rom_uints[307] = 8192'h40040000405c00000c001000010000000c0000000040340000301c000000c40000000013c000000003300050c00043004010000004310cd03cc30004430001010000c000c001000403000000c100f0000014003c00c0340000c400303000c000015c40530000000040c0cc00100300c01000c000111033340000040700400c00300c00c0401000013001000003001ccf4000000000000000c000c400000010004c40104030c00f0101c003c037c7c00100c4c00300103c000001c0040030c0003400001010000c1005000001000400000c33c03c0004300104c000030070000004000000c0c30000011400040140c010033ccc01c030000000300000d0000000c10144003400001001040c00c0030140c41000c0c00000000000001d0040f013001c0000c000400404400c3004000000000030c0040003000000000f01c300c300000000c0703000c0030000004300131110000010303010100030001003000c00030000000003c0d0010f0010300003c0c0300c040030000040010000303000405c040004000010f007000405003c40d00000f000c03c0c00c000100501f00c004500000710000f000130040000c00400001333000000703f30130030410007100000001d0000c030000000c0000c1004304c000c0411003000040000101401401003d4003000000c0c43c44400c0c00cc0341c00c03000000000c033c0c10410c034c1000c301000000c5010000100001010003300000c3001c00cc450013000001000c4310c0004503000300000cc104043000005c04c04030000000000033000003014cc03103003c00101000c00000010300400c0010004400000100013000000003303004f3c5c00c0c0000000000010cc43c0f071c0013000003c340000c30000c0c03004001d40047040700377131300c300700000000000c03041000010000000140c14034000cd4400033030003000000010300000f030c0300000000030004300000001c0003000000000000110100001c000c004100c3c4010f0c00000c0010030010030300401000000000000430334300000000700300130004c003c40000c1000c3000f0000000000400430000030000000100400051341f0d030040043c17013000c030c003000100000c0040003000000400010003044000011001000300000004031004c1010010101003110300053000000014100007004431010000400100000000300010c00004000003503031004340003700400c00030f110010010c0030c0c304001050c44700000300100cc400013010010000030010340000410000c00010003040000000033407c0000000003000000400ccc3c00031d00c0000004001000311001000000000000d40010c03070d3100004310000c000001000f000300000000000c104000c010013c0c0d000cc0110000400;
rom_uints[308] = 8192'hf400c0000003045003073cc000000100003c000004000010d000c00300033401000000030003010c00cc00040fc0c00c001000300303040003c001400703004001000000000d40c0000110c000030c0000100000030050030040c03710000c0003c000c000c300c1003c0004030000c00040000f40403000c0144c3c00c40000400c0000000000000100c00700000000000403030000003404f000010101000f003c430f0101c403000140011d00c0000cf0c0000000c00c0c0003751044000001400011000c00400c00003300c0000000c301400c000000301400070000c0101000004040004000c00304000000c00000001003000000000000000003000c00c0050000000d0ccc100040004003300c00300500300440000c0000c3c4000300000340010c130d000040000c40300004000000000000001110000cc0c007400fc4000c00000000c1f000040400000000304c034003440110d043000c004000c04000430100030000c000400003c0400005000300c0c3005c03001101c0400c3003000f440c0000c000030c00000c014000000000030043004c0000003000000401001304400c400c00c30400001303450000000001300000c40001400c1100400003300140000000000cc53f000f00003400c000000c0004100700c30f031100300c044000f30140000000100d4007c000035000040041cc10cf41c053030004c0404cc404cd0401000f000105c040000000000c3713c00300c40001c10000400001304000400f00000007140000030d400c01430300003004000000f0c00c4000040100c043c34000000000000000001c000000400300c0000c00000300030000040030003040001000c100040ccc001000001041000003000340c1000c0c0000c0000f000000f003c00055c3c0000040c0300400014340000c30701000145040f40101c0f01c04000010c1c0400400400000d00f0001034c030040044c00000300004000000c00000043010c041c001000010000000000401010c00c40c0004c000000000010540000040f000c3000300003000040cdc000430c000005000400d03000100000c00004410300000000c000c005000c0300c3000000100400c110000104c4070c000004000301000040504000400003741400000c40c00700014043000000100c0104114000c1513000000700440000000000404440000000c00003c00000000000400044c0cc00c340000f0d40f000000100c00c01010c00700c400104030000c0404005000041000301c00304ccc00cc300000003004000000d000004c0400000430040001f00c0c00001c0003cc00c014c0040501fc3400d0c3433000147004c000300010001000001001000070170004000501030000003100f30000000000d00300470c000000000c00304000c4d0003100;
rom_uints[309] = 8192'hc04100001704f101000400410000050330153004035130000401300043013000000cc003001000000004000cd0c0cf300c1d0c10dc34300f30000003040003c300100c3d0c000c0304000c03c0c04300c300400530004c0f3c1c000000000010444c11fc30001130000c00313030000700000000404c03350040040cc0444304f000001037100040100000c0010c30000000000c000001401003000010f03350000c0000030fc00731403100d33000c101010d030000c00030c00040311c04f000110c0030000007003400c330300c3100070700c30000000d4f0003d007301403030003031110000001007100000005000d0d00d00000031400000c003000000000f00000053301403350700c0c0040030500013c0c31014f0c0041040c0000000004000d04c003304040c404000000c0030303730000000447110040f3334000001010000003003001041034000100f4000c400040d0300300df000004040d00d300010fc0000100004400c0003000130000000000100c0030000c0000300034333000cc104000040c3410700d070c00000003400003000000000cc00010000031010000c000310070d000c3000000001000004710c1000c000c10011311010300000043000c1fd30000000100330cf1cc03401004340000c0c03004014001500000073c3c031403d31c0f0c0007013c000031c3000000030c0000030c3c03c000040000041c00400034010c00000c01000ccc00000330f03010400300310000301d03c44400cd00101300040000544000c000000d0040031c7040040004d0030cc00100000000c0040000013000c0000001330003370301c003040300003c000c000303010c00d3c00c00001033000100c443000303000000410c13c01030cf0d03c3000003000010000ccf001400c7010001000cd40300100c00010104003503cc003400010000000004cd000104f4100000c0430c000000c5033130004034004040000000003000d3030c000300c301c001df00c0000c310110000101040000000000c01000000c000c07000000000033000cc00c000007400300000000c3010400403501100310000000110010c00310107101000001000004530100c007000013000000300035cc00000c000c00130000c130410003000040c0313304450d10003c0003c0300101300400005004301004000004003c00010330400030001030000c000110d04000001d0c003000404000000000003cc300c000001c0031004130c0037303103000031c000030d0043010c3301000c0c030005c0d00043103c00104c301c3340400411f0c1010003103400000000404000000030730c0100014334040c41300000034003c030401003000014c030000c0130353d0000003071400047000000041000000013c0737000401000030100c00033003000400;
rom_uints[310] = 8192'h10400000c410c1d0000c1400040470c0000f000000001c0040c0c30000070000700030400d31000040010000d0004c3c13cc33c0040000400013010050000003310034f04dcc0010010000c10400100010c000c114c00003040d400000013d001147cc00040003000300300040303300000000000cc000f00004003d30000301c4c044000010001000400cc0030001c0100cd000000040005000000030000030043030000000400000300000c00040013103c04000000cf10c040053100330000004000000000cc00011c3000ccc40040400004000000003530430c10c30033000030330c00000000440003000003003c013431400100001c00000000000000500101c0010ccc00000004433104100030c00c000314d30035403000310000000000003000444130000043c4074000114003113d0001074000d313000033174007c0010340c000c00000c40030c00400c00000000037034c13304d0c0c001004003011404100130c0c00000400cc0003000300043c000000c1c00c0c1000004cc403301034000004001110040151c41c1c000300100300000403034110d000403053c0cc00cc1000f00cc507d100c0040101010400dc0000000c00000003034010d0000300043007000004c00310001400cc0f1401c0031c30030cd300000003000030c000000d130010d4f1000f0c00330000011010d1300c04d00003030fc43cd4000c00c1dc000000001050017004c1041d1000c040043300cc410c03103140430f0010d40304000433004040001011413c000404c0030310c404c1300100400001000300110c0c0c1010c3030c01310d00c40000000000410c170170c4000cc000000f0010f1440c0303d0cc0433c000c000000003000000030100300c0100300030101010000c00c101401c0d40c11c0700000c7040400033011010000313c003140033c0000007431300507f00134d10300fc00000c0c104310000c044000300000000000040301000c00c03000000500c1030400104f1400f0033c0c314300d01174000000000c000410030c0100000c00300c03001004000100300c000f003450c3000fd000000c3500304c00c004001304033c000c4000013330000004000000040c0010005413003d00301c0000130740000011c1001d015040040033174d13000040c000100400f00301c0354100350300c01c00410000000410010300303100f00043000140d0c0000013c017000010400131011000000030d71000c0c003010c3100100c00300f7010000300c7300300000003134c40100000c4730001040c30c0cc00000110d0000033000d0005c0000030313cc00010000c00103404c00004330000007000004c000000000c00000003c0013004c43100000050c03040c017fc000000100043c00c004c0000400c0c00004303000033004000;
rom_uints[311] = 8192'h3300f0401400c00070c040000150c0f000f0c001c01c4f00d0134440c0400000005c704000000030005040377070001004000113040cc01330c000037000514000000f0cc0d300c0430003130c03000004413f000c0303000040031003c0cfd400013043000340c40100430000003cc34004000340dc0030000cc0d04001500000c3000410c0000c0300030001001100c00300000003000000300430144d51c07000011007300011c0cfc131dc0fc0104331f3d00000000d030c00010750030314d4000000000cc05f00101c4300c00c037c00000f4300c000171010c00c004000c000004000400000f00030133f0fd007c0d0003000000300101000000000001300000000000001c70c075c010dc40003014143331f1001c411f0c0700000014003300010100340c04300104000cf0013c0c0344304c0000c000cc3c3000010c010c0540401f700000000c750c000c00000c0103050040c40c4000000cc033c4031c0070004000011040300000f4010000010c000c0c3c0535001030033c3000001ff00c7000c300f1000130000c00d0000000300000430030010c010000000010d00000000c110000300d000030100d50400c0170010c01000300440041301030c000114007310030c030040c04101f000001c34701033030000001c404000040000030043c0f0030331003010000014000f1044c00013d1f3000403003053001040033d4000c000c000c0c40440c000ddd0cd1c030c004c0007144010000000000cc0030350d3100000007001033004c3c00054d000c3c30d14c3440003740003004d104041000007030300fcc0c004031000c0f703cc001c101000010f00000cc00440c00070771000d30400100d0000c040f01000104dcc4300030300000011c003001340410303001101c0000373c100100030374000143300030c00d0000300d0040d1c4017330c430147001100101000000f00d00c033333000000407f0003c00000000040330030030030070054030000004cc0f5c0311444dc004340004c00430f00000000000d0031003000400001000c030040010c30f1c0c300300dc30000f0c01f40000c0c00000f00c00400040000100140c0c000300000c351101004000c0004003100040300c0c5000040401344000107c000003004430000414c3003000700404010000030401040400470340041f000074040c003c3000c101c400f000000011103030100004043040fc400000c010f0004000000440c0f00c00003004030300000000000000070cd00004400001030c0d40000cc400330530341000c1d101c00000340c0001000cc000c30000300001300003000130100404103cc3301c00c03410000cd000000000001301c00370f130f1030305000041040000033000fc03c300110001010030133000000c300d000000d30404100;
rom_uints[312] = 8192'h400f030c00c010000003cc0f00000503c00004000000f0c0434c3fc000c1300001cc0fd0070000cfc3c0c0cc1c00c073c040c0707000c3000005303730001cc0531104404030414040000044c000cc1c030044cc00c1300000140010010040400010400000c0c0cc1c140000f000cc00c00000301000c0001001000400cdc00f0007004000000cc030103000400000300000003000000303f00300300441c5c31041c0c00c04004001c303c441300140014430000300040100c00000c01c0f03031040f3c0014403c300000000c41011070310000c4000c0401011734540003070f0000000f000100500003431c000c0f001000130104000301000413000007d0000000001c3c0000c0c031004c10f0034000130c3000c0c3c000d400c03173004c0c001000010040350001040007c00003000c07533100000005000c0500004c00003cc3fc13000300003c030c001000c3c03c005c043cddc433cf005d000d0130073403f3400350000c00000c4000000443ccccc00d0f05f0fc0030004c34030000004030cc014400000000000541c30001000100050000cc00030c440004704c1100000010c00050034500c00010403003001cc5410c004c0c003003c0005471300000000c001c05c30100000003c3030c000340070f000000000403c00c0c0010dc0350043c04100300c41c0071c000034000014000300f10000044000d44000000000f03040040400300c0c00d31005c000000000047134f3130010f70000000100040001c0070c04cf000040c30334000c0003d410410c0cf00001000010400001130000004470000330000c000c14117430003000035000c01100c43430c03005c00010c00130000c000010c10104040c01f54044c0c0013f35303310c3500000c010c0010c00c303157000c0105c114031000f000d3000400000050401300000c1c00000500400c03c000404105f4140dc4400f0400c10000000cc00104400000000100f301c0c0000033c00004c074010700400300070503100c000100040c40103000000f0c3d4d4001700401030f30400300ff0c130cc000c3003001000053c000c000000000005f01045300000c05000c00000c0001c000105100000000040000f0000c0000000050001c03440100c100c00001005000000300033c010000000000000d0d00040070f4000004003c040043010f011003000304c3c0001000000c1c30033000440030000f0c4473000c00543503000400f7010c3100510034004400000c000040c01c03cc040050c00030000300040470101000000000f00c04451300010400000000c000530c4104000000011d00000007031c0c4d01c0cc00cc0fc00c00cff0c300000437c100001000035334010410c0c00400001c00040c000440000f00003011001700040c1c1100c1100c300500003000;
rom_uints[313] = 8192'h3004c00004000003003d04710c30000050500000c0f040000c4010404000c0403300414000c00430000000070000c01303000c3010070000001100400010400100001010000000d00c10003033301340044000cc4c0001cc0c4000001040c00040f01010d014140d4c01000105000000430000130004001030000030cdf0304010004000140000440401f7c303000000170100100400030040000010440000c0000ccc3003030041c0000000c3030000010000004003004f000003d001403000000300f04000030c1010500341007c0000000110137043300010cc00000000cfc00c00371000331040003007000f04c0c10001000100c000000001030013c01c4030000040c00d00005000cc4100c0c0500030f100c0cc04c000cc000f0000130000000000104003000c104c0304003000000041cc1000003000c1001000410c03c50000100c0d00d00400300c00700041300301000031004400001c40c30100001304300304003c010000010c0003000f00001074003050d01000034c50fcc774304000030000400000041c000000100c0440c000000047000000cc441030c1300100000c30030000c013000133c0300301c740c0005100c00140010070000d0304110000c00c5f013100100040100000f100c40c350331ff00003004000c00300033c010301130013c001cccc3307540cc40c0000c04c04040c0340cc0f10c7100000001000031f0c040010000000000010007000100304400400c0fc0004d01000300000c030300040000c00000000c000000504000cd00c0c0000c413c0000000000f0100000400000100400030000003c01110000011010004050c330c10001000014c04000c00000d31000c000010140004cc000c0307d00004c01330400c00100c4c0000007c100005d030400d0010c0000000001403303400d10000031c0031400400d4001130c001011070100100c0000401c0103003044c1c000000004000c500000103c01540000034010000400001000cd000c04010000100003300500000100414c440010004c00c3000100000371cc0003c04c11c000c0144000030111000130000431003c01400070100100100c0000c0400311010c00000000000c000c0c030c4047000000c070000c0111103c001300007000000c4f03000000000003303133007100430030310040010040d300003400c000c3040030000100c0030000000704000030c00c00000503004dc3004000f0cc034400100000004100000000100303033040000000000010000700000054d0340cc0010004041000003000c0000000000000300c300400010301c150000d04001300371d33740c00c1000000340400000000cc100000500004300400cd0000c030000d0100c000010000030000d1011000000000100000500c1303004003000000;
rom_uints[314] = 8192'h143c0000c00000000000000000033113303c01403f0040400100d1000030c0010c000103000000000405050500000040000300017f00c03040000000c00f4c0c0000c314100100000004100c000c4c000fc0040334000001c0000000013cd0000040c00c0005000c0000000f004030400000cc001cc304fc0300f001044000000f330303100000c0000000030000030003400400011f000504000000001100000100000443c010c30000c001350000000100000000000104000004c4f00000014c0000c0000d04040340c0104000430000000f3c0000300c0000010c0d4003c007c0000400c0000105000100030300000000c0010000000000000000100003000300100004014000501f001001400001cc0000001300f00130000001c07f05404300000c1c0004001000000030000c003c00011f41010000030c000f001050003301000003c40000400000c430000003c00303c30013ccc1c0030000001c010000000003050c00c000010003030040300010000010c0400c100100000007c00333f001000013f00044000100410fc40040000000100010004c700000010000c0c01c110000000cf001130c0000000000400030040cc00000300c00c0000030310c00414001150c000030300d00004430c14000000030c3300100000c00000004000000000000000113004100040100044c00004004010000043000000c00103000c00d0110400340540c00004304030f00c44031003040011005330040000044010000000330000000104003000400030c0fc00003000001c300004f000000033000c0000000300003c510100340010400010300030000000c0000030300040340f003c4000005000700c0100100000004030400000000004000c00f030000010304000030c10100030c03074004400003cc0100413403f001c000130000310303000c0300c0050c00f003030c01d4000c010030001c0001000c000c15000c3040000310000000000010040000040003000000440000430043c0000041100300c0000031003f0000014044000d300300cc000300cc01cc00000010033c0c0004000040000000c03000000000000300c0704000001000000100000cc000050d0303c00000c001c03004001000010103000cc000f0000000000430000040004000c30000f0fc000c4000000000c03703c0001300034c00c01d1000c0004c004000000000000130004000c00330c00100033c003c00130041001c000c0000040003100c010ccc0000043500c300000010c17ff00c000c00100c03c0100000040300000c0000100014000c04000500000f00000c0004300010400400000300000100000c0354304000000301500001c400000440000000d00110000c030101cc0000010001010c4001c0000cc00000050c0000000f00140030c0000003c00001400;
rom_uints[315] = 8192'hf400001304300001004004000010001cc3000400100f7103c000040000c10c00c000c010004100c0000010101f0004c03d000404cd0000000000004c050005000003400c030011040000000103000f0001304003000000c034cd5403300d4c0000000f300400330c003c04003c07c30000000000010c000000c0c000000400003330c44000000040c44000403c0700c700010017000000000d0300c00377100300401000c00c73110c500c01101c000f00004300000000000100000c0000000000350c4000000c10100000013c004d000c04000000d000303331110c30c40000001000001c1000000001000000c5c0000000001000010000000000003c300000011000001004003d04c335040011400c0000000c003c0c00000c0003040300cd000400004c0033000070000004000c4c000d010300110400000003000303000003330d0300c0d400003000310004400c400d00334c00c30000000100000c300c000f000053d03d430300100000000010c400d1000700c0150f04033c3c000c104d050c0000400041030c00000d30300000000fc30000300004fdd00000000100000f4c01cc03000003100c0c30001000000104c3010040cf0c0000000005000001000100000d14340c01010c0f00000dcc00000040000000300000030003040104c0c000000005000000370000f400300d0030df070000c011114c00010030fd0101c0000000003c100000050134100031004100f4430500000011410104000c0c40c0000000000000000304030f100000410034010c0300000011003400c0c000004100010300000304030000c30000003000034000100040c410030000030c30000000000030040003000c00c001c33d3400540001070000000001f3000000000005110400f4030000303433000400104d10040000040000030400c100000c0c000005010040033410c34c40310007030c0c0c000f3c00c10030c0333004c04000c04000000304030f30103034c00d00400c5500000003cf0000040451000403004c0c00113401030400010000c000003000c10000030000040f00c1300c000d00c000c00000400100000000cc000cc0f004040000c00c00400000000c00410000000f0301000c400004cc40011c0000013c0100030001f000050001001500010c00010000c1000000c1c0000dc143000c0004003704400300070003000c10000010c31014000000d0000c030c00070c30004003005f000f0c000000c4050030000c00033c000c04040c0303000d040030c030c07007000400c3000c03110c0700300404000000403010001000003300400004040070c10004430000c1c1c10000f511d000c000000404000000100043c00001004c004cd00300040f013000010040000f3000430001c30c0001f5000300f00300300c434000004d0c030300;
rom_uints[316] = 8192'h4050040000000c0001000c00041f00100c0c03301301c74000f300300000c34000300011300300f03734001c3300000000000c00000003f00cc001c30101000400000144410000103c000004f0000004030000010cc1030000000000400f0101073c00304410c047030000001000001001d00300000c00cc000010130000c400c43030301100003100110000000f00301070010000010303f0740000101cc1d41030510030c03010100003003401000c00057000000030000400300dc00400701303014000000030500000040500030d00005404000004000c000001cc440010f00100000dc400c00010003105cc000000c003004030000000000100d000003030040030cc01040000133007cc1301d00c3000f01c30000100340c000c30003100053c00c01100030000003000004000101000000014000000005000014f00003001000cc0511c100300100fc0103c03000c54700c030100c00f30030000003330fdc100cc5000400003155c0c7400cc0000c31110313410dc05c4000400010330107000140031004f0304000003033cc00000c004001c010034030305000300301011c303c000300c10300030140c0003000cf004c0000001000300033000000430103331d0030000000003000005001cf01110040cc3140430141cc03333300030000100000500000401010c15c3010400c001403013f407300000511000c433070003030000001040013037c110c0c0cf0fc0d10030130000040304173400001330c0104000100000000501300d304c01013000403040010003040000103cc000330410410000440d0040305100100000100000410004000111d00c000c1c33c0000cc7300001041100c0400300001100c1100004130440f003000c000000033000000004c0c3103f031703043010010dd01313d001c0c0005141050000c0c0000030c000c010043f00f00f0011300c0040d30013000000000c1000000003c10030003d0000101000300000c330c40044007c100033000000000c40130300cf007030f1000014001070403000cf0010c00313570303004335000000040c001430740110000c11c100003c0010010000330300510000000040000f04001d10c014003030001310503030dd000000003000113f13170000d000000100100070d0301530040004d00011400c1d00000401100c00000304c3d4d300000c00141500101330100000c033000700c0030f000d01011d0430001c01d000030c1f10304004d41031000000303000000c0030300534000103004000000104000000030000000500000040c000041031030401540030000d410040000104110000000000003001100000000000013f00030000014030000011031000041301001c01c000d40000001030c4000f3040010330d40003000000400007033310111c1000000c;
rom_uints[317] = 8192'h5440400000400100c00000000c034011000300c13044340011c00000414410000030cc03003c000030000030011001c440003033300000c3003300c004000000000000c030c13003100000c10003c00030043000f00004030000133300c0004400001151010013000010100003300030114103c00010030400000300d000001041005003403330333000000005001000100000030000004030053030030000500c300000c00c14030000300100330001000041c00000c0f1000110004403c000300100c04000d070300003000100c0351445c00c01544134c40000104100c403c00000310000030003513034513100c01400cc00c00100c0c0000000100000cc430c401000c0000310f0310341000000c0d0c10000031001031300c000c111014000000010d00400004704c014000c700000000130000c000303c0d0c00100000100c00100314500030000c00040d0c0004040c0015050c300303000001d0053c0c04c01130001c000000c00030100340300000c40c001c00331c1000d00000033003c0c00000303c044000300010040cc0000c0000003000c0001034004034000c10010000000000003030000cc400030033cd0f00300333c40030030743001013000c1c3d300c0007000c0c0001040100001c00100500303c0410000c00400404034cf000300000c0330004110c00103003300000103c0007100001030014130c344304dc00001f0f0414041570cf0740033030c03310310000000110045014000410013043000004034c0001040f3004100000000c040030f103034000301000000000030000001300003010000004100400000000c10173031400101001701030000d100105000000000c0300001010000c34030c3030140c340d0130c01000030000001010003c330c050c0c0004471d010c0030040010357000cc1001fd013500c301130003447d10c307100cc11130fc0010350c003000c40100001000100c0f0000044030f03000000011003415013005300c001cd4103ccc07000001000300003c303000100f030000010005000030000000300000110c14100c300430011040001c0510000c1003000005c03013c04d000c00101003c0000010010c0f7000000014400400100c00001d0000040404003000000050f00003c003000cc010c000300400000070000f00100030003000d0004000300033000301003d1004010d100cc00c001000000030003043f000100cc040303cf5300c000407000f1c01d0000001fc0f00001f0004040c010d303101100c7000310000004c04000000030000000c01c001010c0cc0010100001fc000000c001000450000400001000344130030c50410000010030fc0010010000000000f07401d0000303010031000001004001101300301001c0c0101303000010111000d0c0000010c000f000;
rom_uints[318] = 8192'h403c0000040f100000000c01101000cc000001301000000003304d0430300000003c001c001000000d70001000000d0fc3000000033000000000000140000010000004d030c003000000011c4005140c000003003301c00010030c0030300300010410540000000003005010013000010400031c00340030000303000570141700004030030030300310000c50140000000000000000300c101000300005000010040000100105000000300000c00c004000000000000033504030030300003703131000c0010003144000c3000cc130001070300040101300f00303010010000000000300c00000004001300310003f0010000000400000000031300000010f00100040013400051cc0330c31dc030301f033001003000100c0003100000000010c300c00c300100031c0004000c7c001001000310c0004030430040030c0003000003c00c0100000000100300050f00c04c13330030000000f300301000010004f30004410140010401000300000000c3cc4033433010350dc000000033304c000100c030003400c04031703c00f00300301c0000400040c0010001c00303443d01010001000300401cc013030710000000000000004000000000131c3001110300101000010000300030040100000c34300c003030310033c400000013d30000004000c0c43000010000c30040c000000c005000000000c100000000030000000000c30000004d030000300301100000cc4001400101010000c100000000330000034017300003031300000430040370000000c00c00f40c0000040034f430c003c000010003c050000003500100030031000000001000310430c300013100c300000d0000030400000003f0000013030013001c10001c00000040404000c03300015001034000f000fc000010001737000000330030000c010000440031000000000000000331000040c300001430340000144101dc100303000001000000000403000001030030000000c000f00100015c300003034c00030010003c10c000000000cc01400011430003000013000301f300010300000033010300030401c0c0000d040cc403100100000330c430000003410014300041100000000000001f00d0f30000034003c300000501c303100003001c300030c0040dc000d31030c001c0010100c300100400c00003c40030000f0050400701000400000000003001c0030c0000c000000004c30003000030c30000001001000f00010003010000000000000001001100c0000300c0034000f000000013001400000430030d000000050000401101030001400100007000000010710010000100000000400000000c0731110030000100101d000f0c41c0000013000300f00030000c30f30003c0c0000070010001c04340030003310000010100010050301c74c00131411000;
rom_uints[319] = 8192'h40c300010c013041004043000040c00cf00004c7000cc0000773400140004100c3c03414040300400110040300c300c140d00303c000471c030d00c013000000000701000040c10000000051c00004c01000c144c0c00000004310f340c0f000c03300cc0c04c00c0004c0004134c100400000c00000047001c00003004c0000000c700000010040000000000000400000c1070000c000010300000c70000740400340000303335340c0000003c0c3070300f1400401300000004c030001010000400c00010400f1000000c0c100000103003041c0c0000001c0cc0001500010c370000003000040003000c0410cc00340c0017410000000c1033400c0000c4100c300000000410100004043c341d00cc0c0c004c0c0c00740001cc030cd040001c00000c103c0c300000100c040000000003100001500001005040170430103c00c03000d0010000307c14fc04000f30300004100000300c1cc0040010107c0cc00014070014c0f0d0043030000000034c400c34300f3000d03f00000c400040041c401000301400040000000000100c00c410040014300003700c00c0000040dc000030fd140000c400143030c0cc001430000d044c04300034004010700c400004001c0c40003c0c30000c00003c3c3c1000040c001c074000000c100010000c00c5dc0415330c01c000f44430007000c0000c71c704000c3000c0d00c00cc010c00c10d0c000000001010f4011c0c0004f07030c0043430d0103000c00030dc0030303410000004144404c0050dd0305400040070100070c0004500000030000004003c00001003000c000c00000010170000300c000451540100403014d0c0000c4c4c40000004000c0010003057000c00040c0c040d1030c00730041000000014d00000f00c001301c00004403c003030d00430700010001011c4c01010300400000d000c04303c00c40f00410f1430c0040004131c000c010000c0143c3c0c0000000dc4dc3c0c30000000c000000c0000c74100fc3440001011071c370000000c0c0cc00434100000cc30400000101300c400033000f43034000334100c00051d3c100400000000007c0c00103c1400c05000c000d4000c0044110cccd1104015c0040000040c0c410000010fc004005000040400004d1c040400000c4c01c30040300000f00700000000001014003110040031300c00003030001df010040d7cc00c00c71d44000500f4000000fcd000301c3003f000040000100400041c000c0031001404c0000400c0003c10001c0c400c1004003000007c00000c7c01000010dc10c0040c300000010304003c14140010044c0033001000044c000010dc7d0f0c01304c10c0003400014c400000003400d30d0400040430300000000d0000100004004cc0c0040444000d0400000c0000301c0400d010300d01;
rom_uints[320] = 8192'h310040031030003f0300005100c5400f3040440070c141403ccc0c40cd0cd10043034f500010007131304c1010004c34c01ccc454f00341c40c0030ff400004001011030047000cc0000457f1004c00403504c030010c00070c03c100100f100c10c0d017c0fd00401450001403d410701c3f5000000310f00c73350cc4c0034d144400000c04c030c0030300c0104140ff00c100c010043dd3c011105331c40410cc0c00cc0300000c3c4315fd45f4433c000300503c13c1040003130cf305005000300100f0c4d3000504031030000710040704041f00370c41014014044014151000117d3434140f0035cf0031f40c043fcd500700303c030c04344331f0c0101004c1c1f0437031050053cf37c03f4c3030000314d4c03c40330f0c7c4c010df4000734004c04c01004430303104f77c0333030340031005704370f00c0040004010f03014430c11003c40030305c0741400c00170c4001c550103330c070351c4053fc47c34043f0c341300500c0030007500c44030047050fd07c03004c0403f004300c033f10000013c044d4f10004053000fd11f001f030c004cd00c34307001750003705303010100c3c01130004cf140d001c03004ffd05cdc500540300430004c57000153340001051404010000041403c50104000004cfdc10104001430470001040530530c10c00f040000c0341110400055c0140044015c004000c5f5d344030ccc033c1400d0f10c1004400300045d344c00013c050007330155300f13c0000c00113101c40000f7005710000c3300400307340500000345003d3104ff0ccc000c3d03005143030403c00417f47033341f5c0040c040005f5730000c0f00f01f003003033501c014c3000f3033f3f50d130430000c04103450314d0000030fc7000134011303c504c5d333c034f540350037c403000317007c3043330057400c43300d4f011404030c0cf004044304f3333c00103003c044cc400c0c000000104000f000430150c4030070c1013c33141403c4000343713031000d300444140010f0300c035350030154335300cc30c01014541010f071000101541303f4f010c000104710c30403175000053cc410003c00007fc500041c743d0400fc30f0430c31fc0700000f333c515f31734000447cfd00c30500040f3f0c0100017c0340f0d0100c34035450040007f00303f00f407f040c000000c10c03344074310071c0c05000fd00410c4300170300103710333c40c10c131c330000c44c010030400cc5004d3cc0d3f5310330400cccfd303707fc00fdc00cc0030c03c0f30400110003103cfd113c1d01f03cc10c001c000003030030011337033314c0f043c040cc0c4030040300fc0040c300033c30c015c01d3010550474400507010c3000303043030300c0c04400c41530434010003000004700000c30;
rom_uints[321] = 8192'h1dc0000010541040035c100f03004030050100cf30c0300000dc0c00c0350033040040c040d03f4d4c0f00000f0400f400c050040001d00c000c1c00434fc300fc50701000cc40411000075cc330c00013d07300c4c0300030c3c0344400d0003c07d00c00c4c00c40c0030cc030447f30cc0c0000010047c0c437d05f54c0110770013c307004c00f3000004c00cc373303000300003cd05003f0c430340044003c0fc040000003d0301050fc3f0311d04c7c00001030f0014040cc44c4c0d0111500c00400d00034c5401c0040040000d03c030030c13000c10c111cff1040cd00001c00cd40cfc4c030f0d013fc550300351340f0001c00cc0c4d4400000f43c00471c33c0400f0f033000cc1c714cd3c3ddc000df0404333d0d111c0c04c00003000f53504f100430cd071311d4c30d0103f0dc000000cd470001d474440440001103fc34f010df041ccf3000c7df01cc0c140c00cd1f107100300c0dd440404d400073c01013c3010104c4000f03004d04400cc013c140cc313003000034034117033700c410dc004007304cf443c00300143300d4003cc103f4000700033c035331450011000010c1040f4cff31003057c000c440307107c00f07444005cc0000c30050cc0000000f0cf101c03153c00f00170fd74004c4000403c53f300c304dc30003100730c71cc4701c1c110c03140300f31c30003ff004041001304dc047304301351f00c0c40303700303f00070000d40c00dcf0000030cc4134005030003544000f0004f310540043ccd7074000c0130050031c37c3110030c30404041005cc34004000cc00d1cfc314f0d0000070c14000015c001007330c00f0430000d300014000000030331d00c73440003044fd4017c01143440c101fc4300310c0c0c0c040000430f4c731d300c04ff741dcf45d53007cc00fcfdcf401fd00c011134340c003441015543543cc040c10c10330c03c0c34c1534014030770cc3c4c00000000351c0000000010040143c00fc003f3c757033133f730103c440011ccc37c11c300440cc33031000500c000371cd53401d700400034004110c40c44050013c10300000dc03070111c74303300c3010c40404c3d40cc33000030cc0000000140c00010c1000300353030041cfc3034104f40503fc540c04530c13010300c0030340004040040cd000304c00c33004c0000c00414000430c01400c4100c0040c030d41000300400405333704004dc4d1d300033001150c0d4f1014070c1c40010f073040cc0440434034d0000f0330740c0501c303040f00400471c1d501034040d004100011f0c0040001d41004dc034010c0d700030000cccc0c1f0340d3004330000c004004000100c40c00011c50405c3dcd31000031c0c00010c04f0c0011d101330431c540104c700d30300010c003044001505003c00;
rom_uints[322] = 8192'h5101000001fd04c0001c0f47f500000dc00c011c30300d1010c4031c0c33004d00001c44033000030003000444033004f01040001c34307c30003004340440005030f03c10d110153000044c4c003103044c01c510140103000c075000000cf001f33f30310040730c1403c040c31300000110d300f40044c40c1400400004004d430c00000700f3073000c00100cc700c00000000003c04301c00004fc10000030c00c0000400d0c03000000c07c3000c0040f000c3040003440074340000dc043c10c0001000c0040c00df10310300000c73c0004d10410530000440d43d10413000100140c0100300004400cc7407040c04031c41004f3003000000000010d0445110700431003cc0000300000031405f43000000000413470c0000fc0c000d340f000404fd0001f130001c5c500003c0f0000143cf003c00c53f3d11f3510d4004f00030400133c00c04070c330410c0d031c30110c03c104004303c3c0034df07dcc0040000014c4d010740c000003130c45030c107003d7cf03c03f310340c1c033c033100543000c0414004004700000100001510504c401004103cf04fcc0f001c1300c0000d030000107d000030c17d3c040fcff3c01334000504071cc303c3f5040040031fc0c00c000000434c0000040dfccc50c05040c00001f33440cd50400c0430c40dc10c1c0f0040f403400cc31001004c000c00c0c4010d003c0c004c010000000c00000c0100f000dcc400cfc1000c0c4c34310c300f00440140f0001d001040001403004c101df400c3300000300500f007104033001c0cf1011c701033400cf447c03300c003cc7000c000c400003050c0c0000470307043c0c37c4040c7c104d730d000300c0303fc3110300c1c0fc341c03c00147c033400000d1c301cdc3c00071410440310d0001cc30300010037011000101c7c530100c00d0c000400301d3dfcc4300c3130d04c00000c003c400c3cdc71004030104030040001030ccc030c00cc13014c0ff303c0004cccc100c743040107400c001000dc0c0c10003fd3f7c3dc3cc3c000307c041003000c0c1c00cc0054000c43cc000c3c7c0c730000cc000300d013c03f00000000f0003c0000730000001034040400000c004703043100000034043000003004400003040c010004100004343f040300010c13303107074cd40d0c401030400d01004cf00000f10f134d1334300c101100300f0400017403cc00f4c00cf0010df0c33440005c501c0040300c7d00030051c03300c00041003000c01cc4d00c003500d534f50071031404c0701000f00c1c13000010344313301f307f0c004400040c0c04000000f04300c0fc50f40ff00f074000d3f01434c0c01d100013007530514d04c100ccc0401000030c10cd3d00dc005c0170745c0c0700000c410d0000347574c44c00000001;
rom_uints[323] = 8192'h13001003070070071004403f0030003cdd003000c0300000c3c00440114330000004cc0010c03004143c0001104c4c001dc0f44004010007c4004c03034c04c044ccc003c540370c001031c00143100c1dc0035d010d0cc000005047c400d003071001000500410031cc3404fc3001007c33150400c00000034301c1004040cf04000000cd0015001c0000cc000000c10000000000410030000003000c3fc100311170130c1300304000000c0047d40041034300f1000d3105000001000300c1d10c4000100004040001000c00300000c03035400330003400cc00117c043000000300404000440101c05f0c030000c040345071d3c0100f00c4314000003403743131c000c140d37f030f703c0000403c0c70000000c44fc300055c430c0f00100000317004f0f00400c5c10140d000701040f40c103c0004040405c0c00c04403505001f0300700001d013300070fc7c013400dd014030011ff0044c30c10011003134030c430c0c0cf00c4701c000fc1070010343400c0003000000000c34010531c054f3340f51c0340330ccd00000c400400cc000c33001401100c100f3c500300000003100f440030330d000000344007dc0100c00100fdf00100d0035c4c3404c4130d110c000003000303033000000100140340d430c05001c03c41300400c10110c007c0c00cf00310000c00040040fc004041c40400000c00d30d1000030104c130000377c4001c3034330f01330f100303503300d5000100000d0000100c0c0310000d30f300050c013100077001003c003c0f411001300307c000cc30c31004300c1034300005034033441c3c0c4400c0300303500c3c304c00001040c0710c17c074000c0101040403001701ff77000300f0534401fc400000cd303005040000004d0044d70015f00543440314c1337ff0300c0004f04c500f33400003030f0c0c040c0001133031c4fdd30410c4000c0100100733400d400c0033700d00001000401110001000c70c00f1f7fd007010440000c1040300c00c100c033030401c7000d04c405f1000f031c041040000000c43c0400f100c0c30f04300001cc011743d0f000c00d0000c0430013f001f0003c0c000d000040f14c030130401000004000000430007c4000c0c01000d0000041df3304c333001cc030003400030f0001c4451300004c000404043c00f300430c0c0100c47101033f100c3050f30010c110f504d000c4000033f70404034000c43400d100010fc1c004c100d0000000c00c0030000034300c13000003d35c01c530015f0c005f00c0003df74f400f00040003300c430c00004040100c000c0000340f00404c3043014043044f4fc4d00010d10004c00c03003f310403f0000000c7040c31c303734c000040c33430fd10f3c400005031050c0000c14131704340100c70000c0c00;
rom_uints[324] = 8192'hc0100000c1cc4004fc4000031c01d551330510c50f0011000070050300440001c0c033041014f000f0f0400530343c10cc0400300000003d700c51c00300c0000f3c005010410013000030100d00000001001003c037000337c744fc00000000c3f100000f04c00000044441c0c010cf3f40c040f0d01c3030c00d40c44cc7004dc444f0011000033003000c030150f5d0c10340000010f000d4040000740f5400104c0030c0301041100400d000403c00d0000000130073f0030034354400000c41007031004100004f100f0301f0000175c407104c4000301dd133c4d31000407100c70130c100017000f00050f303000c300c50f00031000400030003000c003310011dcf00d031ddc10003300141f053004001f01000001040104110c0f400c0010041f300000110f33004437c0f004100c010f0f4004330133c1f0030cdc0c0cc000030c40343f710c130104441531f00135005c50103050413003100f1003013c10d4c0043505d05000000007001c104cc373001fc00551fcc4c00400043d04c075c30d1c03300000140400701f00000000000c000410330c00d330400005f000351100c0100000040d014c4030000001c400301d471307c3303c0c33c00c0f330530000f0f40d003030001040310340033f00533f0030c0007007d7c5f1c1d1f4f43cc030fc4340c403c34003f3c00f4170430003d330c040000000d040003500301005c100df0f00cf4035300f50f0031300100c475301331c00d300301107414301010c0001c30034010030fc4d030000453c10c51c040ff103040503c3c000c0730040c4000430005340c30cc4410000000c000c4c01ccd013704550030040c300c0f00011103530c410c001c00c0c03f0510033cf00000c4530300c0300713044001000c7c3cf13050c3303dc4d04300cdd0000c43440c330041003000c0fcc5c4000f134443340004c5331000004007c40f0300017d400c3f0cf1150d01cfc000000030730c0c00cd040004031700403c0055000500030df30001100000040007030c300f33f330005c010705300440304303010000000100f03d00dc1004c340100c0000034ccc071411010f0000100c34330400c303040c504103300c00130c0000430133100005cf10030c401700000c0f300030c00410010c3000110034c01500340f0c0d40105070003000305df03c00030450010c1030001013437705000f0c413c4130c00101400100430000100310cd30040c07033c033055053f04070c04000031ccd00030010030013f0703d301371d000000f043f4100000100107cd30413001cc730c30fc150f000000030f0030303000051c7c30303f3004031d001cc00c03100d3007c0c3d44d000d1000004c7c30003000040fcd300005004430004100700743cc7000000000040443f0c50c430c000343000;
rom_uints[325] = 8192'hfcc4074051c11000034c1100c000c0c4331c00000300c7043110c5000c01c04000dc4154c05f034ccf3000404cc000fc0110004574401071c0000f3c03000c050c307c3704170405c00030c3300033f005fc04040703c30045000c014c15dcc40004d000f0000d03d0071c0c303f34cc0f0cc70f0307f003000f44cc00000d0047cc0f440044000c043c00300000c74d0cc3004000c00c44040731c70033040c7f4330000000034d003c1104003470cd0000410c00340fc30443000c0d071d07cc100005400cdc00c00c04030fc07fc3c0d04400c300d00c044f040c510c0307074100073c0c503400cc003410c4c000403303c000d00c003000cc000d00001c30430cf03f070c00300051431ccf00100dc40d03400c0704440370d4f7c0000000fc41004c3c03cf10143f0c4c0d03000c130505c40001000c0003f0c00540c00d0c535d003d0103030c0301c00c00003703744f3010c540c3544003700ccd0c300314004c040c040d0d11c40c034c3c013c4c0144370501fcc53f0c0c0000c10f040fc33c0400c0c30cc00043003c0c0300c030d0c03500010c000001c04301333703330304c0d000d3c4130d400c010c10004d0c3503040000734133510c0cc30c030034300074c001014c00c00fc0003f00003303cc0c0c0c00000101000c411104100c3c4c03010043c70533000f40003c040dc00cc3000c0530c14501054100c145dd00c4300c10c01f0301443d00d0c440c400003cf40f00dc00cf07300310cc00f03400c70004c50410c004014d7c430000000037dc444100dc0c0471003010040003c400cc4004c0003f0c04100cc003004c00030fcf40c0010100d00fc400001f0f000441c0c0000d5cf0000401c00cc4fd7410ccc30c000103054033c440f00c04c004c014040007dc0003f3dc3f3400f04043030405000c031ccc03430f304cd3cf30c1cd504f10703103711c000c040743cc00c044d104cd0c04040c35c00000c0c040c040000cc30c400040000c00040f0cc0000445000741015000000034c3303c07000003c3041c410c0c44dd0744000c0741004001ccf400c04f40c0c3511cdc0c00170c040000040041414d0f0004c300f30001c30040504cf50400004410c107103fc010c73041cf0d1c34030d004001010cc007305f00003403000f03014500010d00c40c4d1cc300013c00c0c77d4cfc0400000c70cf003104033344001f1000c000354514d43c41504cd0dc04003304010c0040013c0f040d3000000f744cc1c0701c00c0cc00cc00f0c1cc0c0c050c04404c3fc0cf040303040c0c1dc300c0003000f1000500cc00c303034400dc030c007000cf0000304d05007d00010c4c0401cfc3000c00c5c00100c301c0030700010300004500c44040370004074003510f000c0f000500c0070c0c0370d4010d03c0444f3c;
rom_uints[326] = 8192'h330000000003c3cc140000000000151030100000101c0330400010001000cd000100000170003100c3d0c000c0003300c3100c341c11010030000000c000f3000d030441703300370300c0003000d14c33000000ccc0d0c0c070c1c00010300010c4500730000510004010034d0c34c000011030005300cc007310000343d030f1400000c4040c70c40c0000cc440010000000c0000c000333000400033114400c03c0000010011041100033001430c3005c3400000000010533003000c00100053070c0100040101d00001004001c0fc0003330400300000100c01030c04c4004000100c00013000c100000030f0170c310110c0cc0c4001010001d000c0040cc04304f000d3d0311c00000c01c10001040000001001530401100040c030c03301c0000450100071000000070303000011d00d00c050c00100000407033cc10530c1001c000c310c0000c44c00c00053d310040501c04035c10003010100030f07f0000f4100c0ccc00d00010003000000141443d00400001404c10c000033300100341010470000f00010000300000440030c100000c4400c0f0c05c0001c10003103004000000000100010311ccd10330730300030c0c000000c00014350010f0c0c0c00000300000050001000c007100040030c0000f0003000c0411404100f003d00000c30000dc33c073000001000c00310034010c00f040000300004300c0337400011000103000003340d00000140330100c01000104013c310c000d33d0000001f050030400ccc030000000003030000c110d00041c03073c004000c0c130d05c00d10010003c003005530001101100c0100001c4001c5d4c30034c310400010510710310c3011000001c30c33400d143c033300c17c0005d400030c0c00100c0303041003070f03007f414310c15410cd4003c00143030004000100c305c1013100010001103000131010003303f0050111300d1704c400c001c004000000c00003c00c04130c14030401000dc01c0010f043043005000115c000340000c0100013c1100000000100000000030003000004140f0440c00443301311000400003001030f000040000100503304005c01c00050000c0000c00c3d00d000300331c00300010340000100010c0000400000003fc00c004400100113c004000c043103c03400003100314d035000010100000307033001000104c4c01c40300c01010c0000500000000c0107d001000c430400001c0004000003f0000047c1f04c300000f00c4340c000c00050710300000103003001f0010000c01000011040340c10513440100001030010000000100003f00000000340100c000054000dcf11400f001370004000000cc0010030744c00c00c0003c0fcc0000103000c0040f0051d03500113c300000307100100000030075d0030c33100010001000;
rom_uints[327] = 8192'h1c43f0000043c30570130003030003300f010010d000cf3030300f01030000000030d140071100c0000c03000000000c140d0011001001d01003030c0510313303007cf00303100c03000f0401001030d03440d0c04c3041414df30400030c0000d00003f0300c33d00330304071300147400c3001110c00007c3013c030430f3cd013c10c57004c000000d01cccc7cd5110000000f03700d730f00300411311c0cf0310c000d0c000000010c50303c700c40000003410400fc410701340300000d004310033cc3300400004431300000c1c043004c030000c47d0f4d0750400f00100034301010f010000c300003000001f43f3300c0000100c0003cc430034f0c37004003030d1413710401cc3000001c33313d0031303003003330c147001100d700013f0001f40dd03d05005c3114010f11340c00c03c00310c01cc40d0cc3f000c10dcd43c00f00400fc01c1f000003c05100cc01c337d0f104004c030000313040c7f0003440c00cc0001d30000030cf0c4000c343c3f0f3000401030cdc00f043c1d3131cc3f0c00000c174dc0000003000ccc000d3303301c0004110013030001037404f331f04001d0004f00cc004d4040401c030c00cc5c10130c304303301430003d33cf0403034000750d300c0005015001f0c73c030c334443001030000500c354110c011cc37330c377110030304735033c3100003101400ccc00f47140c0c001c0310cc004100011dd00c0110304003c05303dfc3d033c70031d000004343c40d000134c443001040011f000040df4311cc1030300540c3451055cfcf307c000000154cf1004301300100c0304cc07000fcd01510430000c0073cc1c0fc0c03100c3043ccc10100333c07cf01c04d00f000c0d410303300f000d0f0f30300000711c103003cd00403040c00304c3c1d4100f040030130310f030700000307400113cd4100c1130073000000f10003cc4f01007540004f04040303030000000fc030033110000347000001c0000100f400c0433433401c07f30100000330c00051000d0f45305000441300014c404050000304114c5134100003c000000330000cc3d10341c030000010031131344007c0c34000c00c00cc10c0313010d10c10000c05400300c30f40c0cd10c01c300000f003003c13c04030000fc30c0030cc55c333c000c313430030013014100103c103f0000c13f000c0130000f00c00c00c3d07c7005100010300071000011f00f34f5000c100c3104030c010c700003300010300131070003005c0104cc040010001f0011051f3000cd4c3040003c440430040d30f114cc031000f4030d00000000303100000cf03330047fcc4f000f0cc00000000c33dc30030c00c01404c0c00730070c104ddc40450043003033303f0c0535044000000c0c30000000c44000033000d000cccf000;
rom_uints[328] = 8192'h30430005004430cc001ccccf303c447f0d34d3c03c100000110f03000373001000043030010c0014d10001101500004c01000dd40d10fc000001015c0000c4330041735701000c040003101030cc31c033c333144c140017dd0430101005000cccd0147330c07400045c3077000c330d3304141130d04f0300ddc0104f3c000c100010c03f10710073007c0400f0c050030040000000c1f340d10300dc4c44330d310c0100c311474d0c040707031700370d300000003300c700000013000334c10000c3100543003f10d000c0307304f003cc377c0f0410000070c33300d01c113300105031040f70103410703cf3331070730411000040c00c440c000073d343010030330cd40030030dc4030d0010c031304004000314cdc00000504c30004d0300003700d3710c00c0000404304c41c51077c00f0c003c001137100d004f033300c70c500000d03c00300050000070140d3005d4010cc31717104400d103170cc0014000130c0001703047040f01c04110105130403730fc30d30000d0c001f04070440033044030130011d0d71d0004f13000035003d0c414c3300d0c407401d0d03031430343003cc0d03013d00ccccc1033050050330010030fcc330c4c0310fc0010f00373010030003300d0131c001c0003c0040c4470004f00cdc0c304000310001d30fcd0f1001c10ccc0300033c003034cc0000000071c03cd0400d73dd1d413043c333330c0c010dd1414d4104300cf033f4d1c0c0470f4030cf0c14300004403c01cd44cc34030d0d3d04000303411034c43301003400034004c0cc330100341000f0017c0d047c010014f00fc0c10000130300030005c3700dc40000f40000030300f1010043c070010333143030033004c300040100003d0f0c0001017c01f034007c01415505033c44003000400c00010c014d33304300700500030350cc0c034550cc0334c133c0d00c144341413dc4010c100003c0f705c00370300704301001000c000043d0001514001031cdd1473730d00030c100c00030717c1d00f10c1443c0c1011c000c7450400045c300cc000005cc33410400c10034340005c33d4000c0cf300dd10fc115074740000000d110000100c001c30000000104001430304c40010411100d1114140300f34330dfc40c0034300f0300f10503c103104134001cd0037303370043310130013c00cc30040c0c401f3110c0d1400001dd500c007cc007c037d00fcc000051c003c03000007d003074c105507c000c05101030fcf00300f74041403c0507f510057040c043d4f303c0330030770c41504c000103310c0f1100073003f4330304733300c000c3441300073d53d0c7c4c113cc0100c0440100000103f104031003314404ffd0110131010c3050314000010cc00430030107010c0330141010cc3c07d001c0000000cc0;
rom_uints[329] = 8192'h33c0500cc3c3370501310f0d1cc01f044c04401c3137400c04d3c0000c140403d3f537ff14050cf40153000041004cc037c37cf700cd0c43c43300c00dc30c310c00501071040003070003000cc34c000111c043414cc03000ccdf5dc00cf1070153c0cc40f03c07300fdf011c0c0c410104053c0d340304030cfcf3400df1004d00f313c30000f5040043c0000004130441010c0030351d730d1300011f030c4000070304cf11000400040c1303033f51c1c3c0001103100077c05d0000001cc0c5f0050c1300130c5d443300005d7d0300010303001100c3fc0000771d434c000d0010004113000c0700100131714f7340000d33cc0041410044c407014013cfc3000430030104c3c300cc0c1c00f5c0f747531d05c00ff1cdc000001c5c0d1c01130003074113f03400ccc435340100073d0f30144300d00dc530f4f31130f74037d113cc0c04f40f44c30d37030730433c01c30103c501133f001040404d00407400f30047c155c40000030ccd30300004cc40015000c0c00d431030d00434731303f3fc05331050001305fcfdf31100010430000400cdd1013fc30103001034c400c0340d370334100303f0c0100001c4f310710c3003c3ccc700004130310c4040f33000003ccf0c0d400d400077cd000147c140f0000fc000c0d0c11c0103301c11fc100133c31c0cfc473040410303c310cc7540d0004103c7ccc344031cc7c0003cc00111071f0501303d3f47033145337c00f0c0040700110c0cc44104c41003f7c30000310c40cf00300c40f0fc000cc3cff00704430c4d0000003515030f031f1f040010330500140001000303c0c3004000c033f40f003fdcc030003f4d0400300c341f3c440f01c10f400f001d3f400dc05040110014f00c43cd0340001003c33c3030310c0000ddc350f4040413c3000c000cc3030c400017447d0c00c007c003f3c3c1f1c00313dc11f1100050040f131130c7cc540430c1cd03070000000cc0c050100100fc313c03dccd11cd0d41c300041703d40043c0f0000040cf00003000330045030c344d0f70c4170c3c03043113ff1cf00043303701d004311307040c00001d4d000cc0c100c040500370cc03cfc300c150001013d0004304c330d00c1d7310c04344500000c070044050d310cd01f703c33010433f0045c300ffc003331f3c0fc4c74c14c3035003030070c30cc3003007c0031300101c30c00003f04c13c4300f354300f4d30174fc0d00513400f340c000c40100c4100f443501c33c0f04330f3303013130440c0d310037f3414000000131cf0c01ff4cd3c100100103407dc13304004f0f0c4d00c040003003004104100300d33000173030f00030131c134ccc1c0000004100044031c0c05107450355501c0000ccc40f07d30341c300c10007044f4301403541704c045cc103d00c1340;
rom_uints[330] = 8192'hc13d0400c0cc030cc03fc000103074504030311f3311d1d000c0c400c04dc0c0f34f000313374003cd51f03013000d540004073410c300004f0004c4450000004ccc054fd00f01c303003cc04300f303c031cc154711dd00d4000051033013c1c103c1c0c400cc10d1d0f34040540c05cc0cdfc3cfc4cf500100c00fc307f10044070f04c41303031f700300010003f00000c30100001017470c0054007014051f0035001114403700340c41c1d5c3fc0c30c4000004035cf00c000c31100f4000431073000c330d304f03f3c4c0471dfc3c14dc3cc1cc70ccf3f03300c43c0cf73000d00000045300300110453314cc01070f34cc4000530003cccff300f04330c3c13f03c040f044f137131c4c0343c74005ff70d50cc001d040104143333000f5cf003300c100431d05033cc34c010f7300c0cd0c40cc030305143dc57300700007330441550cc050c0013ccd731403cd043030031547003cd033cc0700710000144c4c1f403004317344001044330444c40c14dcfc0143fdf0c05c10700cf047033ffc33c1400f3103c053041f0554005410100005003df34111047d030050c34030d000f00cc05c3734cdc0000d000000403cc507c55c01cc0150755445c0105311f1f3001cf011c300df0001cc34f30010c343c3dc00c4c5433703015f047c050cc0010414d3c34413ddd0431c07004053f05c0003140014f40d7030d00404d0300540c50173000c0000d14331c1004444c00030030fc343030c43c47344f1c475c30100c50100151dc000500c3530171000037dc105403fc004330010c145500c03d0000f05005fc30c4f11170000753c5cc4431004c533c040d1cc30f4100003ddf3c301cc43cc00c4c4c703530303700000003034003430c5f3d31c3301744fcc0300c500070c0511c054cf51474000035fc4104004041f5c5ffc330c340103330033c111c010cfc003305303d43f03d01010013f001f0400c1001c1100c00c00004d03001f0030000330c0c00ff743c440cc5fcd1004044031c000070070103f7f000010340c010004001400111cc00f000f000031d140004cc01c0043cc011fcf4343000507cf300c330317cc40554f33c5d0010445c034413303f015000004034001c30fc07300031435004540751f53d00f0100030403f3f330c3043301c0333d5403c50001c73c10d10ccfd3f000c50c050f300000010cf3c3cf30000000cc000715f1035005cf10f1f7c30f50c070377043d100f40105310f5cc007031c00001300c0003104341c00c011c0040010450fcd03410045c000d04070010473c05307334ccc00c41400c0004300404d000f4301cc00004700d3c00371100f33f3f00440f4100cd4740cf110c3cc10031130dc170050070d00000ddc04c71fc70cf3cc34f00c47005fcf13c10c001070000cc541c030d3f410c07c;
rom_uints[331] = 8192'h330000030c1004330ccc00c41004c01001003004dc3440000c4000c001043047000004140d0c40c403d430c4104c3700cc0f0c043d303d000ccdd44000c003ccfc00007000040c04c0000c0010070000c004001711400cc0441000400c004c0704cc0fc04004054c074730cc4d1005c4430013410d4040010f1f0f0c1c55000303050100dccc00100340040c000700fdc0000100010014000307000cc001c0473cc0100c0001cc0074c004fcc0d3cf70003c30c0004cc00100000300003000c031430433c010404000c00f0000cf0c0f30400c0000330300300ccd0d0cf100130c10001444000410030000c030310304000f43c00d100004010400c43300cc4c3003000407001471f0d0f1fc04410c1c07dc0004403cc000c1d00444033c003004f0000c47400c5cc0000000000000c0300330cf03000004070dc0000c00c1cc003c0c4500cf003500330104000000003030110f00cc4d004f0d014c040cc010400c00411141f7043d0040430004c3c00d31110340c030000f03cc0000040040c00c000dc10000cc1c00000c000031c0500cc000c00c0c00c404154fc3f000cc0730010413f0c400000c0cfc3cc1c7cc30000dfccd00c3c477040cc0c005410dcc0c0505c304c14303cc0c07c0340c004401d004000377000000000d050000c00cc0f700f0ccf74fc0340100c43441c04c07cc03f4c000000033400030c3403c05034310450c7d300c0c00040c0444c100003030400330044cc31310000c3cc0003103010d1c11310cc0000f00001300cc01c040104cc0fc007400c40000000400f003000404100100c440f0001473000100c30ccdf40000c00c3cf30c044003000c00044340401030000040040403054040c4ccc7cfc3300000c030c00340000c007cc4004c0004005f3cc04cc10111cc000444003144000d501044f3ff05d0105c0d34c4011cc0300374c13040304c01000040445100001000030d003003c03c0c030c000c0030c0000000441340cd004cc40107300c14003301050cc3c413f000313300c000430f00010000000ccc00340f470770000fc0004041400c3001f03c004414f00d50c0011c7c000110000f0d040044004100047400031003c301d0c04c0010000004001c00c004440001000000c00013000c00003010003ff0c340d0cc40c71c00000cc5000101c14c0c043c4cc00dc00c07fc0c0000f7300cc00c74400400000fdc00f003000000cc00cd30ccf04004000dcc700c3c0f04403cdc00140c0104c701f04c00f000000040c34404000010f00c035dc170c00444c730113030c0004000710c04c04440cc00c70000c0d00c0030c510c0040700170004c4c7c0ccf3030c000007d01fc00d000041c00c0d4400c01c50c0004c4000cf0c40030c44c043300c003c015f0c4443100000540004cd04504d40500400100;
rom_uints[332] = 8192'hd0c0000000c0000000c1001cd000303c51030000f000407303030100173300400003304534310001030d003003030307c034100c57014030c5010d04c7c00073004c1041100010103000301001041013c107000dc314100014114003044cd00c0c03f4c40c1303010c4313105043730303400300334d000d000403404013100010343130010000cd000000d30c00010f00300001000040003cf300c1400040701d000c0100304c0f0d0001000003003400040f0d00003030300010330f500010000014c00003033410c100071000011c00033001000013f3434c31104330400110cf0043000143400000003340cc10c00c00f403030000003000c3300400001c03c03333c000d000000131033cc30dfd0331000100511000c00000300f000d00000304000403400300c1010003030143d70403000d303000310401000d13033d00030d000330000001000070341dc030040414fc1000531140301100013105f000170d13f0101f04000331dc03000053000041d00730430301300000404001c1c0001734334c3c050f0003030000043f050070005140000030f0c310c400040cc01c300050d30c0100f1f0130300f03300c0d500001c1333d000c00000310474410013003500000c30430300000000c010007007c410d4000000001131f000cd3c03d00500c330d0c0040040c301c0400300041c030700000030000001111350074050c7c0043010c03403030510304100c3150000010c00030110c5000c40113031401d0301c10303f034030c100001ccfc0c000101003100010cc033101c500c30010000540340c0cc573040100130010d0100000000030050030f11010c4103c100011400400010c1300003301330334004310c00401330c13d00f3030050303c0000c010004300310700ccc0033450143c030000001003c31017d100000100501310005145404c1f1f303003c1300f00011c430d40043015d7cd003403003f00737100003000044037314004c400430011f0000030c0c11cf41000f1100001001001040003000041300313403103035f413f400300001c00500071003351c0000300ddfc3001000001cc300400dd310730034c0c3101014000003001f3000cc303000f01c00c5d000000300001400000c00f000c03004c00300d01110000030c011030cc001100001430f000130c070350c3104f0001df0073004000140d0cf3403d0c1003353100130130034500d00101c0c14014040f1c0011c0d0c10003004d03034010030d01400001031335301f0d1013003000c10d3f013c370003dc40000d41401301000001000010300000c100c3000004304040000000c030f001000f300cf3007003310c0f14300001070500030c30d0045031003031c003031100031004c0000300010c0001c444003030000441000100f31c301305017330;
rom_uints[333] = 8192'hd14100003335000000c0c0c300003f30100341300c30000000f0f033c00100001101c00d03c3010040731000d0c03000c0403043d304d00fc3413003300010300140410011001311100003f3c0411cd0030340004cd00cc3f0010010cc300c43010003433100c10134c430c001034040c130304c400110c371d0304000340000000000404040003000c33050003430303033300000c103c04f030300004337000000150300004000110f0043330000011100c0700000107400300001513003c040030000003003000cc4d1d00100001131c0c0c00044f04011410045333300010300007300d0c00000403051000101d0010340d0c130010010c3d0f0c100c030cc03030040d001533000044003010110f07041fc41400030f30140110074400c000c000001f0001300c3013301011d4000f000f00100430070d001c333000011f00000f33370f0000c000041c030105001d010c0130000c00100c334c071007011d0f0030430401303401300003fd04000434001c30040c04300f730103070007c731300c00cc1c0d0433043000341c0f00041c3c000040174c3100030f100c0775140c043ccc0000011d33300430000f0c0f040f33070f330714001000011c7f3c0103010d100111003400003700043c1003303d0c0c04c003300407440c0cf0000301144504303c0cf41f0030cf00033d043c10333d0003300c1110040003003303f000003130000330f00c300c010f3d3f304040c00703f30c10040c3f1001130704010514301100070c04000c00330001011000041700f00000c3f00c0c370400000001003000000d141d0734000c0431000313040000001017000100c5100cf0040c14001c100cc00010f10c0501101cf30300c504031c07000300000000000401353000304c0c0d110441cfc0030c073c0000000430000000010d00070035dc3f330000003007cc3c10001013301c30300037cc10370c10330005500c050033000c0000303c00300000001c000000c007304c00033700300004100d30000000c303000103010c30ff40310c010c00344700343c000034303f0c103d10153c300014030c0f0000300030000400041c303004050dc0030cd010000333040037c01404030c000000000700cd040001100331130dc130043003330c0433040d040f3f130017030110110c0f37100c03134401500303040003fc3000000033c00d300037c40001dc31033c033d0d03000d50040c040004013000000d0d0011010004000400001000310034df0c3c100003101114300110000000300500400d15170c3011007d3005300000100c300dc404dc0300000037003d11000c00333100000c5c14303073303030000c0400040c00f00000011000071f3fc00c0f3330003d00300000311c0f0f700000c03d1d140333310003140005df1033310000310;
rom_uints[334] = 8192'h373c4000c03000c4330405cc000c34370cc1c50040477004131100007c1300030430cc00c3c000cc04000df0031c0044cc4005c030f003311340004c000d0300c0003030007434300000000d0010030dcd00c00040404c0044ccc00c043c0d0004011040000fc0070144c500000c030301c04040004000000c47070050f3400f71d105003f0007040100000c0c00dcc0010c00000000c0d00007dc4004000300c43414c0034500104c40dd00443300400310d0f007403c000000000f000cc00c01100c05c045137441d0017c403c00f4c0040700000f30004cc40c01ff3000010500003504404004004010fc04300700c033503c0c10000c0004c30f0300040130003c0d0307514cc331f700cc000d074f0f10000c00004d1cc0074000050000030300045c1c00003401050f1cdd0c0f1c010f04300430cc004c00007303c01103c101c005010c0cc0034000000403431c004c0073c1005043cccd4001041400300d40cc0330df40414150c001cdc40c11cd100743430f0c053c7c030f00f400344c340d00c47d011c030001c4000c034c441043300001c1c3045330010410c003305104cc100000007c0cc4040c00030c010000044c0c53100f7c00cc0140c1070400000f4000107cf4c00030c000cf00004f400fd30c0000c40000dfd040410404301003cd0000dc30003344000dc400007000073004000303034df00c453c310004034f0d04c001c00c05c4000c0c135d00c345013c0073040100cc0000105400104743c03c4000010303301d103dc110f0040c300403043cc0cc00c30c04000004c0c0707c000d030004c30743400d1c400331d404cc04fccf000034f00c34500c0333031c00f4007c4000003c3fdc0c0c00f704030f04000001101403c000c44000033004070c044f4374f5c300000100100000c13000530040c1130003d07c3030373f000103c070d0140003c3c10c0f7000300330c0c704c44337030440040001f001f0000300000000c0443000c1c1004103c014c0074c5000431303100d0c003400030000c3040400005d100c00cc000347401430130440070000000c01cc0c40c0010d71007000030001df00c01c00001443c400334c100010301000400000041d010003c04043400300500014c013074740cc130000310c00cc0f0c000010f00000030304000341c4130300c0040014300c0c0c004013000f71c07d00001034330f00107000043cc0053000c401c4413cc000c300000cc0050c01dc07c3443c00dc0c003431033304000f0f000f4c301c000531330c4c03400c00054c540cc07d3d4100040f0c000d04010004400cf031c0dc0445000000cf430007700130c0334c000004d0c0704400d3c000000003400c0001410c174d500300c34000c744c04370c3403c0100f31c10f0cd0c400c5c70d0107001304000000;
rom_uints[335] = 8192'h17413c714d1100f0344300c0f0d103c5c01103d00400c300303c0150cc7c0040c0c140030407130c34001403d000d4014101c0534d44c03f0d131cf0fcc1100300c1053405c41113130000c11000f0c510400c1f10ff114043c1dc7c0001d143d0410003111070354111c30040034c53040c041dc447cf50407400c30f00030cfcfc00031171000140fcc04c5cc000034014400100005130dc003010704101443147c03c403f0c303017c000003c0c04cc3040000003007cd41030005400000f5c0301f01001c000030c135c1414fc04041030000310033f4355534043df000c5cc0000d00c00300030c005c0cd74f77001c0100031003f43000003003000311d3c3d004d034704c041c40c4330c1010000350c0400300140d30d00003f0003000033700400d40d0c4400c707144d3430c010fc01700030003c0043dc401031405405770c043f433037c30c0cf03f3c01fdcc0c400c0414d1100510007d01010030c4cf0100030f040d00400c0005004434030313333c3001000c10130004f00000cf1f41044000c1000000c3310c0c4f000401c010010311437c3330031743030d53501d10c07c103c40f040444304d00010d1c4011d4500150340fdd034c5cf0030435330c1400c051c00031c000000330d0013040cf0d00000410000004104410c0c1044c41334dcc13fc01303301f00cf3f55cfdc0c1013c075040403d0d10d04544343c14000030c3003c4000701300013c00303401c005f7c0731dc43c3114c000135010d014070c40005040f00fcc100300d4130304c705301133131c000fcdf33000500000003c730f4c3000011014c0d0d0c43033dc3000710000000d4031c003d503dc41cd0c10cc0000c00030cfc74400140fc413003000c3c10d03030fd000c011403000041c1c01f3154dc74d05044100fc10c14000fc0c000711c0fdf410d54540400c303f70410033514c000d10300cf0d430cdf00304330104c100c7000000404f010c0000c000500c1403004000c5c0340c30307cc03f140f00cf0c1fd300001014f0400000070c0c1dc040c0104441d140c1003cc31300cdc100001100010c0000c440037400c140410430f0c0c37110c330c0d00017005cf3000c00c40000f003130130000000470c70130400000300003115c10340300310d0fc01c3c14113535000d0104d003031d1f3500704f0013c5030c0310c0110000050010100307040f03c50c133100c5040c0f45037010cc040501014cf337f003000c300c3000050031f101044c0400041dc0cc05f0001c0040d7770403310c30c54f31cf50c0303c003433c044000f703cf03004135034300003003313c00535141c1500cc400005000c0f4000131c00fc000100c5400331ccc30d04c0c0003d0c0c04003030300f3041c0071000000000c0070303cc03005cdd0071000;
rom_uints[336] = 8192'h1000000303d3c00100500003000cc01c1000c04170f001d300c31000c0000343c0c30dc3c300004c43400c004f000f50001137c000c0007c100c1003f300f001000d30f400f040dc00050c04c00340004100c00c0c014045c440c4f40fc1c30c4000c300100103440400f7340fc1cc000d000cf0c007c43cc1131cc00007c3010347000f0f40030400c0c3cd0c0030103c004c0000005130753051c0cd4344000171404000c000c43c43004c430000410070fc0005c04c0100c00c034d30000c0f03f0000304f0010014103c4c4f000f44c1031007c00001cc43f001cd4010c10000010304400c000cf0434c0cf0001001544701013003001310c03010400cc0340001043030c050c0001fcc030f1cc33c504041cc4c3003d000010f731003340f0010041010000c343100304fcc00300c00c003f04010004400404fc3c30000cc3010304310300c4000c053704001530301c000cc70c10c1c1c043d1c4c10c00d000cc004fc410c0111f0001050c0000c0043050004044f00f404000c0c500c33fc0104c0000000014004c4f3c10030400010c000045000004cc0000010031cc4f3c0010c000c00c001c3c00c00cc130700033c1401c010c004034c0070d04dc0000f00cd0c040cc0c00001c0070c0350c0c00140f3c034000ff05cc4d0c3101003d04000cc010403004004f7000c00c7044c04d500000c3004040440c434000c01c4c4c101cf40c0c0c07010c43300f0f33015c010000cc0405000c400c05c0fcf3044c0f4000340cc0000010300cf43c4c4110304030044071330400310100040500c0dc00c003f0cc0000d03044d4304c0cc004f340c7053cf0704400c0440c4c0dcfc0cc340530000c3010430c001c10c300340c0cc441c030050c7001500400310cd0c00c0d01400434f0f0100f3005010d00014000411d1040c031c0004c00cc4c1cd0fc14044f1ccc4d7c0c4110ccc017c70005c4c0014cc00000700c70744301004c3010100000c01c403dc04cc0000030044c30330430004344300c00c000c0c0c17c04c304d4c055000400031c300c504c044c301c00410c41cc74404104033c3070c00010c000001c430c0100400c0c4404d40004c07000f14305c70104f41f073010c040001040c404ccc0070400410041f3c0d43000c300c40000cc3000030140413c4130c3c0cd0100031037f0c0cfc400c0c0303c05040040000cc4f00c1000c00410000c007000340103004f43f00103110030040c0000c41ff01000c0c30030500c33440000c0c0f00005430c3000400041000fd0400c71cccc43c41101000c5000c45040034c000400c0c70005f000000c00013404010c030cf1f0c10c040003040150c400c01074000403400403d40000045c40c0000310004c40f1501c00c000f0003000013500304010c1c3034001d00040dc0400;
rom_uints[337] = 8192'h3004c030155500330004030cc70011100500550003400511000c01003f4f0f4c00030c131cc703c005cf0c00c0007704103303010dc0f03dc000d4cf0c0f0dc031053c0300300505000000000d00c00c04401d44cc0c703c4f0c017c0c01d04004c4400f000f00c100cd10000100003f3407050cc4004053040d4001c110cc004d0cd300044c0003c037c0047d0000307004000000004300450c14074d531140c1450f044400c00c300000074d3100737c4fc001000f0003005300f04c3ccd33444703c30100f074c0c000031c05c035303f000f4350000c00134d030f3000d054040005c3cd1c00000c04313343c3c10300c1330fc3000004000c0cc30000c073140c3c00cd0304f13130d5f4300304ff10c0fc000510030c1d1d47034434c00c4c0000100347410c71c00033ff014cdc030ccc330d0104c0033d0c03501c03003fc00704000100dc0c00cc3f01c1c33fc300f004015dd0303c010110c43003000c43300001c3cc00d01414ccfd100c0c4300040f40410c1404cd00410004c504d31500751573043c40014d4c40fd131d0001070100c34144000d0c4004100000030010d10f301d3007cf00f17500000410c00c074000000340340c30004c44100cf3cf4c0301fd0045cc33d033030405000700c34f030404c00c13000c4df0d00f44c4f4103f0c03c475c35ffc0301f0333014330100c41d0403003771004150c34c11dc0c00300301f3130740c00c400ccc30033441000001c5c401055cc40305303333135443000040000407c0300443cc03040000300330cc0d0c00004c0043c00c000004000c000f003cd4f3d0c30341000107c5c000300f017f0700033411000fcd0ccc40440414303c00030c3f0f07c541cf0d0dc003cf030001c10000000cc3f0c033400000030c0c0003007d03043ff310c1c130100c00fcfc33100000f30040101071307011c4010401c3d05c0100cdc13dfdc10c4154031530030f3531300f0000004300003001141c1731c4d000d0341d03440f0c0c304131cc43003c00301430c00414f103033304c3ff300103000f00330041010340c30f000001014714070543030010c0400cd430030c000fc000dc1000c0c00cdc04040c03cd000030c70103c00033040704f003000073dd0d330f340c10cf55c0f40300c007043300004510014304001cc4004340d1c10cc0710d050103000031043f1445003fcf714100cd11731c103fc0714cd70303c4c3000403f04c443c004001c5c10c01c434001fcf0700304d00071d0c410c0103c0c00100403403c01d0c0f7041004300c110101c3c40010c0000011400f00033cd0000f34401c000c0010c03004033cf00c010000100c305c003c000003c0400030300370c0071c744000c30031d0f000404c0f01c04001f4000fc004000000c000cf3c3004f00c5040f0100;
rom_uints[338] = 8192'h3444000c000c0c001c00001c0f001c0010c3030c30003530003c4334033003040037750cd40c070d0d1500000300cc0f4c540175d45000103c00000cdc0000040001d704447050313c001f04f70f3cc30504100cd330010014000d070c4f0d0c1d54171043001cc0f44703014350000001043100013733c0c0c0010000100c30c703441000430000304300000f10000fc04c044c00003c1c0f033f01f701000003340c010000030700cc0c00033c304030c7ff1c00043c11413704d14d0100d01c44000c0c04030f01030004400113040004000007cc00003001000144d704030441000003100010000c0c0f0003400010304c00c0000000400040cf0c00000c000000ccc0331f03003f03031d0441000ff30c0c550100041c31003404100c11000f0000300444001330003405f103c30004400000010300c010000350440c0d40303c4001001f040000004300c401300030030f44c75500f1f31f341d003c0000073000014c000014004c1000c00100cc01000c1105073c100c370fc50d10003f140700004c4f03c35c00003000c3500c003003cc00403050f107100d0701031c45f100d00400130f03300c03001f00c10c101d4031143c0001d10f000f3400c400c41103140c3304051000c1c0000dd010000c0100301d0031011010cc310f4134003140c10104330c0401540530040003c3174c17000303c00030311077170530170c10f0030d0c030f00010010430d07c11cc500000c1f313c01f31cd71f0070cf10137500c00140d010100501000301d0000013003317040000cf1c0110075c0c070011cd005c0c0033070411c4013dd001104f010300c4c0053c003d00411f300f1011030d311c00f03300c00100413c1c040d0dd4c0001c050001c113303c0000340010000373f30135441d00100044010c0f0310400711001c1c01cc3c0304000000c0313000074010005c00003103d4030034000c000f1f374c00000040c000000053000407070c000144000403014c40010101d71c330303f3001c0000001303c3c40001043f000000007d4f0004011c400c00110415030400730000c00c10104300040004040c34c3001dc14c430010cc440300c3000300010c0131c70000ccc0000c10dd0000c000334c400f3440f0c3c344000c00004300000c7f0c0333030001054035401c1f0c4c0dc70000030dc10c1c000c04001f30c174c07c100011000000770f0000403000c00304033c7000f1c40f0300000314010cc401c0c057001d403c00070f700405fc07340030174c033074011171c3c304005fc0c5445c131d7400f0000c00c00ff40cd031cc04007c0003404d00005fc00304c004730c4dc704c310310c00cc030c34010001003000001133070cc53310140140040cc34034004cc300100cc00134334c070005c0c30cc01d401700150c0c;
rom_uints[339] = 8192'hf00700c103010043000040c030c143f5430001304f015c1070f4f3334f0000013fd050050300c1c0d00440400c1007045000031430c017003100c0f0dfd010410d10001d301100000d05330100cc1013133f11000103c3004f0cc300f453010010041301000c00cc100303c4030cc0000433511c0c1cd0c340cd1000004f0330d01c0140000ffd030003c001101c00f50001000c001000d00f10040f410004010c70010000010c400100000f0c1373404c10c00d03001401c00c0d0000403c010011005000117100c040fc1c13c3c000c00d331100043001c0300c31c31d501d40010c1c03305c0f40cf5cc073003f00c443fc0cd04010000c400000c1000f310310400030100d0c30350017f1c431034c4c104103c0750303dd10004000fc3cc04001431c0330000d0d0c471440c3c0003c00700000010000300d3d0031400cf1000dfd10100000c011c33300010fcf01010305001401c104450501413000030f00c0f033400c040540030034cc700000110c704310f1c00433037000fd1cf1f30540c53100c70010003dc30f0c3c0003000310110011c0300cc000004000043400011000013f1043001004cc03400c070c35d0010cfd00103140c00f54011013300013044cdc0f1440034003010354311c00400301c000344404001000113030c1114dc03300134c1ccd104c0000cf40450044030405000cc100c33f01c0f10f510000047d00030301c0f300000c1143f0c0301f3330d17047d7c734030043004303c0f131300100c014001c101f4cd1cc04350c3010134070444033c3001ccf01040c000000030300433c10030f3d5c0c0c3d04c104d0f403170f41300f0000100005044f1cc003c0404001c00f003011003dc0c3000d3100c1004003f00303070f4000031c430300c0c130010f1000004cc34003000d070014434131304350c105c31503f70cc50f00cc003417c13474300ccfcdc543444c1cf07c3304c00110000004030333c3013000c030d0c00000074330011c1f13704c31304013c001cf0f000c0000c0c030fc3cc013030c11f444dc01430001010010c400c0043300031d500143534101004030004010d0010f43004300c00cc1730100050f0f0ff00f0c3113331d3053410000153c003c1340f0c01c000f04c0014000003400000510c033000000034501f100001003110c50731f3c0f3730c03c0370c0014ff50c000004400c10403000000403333fc4100cc1400c00433cf100c703003003c000503c0000300dc1030f30040f00d00011cc103011300131413000c0400004f040d134f011104030000c0100c0010007cd041303030f405003000003004300303f10050c0f0000c04000100c310440c0c0000400303300007cc00041511d101c030003401000340c30c0d403074c1f05c0c3c05011f31100014400000c000;
rom_uints[340] = 8192'hc433003c01107d00110030c333403cc14f0000100030c1f00c7030430f40cc04103077c33c7040030f1d003014c0d01c330000f3043000400f0031000f30040010d00173037cc0043100cfc0300010c4c0c100503410d400010401c0503c30401c3c74317303003400c3410015ccf01c130cf00000d170005001c1c41510100000f401c03073f030033030304004304400c0300000c043c733d03033d0103dc4f40c000001fd74fc7cc070030101d340403f311100c0000cc17400c4c0cc4c034c71f03044007010131f1c3c31d5d0030374f00000300300050010f04410c40cc03400f1d414d033f04dc0700ffc440004c0700c33040004cc030030fcc000c04c04141004041015c01114000003cd330c3f4d10f051700c14030051c0000f00c00107000d100c14f500c30000c404043fcc300330050c10fc00cc0004000c0504503434d033c000f7100c0c70037700000003543c1130701f44000100cd51044400704c737f1cc0d50501f43301000c0400c010d330101c003f10010000dc507cc0700303f00c00700103000430030104001000f00001d00440100050d00000f1710140f7c0104300c003711003f03150130c40cd0030d33c103c70c010474dd0700f0c3300007014300f00331030335000300c003c7334c010340703c010d3403011d5c5c0500100f5003000cc3013d100330f0cc307c310000400d304cc073034f033040c45c000c77c000cc0c0033501311cff00103003c13f331313440c4430711c30f5003c0000cc50d30000041400c341703000170007c010144c300f131c131000f0500000c0cc744340c0c300051cc0000430d3d1f700403f010c30000010cc1704040c0cf00ccd000400d00310cfc44fcc05101d04c100d1fc334750443101003f30c00037100100300430c300dcd133f50cc400cc040347303f011050303c74c373054134344c7c0000cc007140041033d01c0000731001104400fc3c10434000030030f04313010f0c3000303000c553157010300010f04513000000033173400100c13004100050011c5c10f0fc0f00301cc01cf40007d47013cd001004c40c7530f10100d10000c433f303c0d01f7010000047104430101505f100000030330030c11031050004005c41073330300310000130003000300fcc5f00c140040c00f140304343fcf00fc00034f400011100113ccc7c304c7333031440100cc5000304f4500c0dc40003c00000331c1444f04030c40034503001044cc0350c40010f0c00005f14147130f540040f0c3cccc0007440c030c01030403cd40df4030033c150d1c100040304000553d00040003c004c1001000370300c03dc103cc03403f10001fd10700d034c00107c0cc04100f4c4f01031001530d0d00c0410c00010ff401033000113c13d11c43cc0c0510054d01400ff00041000;
rom_uints[341] = 8192'hf4cdf301040040f10fc01030f31004ccc00401040001c4c013c7141143004d0007c30110307000043030001c000fc01300034f1d1054c4334401c403313070300cf0ffc7043d44044000d0c0410003330400011d00c04c00c0030031001137c500c3100050100043010c030401f111c1400340457f5c004d01007011c01150c000000001041103000cc0cf40011003010400411000000c040c00d300303c1011000c4c0055f03fc403031305400003310000300000c00301f005007c0cf003001143301314030371103000014000cf41c3c335c0c345c0300013115d7003010c500000d1010f0330c0c0001c4c0f003010400f50150030000c0001030f0040c0114303017c0f0c0437104043000d004003707000c0f011c1455100003301f3c0004c03000f1f01c01c7330f1c30443710033d010c001030073400d103005c040c10c4dc700c1310c0300c1005c0c13330c000373000405044310040000cf37cc30d151d0cc170c0c404737c0040cf0c30cc10307000c03d0101100040d00c0d4cc1cd73c00013330304d0f50710500c00000310f4000030045040304000d37000015130417c753c3100cd34030c4730303000133f001c710cd51000c010d005d0d000f437f030c3f0c1d03c0030030c071000303330d43105043000c10400000003013cf00c54103307334cc013cc000c31370cc330100435003001005010d050110c10d0430c43c040cd33c0041c71314d50500d000f117f37cfc303df030f04c445f1540d00030000f0400c040400300c4003000170c40010d530070000115c40140c0d0cc5010c0c05003040400330000c1000c07c5000c0013d04c01f0d1101010070403c075044410c00000430000c0cc4f40c014d0c0304cf10030c757001c100c43174005c30c35c504c0001341001400c3100004004310073700d0403c73d04f07443fd0011015f3dc00d1004475c01311070cc04f001304c3c01311cc0403030000c010010310100300300410331400c0513cc5d4c04c40034c0c40d000c30c0000000f0314033c0000000104300c44031004030010540011400000034c000c13d71370400100f03c01040000040001c043c00030070c4700000700300d00f04c03c0000f4003410c4303440000311103c341c0c31473550d00010c3004c044c0c3c40500d1070013430474100c100d1000003107001d0ccd3313c00c00003010100003d05000005100cc011000cc34030dfcd0cc40001030011c30ff01043c100137c037000004cc0c0df011040000d70c40f304504c0471405040d001f00503c01703003cd040110300100003c00cfc00310f0330300077443c0fc31c33500333df37f000f000443cc0001400100000030151c00000170fc301c4f4c044304cd030d300f3054c444100431100000000000040433000d300000001;
rom_uints[342] = 8192'hffc74310fcfc0400c005f1500c000010c00ccc30c340ff00c0d00c04143401f0cffcf7c0005d10405d7000c4cdf03dc00f1c0cf745d000503040c0100000c054700c51144d3400c3d000013004003c5d004104fc7710110c010c00510cf11dc050310700c444304103013c00003734d75ccfcc405cf0d44000c4c0007fc0c440c330ccc0c0f4005c00d4000033c043c00311001000c0c040fc00c0003007f00c41f054f1f3010ccc01000400f1f0000031040c0000c0ff0c0cc3004cf750034104007c4003f03c30c0000030c000415100403000c00c40cfc4ccc03044c40000ccdf0030f04300003443007c404000c0700c4c4cc4130040c0f004c0c44c0010340c0cf00f0c4c3010c0c00cc10003c3cf3c500c003030040d500c0433033010004cc000c0f400c01c10cfc035345d40c01017c31434c00000c43730d14d5c500c374c30100731030fc4c0dcd3c0ccc0000c041cf05c31fc4c07c4cd01000c0f003404344cc4340c000cc04ccc00c0300003000c40400c105cfc4f0c7cccf001c0c071c1d01dd00f4071c0f0cc00000c0f0045004d0c4c001c035c5c0740000001350c3f5d0c1c05c0001c10cc347d43005c3300c1015003f0310cd4740044430f0143031433014000753c007d00400030cc001c0c40c4400000f0c030044c00dcf03f701dc0040010003c0070c4f3004400c030c40c400400004000c030fd0cf000450c0100c01c703cc030001110d3f7f44cf0c00000c0c100f1d134300c0004f0007cf4d400d3001c4c0071013300c74c0d00000050c10104014040000c3303030150f0c1073040c044d004f7004000c044c004005c00400044304c00c004cc00000dc05ccdf300300050c00050c073fcf0d034d00c341501d00000004004c3143df014303301c0004cf3ff30c010745003f03410cc44c0cc010d1f30f4000cc0030030cd00c404cdf0cc74c0040500f00400401500001c0010fc04c0044301400f10000070000740c0c4000c30000050ccc33c40430c0c0030c00330cc00300040403c0330000cfc0000f5300044c00dc1c00c07010045cc5d003014c400cc000c404501f03310cc0cf003c4014171ccc000540000700c4c10000c5cc050300d0000f33000000c300000003c01d0040f34c00110c0c04c000f1450700400c00001400040cdf000c40cc4c44ccc11f4c051c4f0c300001d73f4c007c04c0000f314304031c00cf510000c040141c40000c04cddcc000000010c14c0313c404300cf03c4400040c0c1030f4034c0c0c4cfc0f33c115ff3c00c5c0c0c1014d4040d400cc5f40dc0d000f004c010c00003cdc00047000073050dd0001f143cc000c0f0d0c4ccc34f040030003400f000000103504010c0150cc474c0500c40501c03307cc3c0c0cc00d041404054f100070000500c7003105f0c51310000cc00;
rom_uints[343] = 8192'h34c30d0f14001000f31010001c3c151cdc00300400f3f0070015310011c03103040c0f0010d00073000703c334c0030c300000c004c00000000000015103040c0f04c75f00000c0cd0000010f140013d0310000405c103003404340c40c00f0d333011541c0000001f30f00c0c050c100cc0000c00c00101000434c7c41c00c00443c0041300000000100004300300303d4c000000130000c43010314000011300c4000f003f0004df30100c040004170c450010001533f0011001f7cf3d00140310530000101d01c00c011140d43c000304400000cc033c000c0400d5400ccc14f4000530013030000c0033c00cc400003c00100c330000000000cc000000400004430134001ccc30004404c00c000c0ff0301d003000154400001d04043c04007001004d000cc0c00c4010300003c370100000d30330004410000013d000c00303340400c00d00000401310100004c000c00c01534044431040735300cdfcf0304c1113c000c0000f30103310100000400c10000003104401c350000740dc004111c0d00340040054000040700350f04c00c10700000004000113c0700010044030c30475030000c0c110004f41400c00410404401003c04043c043414c530003000001c00030100300000444c0103c0f003004001d1033030000300050004001434d3d300403530d0040003410100303050034041411004473004cc00c13400040401c30d03f30003cc1c0c410000014034100100150f103c010d40310f040300f3014d0f0c0000040004d0033000c3dc01000103c000300f31c304000007c00d00c0003400000001470310000c013030003033333000001010110c034c1fcf0000401430004000010c0f03040130014040f1000c04103c000001010005c00cc000000104300c010100f00c13c14005031c0000000134000d0000c71314300ccc01111c704c000d03c03007c00c5df03410c730430010c000c3001c0010c4400000d030000f00f04d00000c000103c0510c01010f00000c0001000103cc001f001d0017000d000003003000f00000100343d3304c0c30d7040400c015cc10310000337300c001100000cc4001040f400035041c00310c007000d430000000c310000f1030400031c400114034300000f43c30403c1ccc00053d1310430c7c00044c04037337044c03010050f73440140f001c0f000c030001d000000d33074400017307070030d40c050031000010000cc0cc030000333c3f00c3c004c07310040400d1000f0c0040c007cc14cc0330300034c54cc3001313c00030000110cc044033400744010d0d0403040d04c10040c740100000c000010000000131404711343c00301c3000003430044017030c0430c003fd000307d500100c01000000c500000d000513340c03030c003c0cd30041010c4dc7c01c04001400300000;
rom_uints[344] = 8192'h1330033000033c0500400410133130003f1000cc100001000341300000040c40003c300d003d00dc000100011c30303cff1dc000000c30d000304043300030003004c44100000c01c0007004cd004303500040000031301001010c7310f40c30153030000f3001033007c405f3043d04014440c500c000330030010014c0040010c4c00c101000050040004330010100100c000c000c010d013c3d703344433107f40003300054001000001000fcf33c3103730000040130000c04400d0000303000003f3000330000000033c4000700330100003073310300300403040313000340000010131110043000f003400000413c0f13100c00005d0010100c00003cc003401c0000003400100c34fc31000c0304001001c03000df01013cf43317000c04d000047000c43000d0040410403011443003040040000040003c3300c00c3000101400f03c03d03d730001403000d44f00c0030110cc04100f170000030000300304104c07010d000d00331000040134001c7101f43010f003301011cc000033000c4f4c0c10040c30000c00043f0010cc40000014c40c0c0030f07300033c00731c054000c040cc0030000030c103fc0107051704003c3010000000c0d00401300000700003373000000403100000c00010100000d3400030c1c03000001000730c00d100100f0410000000000501000010100c000c00430303030034033f30000c330c00403103433403000c30cc0c100c0010040340c0c30000000074000010000000d03f000030000000303003000300003030d4c0c033cf0f0050100037f0100431004c030c401c04011003c01c00040010300034171434c00c0130f001301c00301013000000003c01003000c1000d00030c7410345c1c33c1cc030033f433430410034ccc130413010c0103037c0c30ff031000cc0d000c30300010d7340337000111043030d33300330d30010004140103010d00053c30cc30030040030400000004c034300034c0d0430400f00c3010100d33000040013343c000007000cc3304500000303030c4140300070134003d0d1000d00400c1103c3043000500cc1430c000000030000c301000000c3c4010c0300430400353f0101400330c0133d0333304c00000303001000004003000000030047c00c003000000311c130000c10030cf0004303c03110000700343130c3c3344701100c0371f000130041400c00000004304100c0c0000001030500033013030000014100c00141454305137000100130d3437103343fcf00f0003034c000014104c003c0011100c0403001c0071100003331c0143d0300050430fc0410043371130000300040c1400004f3c1cff00430404000003000c000f00000000443300c3c443001330c003c4040c00d114700073300040c310101c000400c01000c7003d01440f01001c;
rom_uints[345] = 8192'h4000030c1003000010000437d010c001f3c000340c4fc30030ccf310470f01413c0ccc0041d0d0141014404c1040c00330d0703cf41005330001d0c3400073744000404140c50c0000033000000000c000003c4d31cdc30f403003330011df001030cc0130034000000d001303c000100300c00000310300004c1f4c5c10010013403331c4500300c0303040000443d303c400100d03030ff30301043301d13304350000000000303400f1317f1c0000000070000003030cd000c4404fd0003044c34c300041043d0000005050100371c00c00cc014404401410044334c0400000000343000df40c0010700d0730c400d3d3c040000000000040c43400100d1c0030300071033035c00000c33010c15010c10dc000031304300000dc0c00f1704400300c00300cc431503c13407d1373c000000040c0c004c400100001300c4d7140010f1dc07000403001c30400c003003001d3010040c1c3c0410000c1c0c3410740054004147c4d00cf00f00301140001000f700cc0000c0c00034713c03500cc00014000300100403000703300c0c000701000000003c0c0010c40c003c4fc00110f003040c075c3000c334370c00000040cd3c04013f033003003730003c00c0114f4f03dccf141000400c00104c3001040404735000301700d731030c0000c30d00f7013c3003003004000334000040ff40004010d40c30010300331ddcc0c000c013c3303144004100050c4f03130c00c400100700343c01c00114f447305c0c4700004010070410c407351040000500c0c303000100007000400500130c0000003030403c7c14c700030c00000100040000150c10d000300734d101c03f0c30d01000c400cd034d0c0001c00001705c0f1000041d0c410003000f1733f0730141c33104030cf310031dd3000347df300000cdc000df041413400101101c00041c1003370c1d4c53030c005dc030100f100000d0403070030701c033311003040c0000300400030001140010004c004c300004000f04300003f130001f001300111c004101031030003c0c300003c0443cf00001000010044351cc401c0000051d0c0c004410003d3430d4cd00001c1f0dc00c03d400500f00330c000c0400c1f1070400300000304c00c110300030000030d110013010c13c04444011001cc04100c0000004cc00100013010434140004551401c1003130705f0010300d3c31d00300000f0430000c0143014f01000c01434df0013403030003c03000010343070010004004003373053000c307000c00014001f0043100073000403c131cf41310041030001011000c0403000400031440310000030300cc4c30030000030100c1030030133300c35400101000030004000030000c010c00000010003c1104730f0c10004dcc401c043707400c0c0017314c101cc503cc0c043001;
rom_uints[346] = 8192'h71c4c0004057f105510040d00404c010c003c004000430d00c3070003c7000d040100ff0c115000340c300d4434001f070c3001030750430f00030c13d31c0000040000400c0044c30000000c400515c1300c53534301000ccdfc00d4f34101043440500700010000c13f4403fc10307401103044310005000017cc030433105305c10cc0037405110c301f13000c050003c403300037030353043104cc3fc0000004044044140344500f411003f40f300513dc300105031cf10c0710003010004d101014000005400d51c35f300011330100d50004c3c3000130300d5f310f404103000504103004004c770c01711040003f00003c3000030000010c1f010c370404dcc45000330c0003c4400f504003ccc50000333fc1301d000150140cc000c4500005304440700730043301300f0f3c0007101cc0100c03003404400040013000041c001c000310004033c00cc00d000471431c300404c340400771004703410440000d0557cc0307440c07cd03010c0c44300034c500013c04403300c00c01131c0ff0010c0050470003c40d00000000c010cc000000ccf440c0000d010f07cdcc0c301305300d0713c4c0001f00000d071130000000045cc00000104d0c3401000f0010041000510700c00c004cc07033000d031c04001c013d4ccc00c000031710cc3df3c4cf03030c0cc410000403ddc03c0c030dc0410005f00104104c000dc00100000c04cf10010d00c1040530031dc0400d340dfd1c5fc00c03550303014c4c350003c00c0405501030c40c4131004c05c04001f01033100c0dc33f0c0000500003504c0010003ff00003041c4d0015004107041c000110040c0d0104130410fc031cc1d3c04130140033310f1c05031c0c10054330010d30c1000011c35313044fc141010c00c300dcfd503c330d1134ccc0041130c1171330370110c41400fd3c0c0704c30cc1034c330c301700f30c001f304c3114007301c000d4300c0004400d70cc0d300cc1c0004d4fcff30f0300344350c4011044040100000c073cc000000400170405333ffc0003c403c3010000c1310041fc3dc0400007330c403007cc11013c0303310f0d0d00010f3d0df1300c040c130c304ff1030005f75c0c135000f100000054043005c0f00f003400004c3c030c03dd00c3035f010cf000cd1c0375014c770d31c307c00cf7007000c1c74043cd00500c33500cf0340000000170310041c41000030135f44411c01d0040140c30ccc34704053cc3434004103cc000010d00414fcc00c101c00f00011404dc0c001f300c0040c04104100500cc0340441d0c0c43c01115035c1c00000d00c1000d034cc0054444c00453c43ccc301035000001010fc0007c340407110d001040010c3004c000c401005001cd3003701004101df01fcccc00010103c410151030033fc3400;
rom_uints[347] = 8192'hc703c0040404704047c00c300000cf55cc77004030c4f30104c00000cd0000000040000004c1cc00000c070f40000f03034c03f045f00c4c10070333c30cc0c0cccfcc1c003340f43000013fc007c00c00c300403f0f0cc33c000c0f00f0000001340700504ccc100d03fc010103c0440d50033001c04f0100c00430c000000c3f000c03cc0004034010000000010c0c00100f00001004003341074c1d4100001cfc0c1017c017340fc007001c0f3000015cc300000c1101700000df40000437c43300c40403400c04d0000fc003c0d0000c00000d107c000000c000fc4c1f0c3c000c5c0c000c0045c00c140f01c000cf040c035fc00c040c00004750000040d0300040cf010100d40001cf040c401004c00f004c33c30000c0c401f301007000d0000d4550103c1c00010401000cc40c40f3c41c41000c000100041c00031fd000000005c3c4cc30004cc354040c00c0100c0400cf04053730003000143333cf0c007307000c0c00040004000010000c0c340041d0040400c034000c0cc0007007414000dc5011cf11000c000c030c000c140c0c01005f0c000304040d0c0f33151c0040100c430017000f000ccc00c0cc0cc171f0c1000c0044ccdcfd01c070c4c0010403454003d0c0c54000ccc000000044000c000003000c00fc0000001fc7c33050c01070033d0c0cc13105c3cc0c00d003440d1c040cc00703c0053700c3033cc0c031500f170f0704000c030001cc044000c0404cccc300110fcc1007050c104f00001c00ccd00430400700c3cd04000404c041c0000c001000c0000d0cd5040c04c00030c000c03d0c4400000300030c040141f04044d01ccf35030c000c4c00710fd0004014df0044c4040c04101003331430000c000dd3fc340004c0c43010400d010404cd00f43dc40c1cd101000f40c004000c30430cc731000cc00000000105013473701300c0c30000c400014c000ccdc007073dc0503001004c00100000040001c0050001010c000004c041000c0c03300c00000440000c0004300c000430400f0c01cc00040cd00dd0400430000500303c03011040110400cc030011000c00c00400000001c70c1c0c0c04044d3000000cc4f13307013f0fc000c0c0c003030f0010004041c300c03000c0c130004004c1000fd00f0000000c0c0c00c00c03000c3c04410c040010dc00c0000300cc040030c004c07c000401cc0000004c140004001c07074c0004cff4000fd4c400c000000003003cd50c0003440003300003000c004400000000c10c43000dd00300000c1ccc4000001df10c030c430c40003404100030cc0004400f04f00c05110d3c10000001011c400c40040cc0dfc0303044044410c5cf4f010c0301c0401c04c007c17000fc0c0c004005c0317c3000c30c00300d4503c0400c0c0d0000c0430104334c000c0;
rom_uints[348] = 8192'h10d00f001c00110000010000100104304d0010f70000034c300d00000c37c0000000305c404d00300700330d000003c0010000030401031341040030000000003f04030c043000cd000010000004041300c00dc00c0c104004401c1034000010d401500100003310c303530c000d03c11040400f040310f0007cc1f01340d00fc34330000000043000fd00300000004000010000000d304cdc00000d34000413003700c0315350100004001000c707c3000070010003343d1400000c0710303c3004001d10c0501c300c04c4330170030c04c00030140300d4370037c3f10c0030010003344400003c1c3c53331c7c0010143c1c03140030000010003101104f0f0dc0070d004c0044cd0070375c000d303303d003c710004d1c00434c0530010f103000771010715400300004031c07010314300d00000c300cc03c14103c400433000001001c3005f00030c1c0003044c300410d53cc700300cc5c0401030311031000071d3c03531400001c41340f7c4c00050000d00c1054030cc0001400c011f00d1034400d5d0000013f0073000c0003010000dc7304001cdc00cd030d4d1c14d000030330004c0c00440007c30430017404c3431030c000050cc00f0c01030c01c00c400000100c0000015004d300053334070c1c14c1030d0007103001c00d401000717c0c10c0000400000c43000001040051010301401000044310004013000c3014031d310c350014dc1407403d040fdf14001c700d4d311d4731000100001d044c1000000c0c0d03003301f00100011004140c070c00100000c0c0007d001c03001c000d000c30300c403004d00011050f1f0700040070c7f51f7304300c3fc70304c40dd100040400003030cc4c1c1100003c04000c413fd00c0004c40d000334f30c4301c0c3c03d004034c70f00000d1300400c40000dc0034c03c00030400004170333433404134f0c300dff07000004044c0010130000000cdc37c000001c017c00300104f040c4004c01000cdc303017300f0c4100000070001c0ccf4d03c0000731000400000300030c071dd004000004000135131000113030000fc4f0300004033c00c34001340400073c000c0c00c0310001000103341000034430010c10f05141040dc004007037114371cc1001117000000130310f010d041300177000c034dd34073f70300c0003340c4c00d30c30000033000d1d5d00001f1c004000c40001c000001d001403001004311c3c1304031004cc417cc4330f10001f00f14d0035004d000c00c3110304103000c30c103443cc0000140000137d14034c0c301c1c03000001000d400d0c0c0403341c040030d13f0330c7c703000770043c0330017c3000000000000c00000144001ccc1dc4141044004c140410f40c3cf0c710330dcc0303d350101d40304000c01d041c00030000;
rom_uints[349] = 8192'h3304c000044300010004303f4000c700000d01c05300c31cc3304d04c40c34030043c40f404407405f00000f00c1d30c3f0d0501000400cc430440031c0000c0c3430c400040cc030000c00004c0c0c0cc000500cfc3cc430043c3cfc034000c00404dc0c100cc00001dc3c0000dc005cc0f43f00041000f451c0f3404500003c31ccf110c1d004400070c0500107007005343010000000005001c301d014d0d4000000f00d000004140400c03410c14c0010005000cd1000dd10107400000c134700c4f30034c040c0400c50103010f040f00030000cc00030c01030431c303000300cd0040044c04c70101070003000103cf1305130003434f0001f00004130503c301f4430f4cf1c543400fc0004c31404d3501400c0cc10c04000ff40301c4053100ccd300c10f1d0004cd003400c000c403340000000000043005d4014004f344040dff40007001000100c3430d000fc744c03c4043f01c0530400f04104cc10333c3cd0110053c434300c40d040c4f000c0004f403400fc3044d0d0cc35301070cc04f4740c4c400004c040c1f0d0011f01c0dc00c53c00411010c1f0c53055c004cc00300c0130300140c300000504101c1c100c30c0000430113350100cf000d03f0000c00f3ccccfc034000033000cdc00007050000000f0cc14c3d4c0c000c4001010cc1070c00c00c0304c1070040000300c00f0043cc3f440c4704430c1011034f410313c00fc04f0000ccc44c41cf004304c04c0c444007004004004d4c304f001000000004cf0300c304c1c100004c01054f0407d00400fcc0454000c0c30103030c300140c4c0410300000f0000400f010f3000300c1c44fc03033001530c1d011c303c00c10c33c0cc0c03c0400305050047110030034fc4cf744c3003c0000cc40fccc4c10300dcc33300c003cd0c30000ccd00000007010d340741f7001c04cf3030c000f3ccc101013700001101c3030101330150c73f00000f0400000403c303c14000004c00c34040500c440dcf00000d0cc305c00c0000c747c403c000c04df03c0003030cf4cd010f0c0d0000c30300030040f000fc033fcc00000043c74043c100107c00cd10400c00004c0c447443003301f4cccd450000413004001d05340c10030f0c00000c00d1cc040301c5000440440000c030434300f7430c0d0c0f71f103730cc04c000d0041150101f4044c0103c040354f035d00440105400500434f000041c10c0f000000431f00d100c700044040c0000d05c400000001003401c0c000133100c1f03351c5001033004cc0dd0c030d44c04c4304704d0400c3054c07403300440cc330000c00074f0c000440dcc0c31c0fc33000c04c000c7d30c300c340c30d0300000003030d003403030303c30000040c3f0c4cdf01030c0030450d00c1000304040c0c333f3f4c0301410100;
rom_uints[350] = 8192'hc10043004040040dd030004043c3340500000041d70dcfc00010000030c00104441344000c0d000003710004c003010f5dc5c0030015003401dc04003140c0404400c030000300000400c335c0000447000c0d40f501c0c34010300330c7d000c00cc30c4004c1441401f00370c000ccc0c113c304004440017003d10000c070c344000004c130d000c430100003443fc00000000000004340400000033000104400fc0003034000c0c00001330001c70011450000010001c53300cd050000315003000440044c03c04100004404340004c04f0000d4040004f0c300f3fd0000c0c1034100c003400034c03dc0d401f14c00c41710cc0070c10740c1c1c0c043c0c0030003000c000cd0031d0c0004000170c1c005041400704000750c0c03c000c340003140c000000f00030cc0c3041cc5cc00d074c0000d00334c44c00cc17301044000003100dd0c0d00c31103010d4f00000000430f3300030fc0c1401c4170c003cf100dc0cc044310c04c44c0c0c14100c00140000403434040003444c0c144f1d0c000000c00040314c43c000d0040c44000df401000000000400cc00c0700030140c04f40300315400c0c000c00100c35c0cc030340c00c00f003c0010000c000040471f040c300410340cc400c05001101430c001004100010004403040071000000d34001034c00010c4000010d0400000043000c00000c000400471403cc000003040043400c030134300d0000010030011330c1414c4340440400410004cc0d000300c00001300000370fcf00000c073000001034004ccc003fd00c001004c00440030f0003303000700141c000c100040000130040c0c11c04000c07030100013540304f0004000000040000c100301400c000d0014cf0744400ccc10430040000c030010004340c047fd1c00d440c0c40000000c0fc03c015013004040453c10300c0003c1c00004030000037410040303441030c0c04004010004cc000007000304000c04445340700c100d00043f0734cdd31c0ccc30c000300f000373007c00043010050c30300047410d403d000c130401003cc003000c1004f500001003fc040040c000c040004400d33c0c0014000c30103004070100031004000000003c1dc0000c300004000000c10000301c1004005040414c10305007103000c0c0041c4003330015000700443cd44cc03cc1400050100430041100400400447004113c000000d40c3d1cfc0cd0cdc00410004d440100100c1430104d4c000000f00000003cdc340c03c000400453300cf00c30707040f00c400030040d0003013350001000100000c000031cc70fd0005c100411000013000010000d005000103f040030c4344f000000031030000c0c1c401313c440003000031f1044dc04141c310cc000000c10140370133fc000001003c33330404100000;
rom_uints[351] = 8192'hd00d0000d405100373041c01001000100007110113dc3071c01f44340d101300f03c470430040033c031c4447100d44c0370d013150700344c03003cc03003010c10043401170504d500c75003003000073c0f10fc31c1043c31340c140331c1000f0c0f30004fc11000373004cc3053050030000c1df4d0000d3710c00573c30030304000103401044cf103130000030d0c003400c04000d00c70c00c00710030c3030701d03c3510130004d00400100c0d0c1000133f3c47070014dc303001035001fc3400f1000303001c3c0031c1d1317450010c0030033703001fd304fc0c370004043134314f1400144ddc4314110034d000cd0c31d0700000c300000dd3330110df3c13104013070100c3330f70c3300330130c0051040010c05ccfc0030ff0005f41ccf003ffc0103030fdf0cc41400c040470c00073d4f013113c100003131313c0d400034c0c4040c031005f3c00131ff101cc305407c333c77cf0c03d0310303400d01140371d3103730300334c0450c401300010c73d00401001c743000750100c00fd1f3105373c333d31001500cc3f150104010001071d003034c0c53004c000317004c3101004fc404c0c4f3353130440cf1c041cf0007c43405333c04c04047300313f00f04035c0d5f0400c0f3343f7000303313c4f004373101034f1335300407c13300d070c3c31001745430030fdd0d300100433031c403100133d4f0dcc00cf0f0073cc343c003dfc14cc43c3347031733f07cc044f3c11fc40c0cd11300000c104353c00300c33d00c113134d00110c0040300d35000104f0c0300040c3c043c34d4c400040cf315000130fd710001004c410c33c43f000000300530d047c0010c7d00030cc0c4df3310730001c31070c00c303501000d10043cf0001110c4d40f00d405c0cdcc3d037c07373400f0330d0c3c1000f3400d004cc1fd50d0c00d3740531001033f110040340103ff0d11110d140110c00400040100c00c003d0003c030d4040c0034713cd0c0044ddf533334df5330f000fc03d4370c7400353d3d0c0003001f3ff403f100100c0144110430000031c7cf140107300c3c0f0c047300133000414c3000fcc0043c0300040f333d043073c000fc01ff0c3d01001f4c1000040403c0d07330011005fc313fc0000c340cf30c00c105cc0301c0c344f000004cc03c31010443ddc01c0dc010001700350404171430c4140030001000ff4400071c03000f00c43d7f113014000fc101d50c3f034010000cfc3cf3000c0c050100c030c000cffd71003014041000c003013334004c0501003dd4131f173707400335000d730cd50340ffdc0070000317c00000037344334700f40c0c3c4710d0003c01c030000cc004300010cf3001003c4104d7301117430301331c011005d4000017400300003f040ff100401004000040;
rom_uints[352] = 8192'h414043000d0101015c710000030300c1730040000003100c003dc3c074000507030cc3034c0d00c3000430c00cc34f10d70f010f004033f0c700404304074f030c404030003004700100030d07000434c303004d000341041333034cc14f0001c040c400030000000500030c00040f51f04304000cf000010310000c0001010c3cc0030c0000000c0043430703c0c10cf3000100000c0d004cc00c44cd07c70cc03fc100c00113410103c100410100330000174d00c0c0000f0304310100c340017d0d4403037c35cc0304350700f3400103c7f1004400034fcd0f000d1d0c43404000c041070700000f0ccc3000034c0040c444c00c0cc0000070c14c304005cf4030114407c00107000d000c44001703f0c043ccc003040504403c41c0330304400300007c0100cc10c3f1c10001c0040003c7c0c000004400010c000000000701000100003c0017cc0100c1410300c10041003473c3073000073003d05fc00010300cc004300043d334014031c74110000300440040cf10003700c0c0dd0030430f000ff04001000100404000030303000303000c000d01370407441cd0030cf01000f30040c03033000d0cc00003cd0404c3c0030031cc40f7414c7333301d0c0000d00c00000c4f4000fc00c4c37d03c300070045c300030003435100c304d34f0100c00173c3405c0340300504030c0045040f3300350c0300c0000041d300040317f7c4c0000c0301030c070343c710300040000300c44047c03000100c01cc1344000cf4004c40030540c343001c0100010f0005c130c30000000c40044303344003010d1334733c0c00000c01105000430003c3404cc10100ccd14cc313011003c03001d30d0000000007c000c71d0700300c410ffccc01c1004077040343314003040040c0174340c105cf5400c0410300003730c703031300010130c340c0c4c40300003300530303030743100003c0cc3407f003c04d700030450000cf0100000030000d00300340c4000c0004340350c01340040100c30103c303004300000c0c0000c0f70d000c00c37304d10700f004004403030cc344c0404f440d003f000000011000c303c10300d3d7040701003101314700df00000c03dc4000c0d5571300407143005c0003000c43d103c007c100004c0330c3340001000c0c03f0701f000d00df000001030000c4c430c30d00c1f7430c40303c033050004403300000d303013c1413c000010011331f0000030ccc34c00300475d14cf00c3047000030007004713c3430033c001000c40c31300d10071d4030c100f00434cc0c4400700410d3c01c047000000030c054140c3cc013003005100c00cc01405d330c3330f7f000443040d30000cc040c00000003c3331404c3cc300030300c7407500004030fc41c0000100034cc001340300c0df0171030300030001;
rom_uints[353] = 8192'h3300c4037f00c014400313d4f0c4c0c014df410d10c000000c5f0005d0c031c000c54340d71401c4000000c504437d0f71010040040c01c0c01c0071300c30dc030c04d100113700c00f01003004073000cc00c5ccfd703d347011c0400540000c0300cc00c130103c003410104c300c3fc00c00030000300cc43c700f03c0c034474c700cc00010c0c000c0300104003c003000000003000cf071c00dd07301f0c510cc403430300c4010c10d4000500c1033000cc13f7c30d00f0330c0041cc710004400031c01d0c0001d0c0530d4040c3c51c00c304f004030c40c401c0d3330000401447114d1014d00f00cc3013403c000c400010000cc001cc000c10010d0ccdd0ff3c0030c30503000f0fccd4c054c00003cc007000043d00c31303c1043000301c0d0730111c71d04010003f00401701c0400cd0001d044cd47df44100403010003cc0c5041c000ccc33c307cc1c33010340c3f34550c0c0cc0f74c051cc000d100000f4007c010304030100c00400000d0ccc077d03c310043114fd000cfcc70c0001d10003f0030303740300000f1110f70001004dd434003304003d51c01310c0011000400c001400f103043104cfc0000f31f00340d4333c0000c50000fc0300700cc000101c000300300c0000c00cdccdf403430dd0003300333d30cc033000f003c0c4000dfcc0010103d0fcf0c3001d54f3c7c3110340311007c1c370c30c400fc00fc0c7014437000054c7cc0031114cc004300000050040304501d01531c3003014c330034f00047144000c4c00f7134140100d000c131433c3000c1f0c00003041cc71d0c1c7107300c0cc070c00035d0c3c04c0004cc3003c03c3000003037ccfc41d03300c0c44f4300d0f330010710000c73d30100fc7f74c0c530005003404d45f0041f0111cdd0040d44d000340031033015430c4c003010c1000c300007c33470c0c0103030d50031c10d00dc04dfd05f040003fc01400000001000d0000330c0000c30040340007c0c040f0c0c00440c0073074000d0741410c000301040d01d3404003104ddc00cc30000d30570077c003c0104107030c7c000c3000034730cc4340000470005d3d3300c004c04430003f00430700010c001030c471c0c1040001040c774fc3000c11c300d7440d40000303c0f3cc30c35d3000ccc34075f40003040040510710d5c000133f7103c45d1c10037c0f041010000774100001030c370430000031000030304300000740073000710cc31c40001c00050400d70430f0cf04100410107404c04101f31030c0004c00330c3fccd150c300000304c7000304307007000dc300cc0c3303003c0c330f300007333c0f70440033dd301cc000f41f10c0d0000310d0103001430000011003f4c0c0143d030c031c71004170c0000f743111d130d0034000004cdc001300;
rom_uints[354] = 8192'h3000100400c330f00014d0003331c337df07d333003cf314401d3d4000700cf30c0340700d00000cc40c0c30dc10c0400015350113040c3c0f301c10c030031300dc11cc01000c0f730001d000001fc03d7f3c003f5c31070014304c00010170010044c34030043f03000c00011dc304031000c0007c000c000071f0d3007c4001100c4d0030300d3c0c0030010d74100000400000704310cdf3140033303f15d00045f00c010003300c370c300003751131000000107c00c03d0c00750000d4730d101c0c0011000c0340307400df01004110300133303c410c007f01c4c000000c11130c340000fc3410031c304c0000c0f4000043001ccc0033c430d300c331000c30000330fcc0c00130000c0c0c1103400000c070010c0000443c101c3010d10000004000d0303000c03000107030c000d0300f1300f0303300300100310c40300000030110fc1034107010000410340300303c4443034041f0f000d000005000303000d0314000010000c13cc3030c0c331035000030ccf10003043300f30f0cf0c0350331103300c07c1ccf105500431cc000010003dc0c57000000130c3cc40cc773000c001c043101040c73c0c33c0ffccc0d0033003400c0415341d50310103f0c3043004cf300c3300c3340000c04010d3df00c0c0000030100500d000000343d30111cfd0110031f0cc03d51000f3c04101c3c00110100300004401044c1003f710130c01030103ccc7c000c04303010303030031004ccc34d0c01f04434107f3104100d0300c7407dc01c10f4000400003c073c30003d003010cc0c131c00443f0300dd531d0c4300001410300070000000011301003030cc74f330003c33c40000013c330410513c034c04f0c0045c0143140c0c0000003317000000cc030c030c0011053fc3f00df4003d330c0c44c1cf00000407330c0033d1300c303c30f00001f00011001f000d30031304033010100310d73040100cc040030c0131001030701050400000000c1d00030f11000c0c1d00041c4c30173040000300730300000031d00400d000004303ff43530330031030c40001414d1000c1d0470300003f003030cc00000010330c7c0cd0001c10110440503010501c03cd001c0c000407cd110030300100707013c34f0030104c0150c0731ff340100410001c031130330170c0100cf30f3140c3c01c03c430c00001010c0c37340f10000f30330000005031c4300cc01100033030d031331340140330010100003003010004503000c00d10143d3c3030c07044f00fc0041dc0301010000d14700331000401f033003c00c0001711c00c00000004401000c00c330c00000c73033c0f3c3030c0c0001c00000c00c33410d000000c1000700045070ddc40c0cd101c000d001310030c1c00d0140c0041304c0c0c0c103007001140310000340c0040;
rom_uints[355] = 8192'hf40c3c40c3f30f047304144c73530070130f300c0300033cc01000d304540030c0000c54031300c1c07030133400010cc43c0cc340300dcc0003c330133300c001c47010300c00f3100030401030143f031473c0df01303cf03d4374300f410030001013c0f44040f34173100c0f0c405d30003f7000c0c740c5003c00c144c03cc0c3350340047131000030003050040010300c0000004cd0040003357c3d0d40c014001c304000000073c0c430f00c11313f3300c0f13340c3000131000c040cd043d0f01034000444c0104f1c13011c043ff0f337000000400030d00f00300430030537c53c300440050500007000010c5104c00c000014d03031040c00000c04c0313075341c3d40cf0fc41704d00d31010470003c00350c101c103c04130373040034341010404400004171d0703044f0c05411fc003010401d0cf0400cfcd0f3d430d50304c10037fc10c1d44430c73dc0300c3d0c0f43100f0440d40cc1000010c0c051d14c0f14070400c0cc3000cd0540ccc001501333040030033d300c1311cd1410000514050cf000301c000011f340000001cc00c03d40300010330f73034c0030c030d0d740000cc70400fc303400000cc100c40c3000f4c40c0101104c3f00400100743300030300010c073301c1743030c13f371003f43cd7c014c010334f4f007477c0443c31c00c40010113c30000cc30d03cc0014040cccf105cf00cf00c30103004003330cc304cfd4c3cc0100040004d040033100f443070c070c3004003005000041330010304040f001ccf30313303d411107007fc103c03c01011000033d4013cd013330301d44c3c40c0c100051770033001c05c0330c3030130414041100c0cf30043031d01f471dc54710444f77c01100000c00000141305c030330c130043f30fd70df0c3f3311001c33034c101fd30100f4311000000c1cf4d0017003c3404c04c13c3000c0f70403d004c0030300010c333000cf05400001704c00cc4fc40c00037000000340c3041cf31300130c0034534cc00d40300041001000d010cc4130040f77037c40f30c00410c43d43d0300000c500fd003f341534140000003034c030f334c10340003000010c011330340070c534000010f000004134000003010010c000740400c00001340030034000417c1c71143cfc000470c100c410cf01303c00403c34303100305c100400300cc10f00d0000c003000000f0070c0c300000cf0c0c3141403310c1c3d004f0031010055103d033000d00cc111043c00140400403cd003c000f010df107c7430700000031f031114cf3000cc003c14cc3000c300141d00150074304001700000003137300434501330cf0c00400cd0f00c000030010300103000703010c30143300c01d100000034000010043c330050d071c10c0113104071cc00341030df0f00301c;
rom_uints[356] = 8192'hc00304005040dc030c70c0f37f4040110503000000f050d03040000c010c401440c031cd03c00004c41040300043011f7310c00f5001400470001015cc33007001c0400d00c00030d00000d1010050370030c0404001c0000000000000430410000301030f0300001014030051c31031011030c70000013100300c103030cf0f1000000c000f00073fc000005c031073c0300000000017f30c005330004d1055400035001c00c003410000711c0040c03003f300005100301103c03000f00070000303300013c0f1003441c013500400c0000030d0cf1000011440c0cccd00300c0030100f0144407001070c01c010000c3030313300c01001000c1440000030c00c3000f0013010004ccf1c03311030004714000d30400043300007c073310030c0c30054101c0014ff0401031305c03c040053f011410000400000170f0000c40100000300cc00404303c51030c41400374434c1541000445f1cc40c01c3303003c010313d01d0511034f01003f110000c114770f00500c140000000100443f0501401c434300330c030001c00103013005010c00030c3004004043f00cc4dc311d100c00004f3f17101000000ff1c030010f310fcf0703c3c0400cf1c000010037101c454005130cc0300041001c34140000000f0007000cc1301170c0043400c4c000310c04543df0000f0d00111300c0f0133100070117f0001403014301010d07050001cc7050041f010ff00011044400dd000000170c07030114100000043001030f000000003df41300cc3003f703000f1d1010c33010001cc004f40c03074c004c04041073c5310041111400340110300000000c000d000c0103355d001004071000d1fc000c010100004000045c031f101407001f3030000007371400c0c00051000301001400310140c4dfcc7115004c0304000541304c0301330c011140000d0c14350301000000051cc1300f054410010c410004030100100303000030000003030400000fc14000140110f00305330c10c00300c10c03141d3350030c03030544011540103ff0400004100c31f40c03c333c10d400010cf5c171005400004000cc0f10c03d10030033c000000100000100000000044dc0530003fc10f0c0c00c3000cff014301030003170ff31033300d0007000d00000f0c300530f34003000114100033c530053c7134000305c7cfff015101c03017047c10c41410c4d000000137014c3000000fc0c000007f0d500c0f0314000004c0030341057c33000f030300101f105430c0010103317143000000300170000c3100041000700f510d1d1003000340f40301000d5001cf000c340c001130000c0d140007cdf433c0040530303c03070f00000c34c0000003001c341003110144000004015110440c351355003433011011151cd0c5000d107cc04d1c0701004430000;
rom_uints[357] = 8192'h1c344000df1c33000013000007001001010701444cfc4f000010c00cf00c101000fc03c0c03f0140101100030c00715c0fc7003c0c3f01310400731c0100c00c101001f30c73005c03000c004743003c330c00c433511c40000400cc1c030f3040f4003303f01070df3cf0043d140310114040c343ff04c000f403ff03c01c00c013f30000430433300000c301f347d0cf400030000011003c040003c30400330f0c31000044cf30f01000cc000104330543c3dc000004140c30c011037c0c00c4330ff3f00000340f00004730c300101c7f00350030c30007f330fccc51c00533030000c04000000000515d10cd010d5013441cf0440001103cf43013000c00330c03303310311cc00c1133c03500c30c51113c00dcc03104050030113ff573001d000077c03f15c001013343300dcc000c001f33011d00110010033ff304c0c330c30fc01030110010c05103001451101111cc0cd437f704c030cc100100440040cf001330c00cc03c3f4cd01cc3301004005c00030d15100dc0fc04105c700cc03033300f000cc04c0000f33300373000301f1030dc004c003011001d041004f3410033c3cd00003430cc1dc013111c01f00f400dc00303c403dc00300433c0740411010031f001cf000ccc000033003310c4343330000f40000f00103d0403400d3510000005031f110073343000740001c0040400403c40000c1f030c0c331033033401331d00ddc110c03000d0f03733003f0031ff3003141431307c00700000c0444f330000c0011110c0c303d140dc000c3f00cc10333f301c00131fc000d73003401300c0f000f00011007001003100300c430111cc30c30f11030003511f30c503301700500c4140000c30014f10153c1100000530cc301000473130fc1100c4003000f0c3000c0003010300d1013300331c030073040004c00f1cc1c700003f0033fd034333374010f17400c340ff004c00110140c00c0d4000d0010010cc0c00000f034300000033000c00f0c31537c14577f00c1010140010c00300010137f0043c11f30100340100050000fcc3013c034033103fc0370051c111001c10300000c3cc000041030030040710c001000c01300100d0c303040c0400c500410c37013004033030003c00113c045030300000c00104035f34cf30f005fc300100773033347cf0cc3cc0070c0c3f0c0c0051041d3cf33304c050f7404004d007003f0004f70c10040000370dfc1c34c033cf50c1330f1c3300f7111f043ccc03c00037300f00c01dc0c303100f1300100c041d000f0f0103c0000c00d0f100ff040c0f07cf0c035d3001140300500300150000301c00c000c003044f3001d7f0000ffc033004d430000100010330041100010c0f303011c334304c1131c01001000000c0001c1f030f11333431f0014103000cdd100f113f30005100;
rom_uints[358] = 8192'h304000010370d3007f40300f54004013770003c001107cc00403340055f1430030cf0d04330330c040140000d0000f3540c40cf1d14040d001000340f500030d0100c40c00f0703cc0000100101014141c10015f311f1030c03030c1c011c003c305030cc0c00315001fdf031034001c73c7c00fd3d043000000c0d0c747403073c30cc500c000300040040103c34007001300100010350cffc00040f04144cfdd303010000300010310304f11c404c300013c0300300c45c30d0000df0cc15403cf00004304d753c0400c1cd0cf1144033133f0003030cc03f3040500c50cc330c3000404d0c0103103c40544cd0330c33c34d4100300c000c4001014700004cf3cfc005003000005c400c330470030c4350313c0cc103c3c4f303075d3744c00d14400f07000f7c075c300350170010734c0c4c0c47043071101d0110d301300143fc01c777c00cc00f0134070c004304317301cdfc07003311f30110014030310ccf00f40fcc143c000001040c0400004137000404f74100c0c4004f01f3030401034c030cc0043d0010fc0c014f3c400f17440c00403c7c341cc00530c44c5dc01c0d0c0030043030000f3f00405030700f4d4000333c000c074c13170101fc477d1403140030010c0c0130c530c031000c101004c00000cf0c301c433c400c14010f0dc10c301433003fc0c7000d0c0d543310043100c03f0034040034fccc30d33f04fc010043040000c3cd04000000c3303403c1370cd1040f540cc010030101344030101c00005007501034000cc000040d34703f003110ccc000113cc05143070c34003004775c1313505301407300000c01030015f000303c0d344134c0000f3d0030d010330c005c340c04500c0017c040001c071d00cd7d37000304033004004400030400cc07cd075d355c0107007dc7d5340f0d000504101c0105f34c04013d3700050f34501033051c1d340c110451014c00c50300c0343403143304003000c0c0f0001401453f0c0004344c41310f0cc73407100344000054300700041430330301c0400c0ff00c150d015f133c00300700310030344404c4410c30f1c010030150000f1f00c0010cd0100044053030300303410c0d004d0d005001cf1003000047010d404000000000000010074c013d04300c3010c3000f13c4070d0300d3100cd344c000010c031cd1cc400f000031730c100c34041c0c07343c40000004cd010100033d0740f044c3174c00343d7c0f001d103c0330c040cd30041c04310003040c003410070003c3c100430c004300004313001307103000f00431345c07003f0400350500c0001f3417004c10303301000054003400041040000c001f30103354453410054004003d000070410d03040400cd00fc40000135330f03147300301003f40c004100073400c04340374c0c07404c00040;
rom_uints[359] = 8192'hf00c3300c4c1000001f305317c00df33f000400c0000cc03000304d0c4c00100d000013fc070040374440034cc000c31033300c0f47c4c300044c0341c0000c000410c0c0fd0000d0100cf043100013340431001f0cc47ffc4c73c100000771340cd035c00c03c30000c0c05000c0d0004303c4d40cc3cf101fc05c140dc0cc0f73031000cc000f1000000300000404100730300003c70000d00f1f03053d30c30033540540410c4300c000401d0c00000c5c00300dcdc0503d010f0cf0040f403137030c0003000c0000001cf103501341c0cc140c0cd04cc531c13cd70fc00003cc030c1c0d000c07f43c0000033ccc031f345030c40000c040c0700000014cd3cc04040ccc4030040450c00000404143f334050433f1c74c301fc0414c010014c0000c334130f0001c0110407f303fc07000430403000430c00347f130000c10031d40cd1d0040d30044f403cf4c0430cf30c003303c733d0d013007f010003d4334100cc10cc5000c43547050f7f0c540031c050010370d0c0400dc003c00c040000cc407f0001040100c03153cc0f0003043303c43054f0340000fcc00c050f74003700c00001f034f0d51f04f114cc1054145f0030fc010340001d3400000000104c300c300c003cd430001f103c40f3030c1030340001c0331c141f3110c005300703500041741041003000001c030003550c0035c004c000100c1cc11400dcc103335004c40c00040cc500cc511c100733010c070003fc001c03c3100010031c4030013004315030f10401300531300074f30c4d343cf4f00000fc444000c3c0371cf0f000cdc000c0c34cc0303410300d14700404f144030c00503ff3033503cc3403040430007c00103100f7dcf3400f0000c00cc150001030c0c030100174300345cc00f300000503153f0104444035f435c040c73c033c0030330041f44cd0df73100030030c11d0c054110ff0f41f40340c4300f3c0004f04001301504c0000c001c000d0003040dcc000007750034704711c00ccc70103fc4000000c3cf000333c34100ccc0d3f00500c4f300740370c00c00437010c405ccc3f001d4033c043cd04000f1000c000744710c303453053103000330030000050d010c04055c0c00030c4435030003c001c0c0c15fdc5000710430d0013001c04ccc30cc0f0744410ccd011100c3410441004c01c00700c1c435401000f30ff0f43c00c3f301c00fd40001001c000cc5f00001147310f74ff440c100100d03d4303033f1cc0000cc0cc0fcc1c0c0d31001f3400fcc4355000c101370010f00001001c50010100f30f400010010000000000351c04cc301d40400c0400c0005fff015505f00043d03f0000c1c0ff04300d30033303007010530c301144001c0cd010dcc43070c10fc310570000011c3301f300000510003344740c4c37cc1c0000;
rom_uints[360] = 8192'hc0770c0301340cc1303404013c00103c33c000100c0300430000070403d00001043003c0c0c400110041000c000c00dc0333fc37150004310004130c5c0300003403730045c0013c000000c100c00c0c0401001c00cc0d0c34f1c3445c4000400d03000cf434030c04450c0334c07303300d301cc374c440003c700c04415c00fc04c04040c401f3400c0c000003dc4100c3000d0030030410030c004410703001cf3300110c330403cc1001d100003000053300001c00c37130000f0c000001c0d400c00700301140343031c000c57430f70400c13430003c010000d7310110000c04014f0d410100cc00110070c44000c00c0f05d403c04c01040d0400007d03dc0140fc41400dfc1c0030003340001c1f0c5d0c043044100c0c030fc4c7c1000c0700073d340030435007000c014c30c035c3300d00004c00cc0cc440033004c407000d130c000c000000033030c00f0c4d00c1014410ccdd05101d037007c0114010043c003c4cc000300010301c0000dd0c41000471c347c100740d004c0c0cfc3104303404070c00004d0010040c0044004c0003701000041000340d4c0c0d0000010000c40c34ccf40010141c0700100014cf303304400000c11c0507c10134011030c1c407040310ccc0c404040000c143040f0000000034101350047004c00ccc00c5c0001c10007400c304d0c0dc4010030001013100004d0c47c7c10c45037010c4040c040f4403440110cc01c000300cd0c0cf0030fc040045c0041cc100dc4030f304305040040074f000700f0300c10403000305d1040300051003004401004c00c30cd03014dc4c41f0c30c0c00043c400005c404030c03c7c0503033733c7050070c0c1cc0050c503c00004cf40c0d0047f40c00101c40050c00000c0000c045474370011c004c3c150d0d30d03d030104c00400010004007c0000f30501f410c0000c0701040fd004cc3c1d41c10410100cc103043404303000500004001f000007d034c00500400700030c3c0c015004300d31c03430300c0004c011041033000000cc3407c40c3c110c1100030c0d05043503474d00303003404404071d10000000c4340d410334000001004140040c0000c0c000000330500c7403000cc04000c0d40401005c0f000300cc5400350004003004004100000c401330c30011cc4707c010000140010c057c1c0c4f4c10c00000004f110d0f0000530d050000d54d10c01400344704041f370304dc00c33340cf0c4330c0f740004133004d00f11d04100004777cc0c004d0c1430700f4cc330f03100000344cc5743c11c0c0040000000410000f0030000d3f004000040000001c1c13f0000304700cf03407001c0f304d710440400104010003c040414fc3c3c30004404c1001440f530031050d000dd00431001c41c3400c1005003f0c070104404030;
rom_uints[361] = 8192'hc000d00000003c4cc400000c30c300000014c00d01d101000c4d0440000c0100d00700c0343c000000004400401c300c4d0400c00c0004034040414cdc04040f10c105cc030030c1000413743c40710000104c3041c3fc00400d14100300410c0c301040315030c04c030003040000c000340004104d00004c0c4000c4310d0001000003310013fd00001400310000cc007c0c0303030d0101003c0001040300c0c013d000333000010d0c5c000000300037074740dc00034700030000031010040c5c4c0f1c001c401003d4cc4c043010000000104004040ffc0c4c0000400cc154c740000f0c7f1007143c000c13301c00000004000000100403000f000c03034074c704001000003303001cf4030f4417317d33c4040007c7030700373300531c000c3070c30000c01041000404000300f001005c000c0141070004dc000500070d0003014c0130350034040c040f40c5113c40cc0d0533c01007050d31c0c4010f0073c0c40001040030300f03015004c0c1c03703100000c0150003104d00c0000c5700010c704c571d4c00c1000000c00d40c40000500000013001c0014100303ccc44031010d5030c1001400703340401304000300c310003004c030007000d431c510003c00004c01dc0010c53453300010c000000030d0cc3ccc00f0040c3000c10043c00000f0c075c5cf103014031010001400c44401110004d434137100037c00330000d310000013f00001cc50c00000c0001000d400044c303074c030000340d303030000c0f14300000d40700043430cf4c33000003340033030f3000f0f04c00c0344304c00000001dd3c5750417c311011003c40004007004000c0400f10c00c10047100c001fc0cd03400c0300730310000110311c340037014c01304c575111013c4140c00000130f30c001500001000cc1c71c141507c3014c4510003cc7001f0403c3cc403c0004d1d000513314d0143033000cc4000c000c0d40d00c00144d011010c4f03c14c1030310000d0c0014000c300010000c37d0010037d0030c0434100f4c30c10c0c11004d1055300dc113d0000004004cc40d054c1100cfc00010c0f1000400040c400003040d0034c4d34400000017fff0010304070f40f00c04004300f1333400451037110f0c00034033103c3c0104c3c0000c4cc3030d001c000d1311030dc100301043500001d000311c0037030001c0003d30040cc000700037c0c4c40703f7c1d374000c405104c3d30005c000101300000c030735005d0c0001c11411f0cf00cc0c0310f34c740004000000f310dc0cc70400000015001100300f3c000003030040100003c070000370ddc0301f000d0d34030004c0310011103000030400300d0dc0d0c401401c00400453c4c00001c344010010c050530cc00043000000d3071d000130030f0f;
rom_uints[362] = 8192'hf1cc341343403434c704c0007003401300c0034c01404300c4cd1f110cc013c00031f0377cf3c11300031011d307f0001d0001dff051ccd01400440cd030c000c4c0304000d0400040003c14c40c433f40404f4330c70f1137037cf0fc0c40404cc0ff0130cc00c00c01413d0c3000f4c07000c0c00cfc14000f040401301cc300f3001310000400100000000304700d43d0001003c04c0300d00040d0c1500d4070d0401031cf0ccd44034fdd1171c4c40c00400070100110f00010c44cc000013000cc00c1f0103401033133114330f00c4330f153d045f5701c0c30f00430d0000cc047cc40003cc03cc300f00d040000c00407c400c14010cc30f00100d00003040700c4c04140110c4304f030100343000131710cd374040ff3317004c4c103c0003034330143403c00c0400031100031c040c030c04cc700004305f011403c00c00cf3100440d03d07c00100110c000110400004507cc0d341400304f000f100003300c000014d1710030c50d00400103004c40030430c01000007714130433c01c0500313c010033c1001771310010c3300000004400703c0000150001d01310000400130c010000003401cc070d0504d4044313000001013cc15c01303030001700051c0f04000cf30004101010040050c0054005030000d1100500110030c330d10553df30300d04c10104400c3c055c3010330503c000d405c03f000000d70351100f11000f03d411c1d0071000100111401f0c411c4cc53c040140f400000c140000001c3c0405c110400043330c00050c10303f000cc000f7d3100511003c00c110100101c0cc0000041cc4c0434fd40000757f03c40c0000ccc711f0003d03013750f0040cdf0010030c440011c013143cc330111014133030000035303c0314c10f070c30343c3ddcf5300000330304003000110001cc0c541c450c03040410cd0300c31c0c1000411007c30310000f03004cc337c0154000330c04df1c00fc00cf3000c1000005c7000414110500310f040d0c000f3f1cc003003c003d4303403035103c000004d41000c4cd00035400fc150033c1051c00d4330443701400d3fc000110c0330100141111dc1343014011000c03c00c0010c53c0c0004c4010104040004c3005d14003003400f30011000400074010100000d30c10f004c04540000d00c00301100fc0400c0350c00c014100430f0c4c4350d00113c03310003ccc40435010000700404fd04040c730c10c000103cc115003c110000fc000c0004011c171cf7370c0ff0cc3f1f000000cc300005c03f000cd0313f110400d73400000d11013300c500473f01fc00d4003031d400c4c0f0c03310cc1441d70cccf03100d0303001c10cc013070d0f10c0010c0fc04c1300d1c0c5104030c4011c0050330001c101000d00c0404000cf003ff3100c000c0001;
rom_uints[363] = 8192'h33411003c001000f0f0300ccc31034c10f0000f31d01fcc130fcc01041dc130fc145101140d50c1407330f0301c3d5dc7d430140dc5140070c00010dcc000c007005dc01cc010433c1000c0070044003001401f0cf51d1031d1103ddc00040070c3350fcf000301f0c07cc700433c13313cc040f14013cf1400cc71c00c100330037500c003c0050c00c100c0710c0df04c700000070c04003ccc3c03041dc1403c50007100313c405c0001003d3f0050110000000f3c043370f101dc1100010c0c1300100031501f3433fc431cc13130004d03c10ccf000031113c130dc00043f00000c001dddc0c04000c0501101003fc003100050000005014403044040cd01303300001144101340d000c001c03111df10140130713ff0504030ccfd31c00c103000307300030d5030400313501c40041000500030001f0d10c001c010130c0d01051c007705100c030001f004300344005531113071cf1301ff30044003fc043030f005040f1dc0054004000d0000cccdc04c10303043303f454303040c143331034053015347f1f4001c003c0303000004031014300c4c3f0011304030c0115040c03411cc4730c744fd1300101d0c4dc0303330cc0100131000c04dd1c03000000fc300c000340400040040c07440300c7c00111303000d0c04df00fc00000050d350000df313df1033370053d00cd03df303000144f0cc3f0454310d010303f100430013043044010003004003000001341c00133004303d1f341d5f0135133070f13000000003001f00043f000c03000010071104110131dc0000dc00d041030450000310007054400c00ff4330000000130100d04317040100c140014d4700c11730c300033d010010d11d0c301010300110003c331c141070c037c010434734000cc001005c1c0c010f0013cdd00300c3001000103f0c0000c001435d4005f03170134310f50114c00003ff01dcdf00501073cc000030000430c00cf4c010130030ccf07001c1400173c000c44103c31000c10103c00d00101f0f0100431300440303fcc00030333fc043040015c30c04000000301440310f40003401c0003500c040d700f3c40000000400f0401c4d00331003d331000011740dcf13c04c0c31010004cf7c010034c00d0047005000cfcf4400030341031301c33c000700d3000c01300f303134c330001010d011fffc00cc17040c7311c0130d00304f0cd010000010d114004030304c00033000443130103303c010cc0170d03703cc1010004500043f001fcd003030d31f00303003153c1007c3031dc00131345003c034d0143343000054dc1c00f00033ccf303000f0c00375f004111033030101300340301440c5003c1030703013c003010000c04c011c33004100c0c3cf73fcc0330303400000c010d03c004031100001011031f0c0cc11333c00c0030;
rom_uints[364] = 8192'hdcd10153400371500030000c4c0f00400f000c0d010303030fc30001fc00d303cc30c4040c00714ccdd0c1cc300401cf30c5031f0cc00000400f117003d0c0c0140030334130451000534f15400cc030c1000c0004d031070354c14300c0d30400430003c003100010f3010c5df0c507c01c00101f03ff0013133431730000c07f0301500000500001000010033030004000010040ccc30d30f3004001c0d00d0043010003000f00103c30c030333703cc00000003434d000000c4c7c001c3003f001f00cf0300000103100000c1c5c0030f300313f30010c101010041c47003d3000cc1c0cf01000040fc15100070033c0c0100470001040c100f40730000c3c303f4c40c4030000170cc40011c1011c3d0d0045cd3303f1770dc0c434c0510c53300c03300000030cc00f7c000c1400c00c0010c0f033000f10c4c30d513cf0150530110100010700000f3100103f33dc04cc303031fc0cf030c0c011dd000700c0313004315c4c300050f401c04130001701414400000140c0300010300014d000c070d1f4003d043c0c00701033000400010407130103303c4000dc3c07031533313340573031f0c40445010f07003017000c507034330040cc10103054f00f0410300100f000313000d000400700040300403cc00007100004031400c000f4d014c03011443c13000c30cc300c500cc0c3033400cc37c03c00000d1503f0c17003fc713fcc14d0c70f0371c0300f30070f3d0340300c300111101f30103cc0f000f07410000004000f40033c000174000051040003000ccf3c00013d050014d30cc14cc00030000c0f0c3114f001071c0000dc04000340403c00757c53340000cc004034fc30c00d300c0c5f000041dd40c5d01004c4111c050133340c30000101000c130000304d1c003040301d0d0f00dc30cc0c0133303030cff030dc0100c0fd30704c003034370f34031000c3013c001c03101103d00c34000f0cd0070c10000113000003010c0c40c13403fcf41030100370010fc010030c7cc0300004cc00c3014c00f40c4000f4000c3c00133303400c0f00c000003cdc003430143001c40c00300001040f0f01f3033001000d100000000df500307000f013f310000dc030010c00305510ff0c001c05f301c0303cc70001300534c1f4100013f7030c3040311000730417000733337400301c3040070c0dcc00000ccfc0c00dc11ccc01300003fc1005cf10043c00c00730040001530300140340133355c1104c3000301c01040334040074001034133430c0011c5000001d10dd53c03404150000000d3c31f0f100045d40010c300d0307315100001400000004d00cc10413103c00034037f0100300003500004f77c370100004105000c1100c40001304000c304d3f303034354c7c4c131c0cfcd00001500053033070300104c000000;
rom_uints[365] = 8192'h1144000c100000cc0c000000c0440c007c4000f300100000d000c410c004000030004070300003331000443340031c0070000034003000cc00004c100cc00300011c00300000000000740c1044000000cc0004d04400d0104c00000430300030310000000340400040400c4c01007cc000c00c0d700cf100443c7c013310000c0c0004c003c00c04c000c00040140c0000040000000c70c00040000c103c40040400c30051d0d1000000000000300004000c00003000000000030c7f0c00000000000000000400001005c0704070c0004c0f0000c4130040c00330c170300003000074000400000c1000f0000000000c3005c00c1c0000c0c400000c400040300c0000ccc010df0030c30040c4c0070c10c100400c00350f100440d3c3340c0030300044300300401031030303cf01d4c003c00400400c1003000c0000cc0c000000007c001003144000041011353000c000013000050cf303414c0400cc004040050d00c00c1c0cc0300403000000000341000c0df300cc0000f310ccc3400404030c0000011001c0000000000141004c00000401f04c0c3c134000000cc0440c300c44f0c00000c4f000004c0300c01400c40dc0314c40c300c0700d01c04007c00c1400410044f000fd0ccc00cc404000000c30100004000400d00c3370c00474004c00014c04100750000000001400df000040c0040040000f0c0c400134004c00cc1c30000c00000d01100c1004040c40004f40c4c400404c010c3000704000400c0000000014000f00cc00140c0000000c0ccc004c40c430c00c007f0cc000040043c00000c00000c40c0c03040c000c04c0c0ccc3c00000f40cc34003000370c040000cc40430443c40004400050c00c70c40303c103403cf04000000cc140010400010004c0730c00c0143d3f4c00000000f1004000440d0007c70d037c000c30c000d007304c04c0004403000c7000040401fcc043cd70010030034c00000000000c3304003010f0c30c0000dc0c010f03c0cc01437c3d034c01370040000f00100d00430000100000431000cc0d00d0010c0000c4000315c001500c0000440040dcc00003d7400c0000c0c04c0c040407c000004c0030004000410f00c030330d0c00c4000000000040400400c00107c0000000000c001c40000003400f4f0c0c000004c3004f0f00c000004f4c0c030000004c0000c4300740005fc00340010404070000000d000700c000000000dd00030fd7000704c011c01d00040d1000300cc04400003c00c1c4404034544c000c000c013700f0000003f0cc10101000431700c003040440304000013000cd00430c0c0000003341100c000030137f0c0f0300d103000047300c400cc04d00cc40c3040f1c5c04040c4c0007000000300000001031cc1c0040004c030330c000fc4c0104c34400000000;
rom_uints[366] = 8192'hcc30c0c50130000033000000c003013f3011041c030414000343c13c00d070f4130331f3c3713310cc311101c15cc00014cc440113400010c001400cc03cc01003004050000515000001144cc0001cc7101cf01010c00c34303dcdc4c1004033c00441103003c00103c0000c30f0d1f004003c300303011003d5003d30300001330000f54f300f340f0000470c13f350033041c00030014f10c4300c0ff0304c0ff0440040403100000073100c3414f03f0435300110d13504000d0c3010304000111d40000340100f040003441c0cc17cc503000f111c00013d0c0fddf3000113f0003d30d0c0000df0341cf003740010017c000ccc000000100c440000300300101d33100c30530c303433c10400010ffc100d705000351030003fc0001c10c304c00144c010104c33c0040d400ccc30734d7c0131000c303cf443d030103700405051cf00000304300000f300010033cd03c0cf14040cd141c00401005d300430104c31ccc00c3f150057f4c4cc3f01f004103c3340000d0014400004c3d0311cd40c70430c0f4410043ffd1700f1000c000cc00c0071704040f00345074d00c1f307100004c33030100c050000300c30cf15034014400010f34000c3c10004000003c010075cc3c0010c30100fc050040c17dc13c300101001501d35304403c5403000313c3c10c31c00340c03404c10d430f0cc034510c0013300304343403410f343000c010cf000c3003d03f3d0330c00cc3f0001110f0cfcf010cc00100c70003cf0440007c00113f010dccf03313c0c3510000570fc100f103c13c10c30c0014cc1000c000050731d30c01c0d5c3f033311003dc0107400333c30131100103f00c003c41000fc30004c0cc00413013454047c0c0c0df0037ff0d0400314c143c010000c0730000035711d03c005010444c400c00d430037cc00050040c00c1010dd014fc1104300740000c4d3470c10cc003030cf034000300c340d3000000000031000d55400ff4d30044000103d307f31003c1c441c403d34530c400ccc300003000104100c00101344073710541013100c1c10d30c0c00f47c04101417333c1101c3c000003030001f33c710300c30054040003000001c051c7300000c4c1030fc1001371000055110003051000103fc070d444cf000430701003cd41f000d0010000c0043004cc4d030f400013c0c3033131010510030441400005c3c310c30010340f400030400707000c014004d0c400c4374cc440303000f000d3fc0300d007341c030c3001c01f534c017c103333d001c0d730cf0c0000c0104d000d0c44400300104013003c7101cd0c0d300070d740404000c30cd00004d1407c47750ccfc0c00000010c0000030d0000010041000144c044030df00c4c50c341c000503001310010f14040040f3001001cc0d4f0c000005101031003;
rom_uints[367] = 8192'h5010000155503c0400500434fd10013010015034000147700d0c50c00300000000c1035cc1001030c4000010c0100f30007c0f0541d500f30340301fd00c4530c400c1c33134c040000050003004f1c03c30300cc50c7ff1401503300030004104d11c4504000134717c34110300700010000ff1dc0000100c7000f0c01000c4c40470c00c30000031c0f0300000000c0c003000007004000434000c745c010033030c3010c4c0c110c0000cc074003000f5f140000c0c000170330cf00030004110010450c100000100007f300dd0c00014c4c10441c1f00070033c0c1100037400004733c41443013000300d37d0c1710cd0007401040010003c0c014030c03000407c00cc3034d0410cd001c0013fc003d14000007c307c1040dcc00cc3c100d000043000034507f0c4307d41300c300051010c0c0000c000c415f3f410001d01404070500000d01004d000501003030c14000100730dc0030c30fc00c410407f3d0070400034c1150413414c30c00f7304400300431c4053fc14001044040041c0f5400cd00c40c00040f00c4053c0007c0000005034400d3301d000f0003d3000077c01003044c01111d0433310500034f43c403040000cd01000000cc00007d0001140710010330c000000400300f0c100c0f0404c00c100130c3cc000040d5cc0fc4c70013040c40330f0c40310300fc000c00400f100cc304301314d10007000d000500113300000043044d074101fc33013314100310c1475c13003311000cf44710c30070ff4401c0070301c70400011045010c40400ccc00c7c401c1013f1007f11000000740014000000011c0000f01d0003c0c04000330300113314cc04d1c03f300340c5c0c071140c0003311c30114c40c034000cd400c010cf1000040c03003000004f0c0c0010033f3d307034744cc00454703410c300f003110dd110303110000430dc5530100d3c0c0d4004457004003c010400d014013000300010000013c400030100cc014000c0d0f010303031000c03d300003cc0c0001000040d00000c13c4d0001011000d4471f0403d00044404303f300f500c54c04000053d14330010f0c0fc003430f0341310100c0c40c413dcd430f055f1130d34034fc00050c47070010101041c03133040c7c03400cc50ccf070730000034fc040c415407000743010f0000000303003dc070000dd30410000001c70cc751010f1033044100fc0c0730100000c1040f0d50074c0051170400c10fc1103d041fc101003004c10031c0c000400c00d4c03704417d0f114010077c3cc031c0000500110451ff001004f1040c400f00010c0cfd000303030c40000304cf070000435c410f0003cc0d3441dccc00304f330000000100c3370d0d010044034000f01003c4410c0304144303000d0f100c40100540300d310100511400740003;
rom_uints[368] = 8192'hc0f71100037cf0040000cc000034c01c0dc00010400004010df0000774fc44300030cc7c0dcf40cf1c4c000f3c0f4c003c0040c00031c0c0cc40004313000001301c1435c4c01c30030030d015004c013003cc7c104000004400033000cc04401004f41fc10c0045c301340005c0fc004c040c0f1c304404003d0cd010cc7f0c37c3f10c00f0100c0141407000f0404c0c1c001f00c3000c3d30000f3f0130f40010404c405045cc05430703100000d5c0c540000010304010010000fc00300007d7dc433c0cf050100004d0c7000131d0c00c0411f0f4c7c4c0030000c001100000000cc0403c40400710f0440c44110100000d01301000dd40010004304051c404cc10c0740010701400cff304c000005004f3d71034140004c0f033430d000c30000004c40000f0040005d0dc30040030c007cdc00100c031041cc0c5030031000cc0104fcc000350030c4f40c75440330c00043cc1704fc4c30cd0530300040130010c0c070f70f41cc1c05c040300c030000043400f103d3300040040001c01d1c0c05ccc00c47c0d40c0c00fc11000cf0c0000c1000f034c44c00000001cd17400c3cc4cc000c00ff0fc1fc300100000d40001c13c30000403c0c04440c0c0c4034f000f4000f00c0ccc0400c014c30c004ccc730000d0cc3d037300c0c0c0400cc31c13310d000000c4540004c0c0031430001cfc171000c410c0c5c1cc00c0c1004fcfc044007f333cc1c047c7c4df0c11f010300007017c30c10d30c400043700f0f1100030c0d00d40004d3cfd40c404fcf401cc000c100c00c140034003041c0c43c0c04f0403c5304700043c0404003411000700000001c44d047544004030c1340c00cccc0000c07f7054c00c4f000ccdfcc0410310300c0df00fc0c70c43000030040fc1c000cc7c0043c30c14400310300001300140f01f10f00300003400440000c0f470fcf5345d70000ccc0140c5100f0004c1040003031dc0f0340000f014f30dc00f0440c4f004410c1f344c0cc00404c7404704c043f0000c00f513100d00ffc0c745d4c0c433c001cc30c01004fc05c1c03440440000100cc0f4c00333c000000d007000400130003000011500043040300f0000c4300000c0ff030cc4010001c00444504f0003c3c3004d4104370c40000c30c003d5c30f0000104c000000744cccdf0d000c00010c0cdd0c00c00cc300cc0400400c00401100c33c40dfc310cc0301c000ffc0c04cc1445f041cc000c0c0f00c10041cc4dfc0001cf0c01334c0c4f0c0140c330014370f3000c100000030144040c45700c4000134c45001d04c3c4003010044134c03000c00005cf000404314340033c4ffc3c4f4df000f0c4c0dcf100300504c0c34c000cc00c00c0f00fdf030d0d000000004143d300c1cc00d00c4040f3004c14044043f44fccc1c04300c0c;
rom_uints[369] = 8192'hc010c30000c00300d40100000d0000070d00071110000000c0713d34ff3c000700c03307033d00011fd7000441c0c7000c000f3140c0041f01000400070003000013404003c00d03050003370000500c03001000101303000010300300410c00000100531003d30003070f04c01001130041c1100003000000c0054040c34301cf010c10073c00fd010000113c0000043c0c00000031000cc101310104437403000c3103000d0c0100010c014730300f00701000003000d0300300034f30030001c00411000100500001030400000d04010400c0070000003c0400340c430001000100305c000501c00000310337100c01000d000403010000041c40000c003007031c0000330d30100533000c1004510004413304ffc03007c00031d01410110003000000c1c0003040c044330000331c30000444710301030c7c04c0010003d304000111d5030030330033001c00001403033d10310001000c31f031010413c007013c0d00304f03c031c100030103005004001fc003000d13c0010c0000030d04c03c0c010d0105c10c1304035313000003110000cc00f410101303300030000433010000f01303010130c3033c0300cc0140f00c00000010c13003035d0000100d070001040d1330c30110001c7ccdc0040c10040c1101443401034007d4ccc004040310001004040c0000301c3110003ccf00000105f04100c0000031d5300000cf030cc000c10c010313c010133003444fcd0d13101c000c1d0410c701401030c10000c13000000711c00304104110330d000c100f000300717f0000075ddc0c073113000f031c0000000c000d1c15c1110301043140313000040010f0003000000400c004030410300400c00001c0c15730337c1344c0030000000cc40040031100040007000003044300103c107000cc00753c10c0340c4013103100400100303447cc4c3f0d401030c0fdfcc0010104340100c30f0cf000000d000304103c0d00001401340330000cd30037030d001004d0411314007c3410104300c000100c0500104c0033301503000c0c000307011300000103001300100f0f00010313c0c035051043003d300030301f14000f300c003000040330cd3711c50004030043000c00100c500c350c100433c00001c13d0c0d00c15133f7000107373c00000000100334c704c101f40044c037013070055f000f0c01300150050d0005c01003104000007070000c40000c00000000f000f000cd0c0c003000030010100300cc0c0011110df0034d0c310c413403301700c30c00333103004300040c00cc4001300733000c000001041f410c004030000000d100003f1000cf01f03110100331310cc41400135000010000000c031d0040310030030dd0450c030300750304000d003cc30c3003700d0130000400004000cf0c4074034000c007000c;
rom_uints[370] = 8192'hc30cc004d0fc1703c0cf043c03103d103345300c4c1f04003444fcfcf1500c00c0000400d754f0df001d00500cc00334c345331330400103300cc000f0003f0f03003c50004c00d7130001ff0ff010341cc00cd3cfcc00335f04c03030cc441011140400c3103ccc0cf0c010f3000c3f0f034045703cccf0c044dc4c3cfcf003fcc3d3d01141007c0fff000000c0470403010c0000c04005c30c353003010c00300f041014077407000d100f0c4d1d1c433cc400007150fcc0c300105c031000114400100c0cc401103001100d10c0f0c0010007c000ccc0305c00403c0130000d033001c0ff00001cc00001cff03cd014354430c3f500005310040010000030cdfcc3000f4c0010000c307430000333d400f0cc0404c0000c50c03dc44031d00030d100300f0410404303c14707f033041700004f400000000530073fff540cdf0c0c44c00cf303000d00f000041305000cf70c101c0f53f3001dfc5000f00400014003430401000cc050ccd0cc103334133d3130033c0000007cd03030d0c3701f1c00f4317cc7c01000003f37c4f300000c030c000000c314303cdcf00000035c05d0cfc30c0dccff00d7fc00103d400000cf1c3074340dd0c30044003cf00004305000000030fccf01035400040cff0c00711300dc04031fc00100017c0550cc14107d10010c00d0c5cc7f10010f0000340f40cd00f10d003000030cc0f0d0000c3c30105d5050fcfc030330000fc0c0173c130c3cc3c041d1c00d30f304074c15c0000cc00c00030c0cff3113cc03ff340c0cd0003f34cd1c41c1c0400c0004f03f10cc1104f43013103c44003014440730cc00000004c0131cc70c1400dc100c313c1504101310fc40cd05003c00001101f01c1c0f05f3300000114030001f011331c00cf03c45300f0f00c00131730357503100000011c3003f0c0f0340dfc0001c4c11400000574fc53000110017f030d0000ccc410035f330f0033c30040c0c1000fc003df501fc100330c00000540005c3000003300104000c04fc1700cf0031d0043400070d3410474054ccf0001730cf4004fc100f01103cc0f3143000101d011003f000fc01000331145c0f103004c000c4000000f30c0cd00400c100040510330503004c0130c000340005354337003013c005110300c41005500c3100c053c353014cc000c50c04000000c030377c3c4f00d000400c3034d31c1400cd0cfc00c157fc0c0010000430f0cc4c4c1c3f51c047330010f543d00037c0cff0ff0043301400300f3fcc0c3000c34cd0d3310f01c3007444133d0044313000f3410c133004003c5340c0003c00cc30fcfc0053000000100000003010003d005cc053ccd03001110df43c000400cc1300003313410c40c01743cd000c0f0dc00c050d00f0047f003c34fc000501c030004f444c03d00431c305004107;
rom_uints[371] = 8192'h3304c400c0500c5c00000033c0c0c03dc3f0000000043f0000f70000c3c00000000d104010d00c4343c00401310444f311c04f410301c3c0c10000c440c004c0cc40c30100c1000c0f000000c000c1c443100044f7c3470c10c7c0c04004314c00010747000100004307f001c0007c004fc00d010d30007330c070c40373c0017010470f4c0300113010c000004430010f0000400000300c003c0333c03c00c430034040300c0dc04cd003c3070fc40c00c401c000c00f0c000410004f00c007070004c15000c3010dd0004cc34410000030dc11400f33000001d0c1ccfc30514405301c51c004f0013000cc03713013030cdc4c444000c010f15100d0000000c0c00300300f0100c0043f14c0c00c41c0cfc0d00c0000305700030d3f47d1100d03c40001034000c1c10f010000c7c4131c40c33104c00004040d304145d1404404000104104c03c003000f00400f030cdf030000d703c013d1075fd00dcd0000070030400014011f03c0041fff03c0000cc043c33cc3c30d4c03000c300f0051c3071050d13011c40000040c03cc77d4000ff004000c0c33c004c0540dc0003cf10d4c371000030c04c1d00311c0cd031c040470c004000000ff00305004004405000cdc0044c0004704c0c0000050403c00c10c04c40300001004003313d5cc010f100c3c04c0f3030330400300f0c100c0c0c33300050307cc000cd00dc410f0c4d304130040cccf0050434cc1d1301300033300104cc000d4100cc047c104411400c50dc10330ccc40043014304507d4f0c0c1c0c4140c001303000c1070c031030c400000c0010c4c0c00c3cc0d000d000003314c000050000301030c00fdc010134470043733f1f30c303c00c0003c01c10c1ff4010513140330000040c0410f0c00703700d00c004cf00431044107100cc340fc700300004c4c50000c00cc00500045cc00c400001d10fcdf0c3130304003dc3c3fc00f47300033030000ccf4f4f00010005c0c4000c13034f00054c4cc44d0c4d0cc4c0f00f4114f0c000040cc1dd0f000370c0054103c005070500c3c30010cc401347004c313d000330434431000003c00403cd00cc007c4f040c040d000300c000ccc0030cc100140c001f03c04004c0034c004007cc0c0014c0001cc5300c0307c04001f405c00043100d030043c1cc4005340c00074110c104c0403f004f04c0c11000c1d0703030f00334d00010d40c000d50c00041143f005dfd40cd000d0000c040d540c01d40331c000055c1070011534005111c303f30c3c01100c011010f0d00fc40c4cf10000010f400030d00040033c7d033001000730000010c30030000c000cfc0051c33d104c0445f00014001000000070c0c0000334c005507c030d30d0703c0c003c300c40107330000000030530305c33c0c30330fcc00034310c000000000;
rom_uints[372] = 8192'hc000c00c3f3000cc73503371513c003701100041cc07034c3100c00005c3300430c00330df1c001003fd0034cc00070cc01cc0001fd010dc3000c0c03d00700011100cd31104403033000fff4440100473004c3054f0f4c040cd0fc11c3c110fd047f0340c04300c0c0710041031000c0c0ffc4004f044cf00750c0dc050c000044f500c0000c0f4300000301000043c000000000004cc5dfc41fc0430f5cc1f04430400f030cfc410500000433c005c0414cf0c0003130cf30400304c04fc10004fc00500000044c03000440010d5053473010700cc0010400300c0073c00450340401c4001c0110004415004c4ff7c0000fc05c0104041043c01c3000c00450443f4d004c34450c07cc0cc0cf5cc30303c00000010cc7043440c44000001c41c4d4c00c0c0c04c04300054c7c0c530cccf33c034c00c00003c0c0340000030540070c0c430070cd0030000f00040cc0f4cc4400fd041c00ccf00400033300041143000000000c0f1d040c4015f4004003301030130403110c007f341c30f410c333033d00400d005c000303cf1c150030040f00c100c031c1c100500c300004c030c1050303000301410dc40f300cc303033003fff1c043304cdcc003f50c40000010000cc400000103f00c07041cc400003c00000401f003000c40000307344c03f74000fc70c0c33411c043f40001044f0077c00007104034c00034c30c5f000100300451000054c0cc3404cc3c07010701c3044400030f3410d7cc003300c0cc0140510c00300c305000400c33031000040011004000c00000ccc003300110d0001f4c5300c0c7cd0c013000f00c5f41f005000c4000314c03c30301007433000407d4330ff33000c0000000c4c0040003cc031104000005000f0400014040040c0f1c00300c0f044f131f04d134574c0c305d07c01c0330005c0110010c1c4dc00041740705310c0d34f000f010c00d4c330d00041f004dc401c000c01c4c51000000001c000001300013340f30010c30d0005f0374cf0c3f0f104004c4300050c0c000c00434001f030414c010000000400004000017c153c33407404c0f030c010c0f033300f330d0cfc040440000c0001003c40001000001000fc0cc03c0040cc403030101c40041033130c40703f03d0400110d00043c003001003f0333073d314300000400000c300450010c015fc071c407dd4330000100c14f34130414c1001007c43000000f000cc35100000c004470004cc000c700000c001f0c7dfd000c015c0c30001100400014c00034034c34fc0000434f300000100004cc0c0000c050003c0c0015d3c01033c300c000001000cc000701000f0ccffc00004f0c040dcf01004404071411300704000030100143f47d4304d030450c00d30301c01010c4011c001300000cd033030400005040001c000f000c31cc13104;
rom_uints[373] = 8192'h134c0d0013440c50100011400f0330300c140303340d4010040c30d0cf053fd3047cc5010cd0000c141500001510c0c00d1d34ff0c0030507100000cd3000000f400fc3d0001dc470500c03001c0000000314743011c1c031c1d1c0130c31c000431000d0f0cd00013fcc30010043573307c7f35707403340cf3003014040357cccd111004410071c0700cfc1c013c1c103f000c0007410c3704d4c0040100ddfc1105d30003d0007d000010d311013d41450c7300301174f0d0000505110333f100007d00000cc77030103d305504013c37dc03001000701c04100000010c4ccc04c00cc0c0130000010005743503c4001c0030d0d000071400030f404c000f01c307100330717c1310d33013f400403041443c00310c04030c00410730c05fc00434001004330471d10c000713700000f0110c3000d0300503150c043c4004cd001d33101407400c1173d303430431c04c0d0000031c315c001cc703703d10031f3c31f7c300c03000144c0c10f5004c01400003001c0c0403003d7410331c03cf4df01cf44c00307104104c143d101010c03017c00000f31c140c30101510103d040c0d0c3cc4c07c0003d71c411130003110350cc10140043c14f1d00d343144340000000413073430001703304050fc004f0dc4f3cc00c0033c35c053c4c403430403350f1001c0c103700c040d07000000c00101300050c0374c00410c0c00c0d410cc3001033100700dc5d0071010c0300c7c10fdc73cc00f0000350140401313333100300017dc000400f44450c1cf00003000371c1f0441140014df00303c30000f100040c40f0c3435c0000d13143350fcc400010c0c3f0040433331000000d3ccd013c010300300104c3000d4c4403033c70130101c00310000cf00310033f3cc043c7010030c4cc014f33071f0c00c30140c30100d405031fc7031fc3c403135700c0f4c5d010cd70033cc10130cc0f0cf034500dc47c0000c333400c0310000c43ccc00c4073c00c740c01013051cf005317531f41310101337dc000030c140001c14c3304134001033030c00030c01d0000cf0ff34cd34300013100c407d000010131000c00005000c30f110103100c04d114c00700c00111310d700c1173404700000c03400373c000010503000c000741c0c410104fc33c40003001d3c0407000030f033d340f001d37c0c37031700d03d4d13003c000cf100103cc00c140015df70f14001300033000000003130303f30f3300c303c400041cc100cf00030031fc43cf04c330000cc1f0003fc431c3cd00d10d05d0d00d00707000404d0010033340000c00c40cc0037c30414000007340403000cc030400134d47004cc01ccc00434010c30c0340d0f300400401041f0c3035c401300000000104c0001c4ccdc4c100000041d0700000431414401303100c1c000131100;
rom_uints[374] = 8192'h30000001103cc0753004004f0041cd403c001c00c1c10c0133c4000c0d01000000c144cd304000003530000f307000030c3c04013100031010c0005300c00d3034000d0300001000003dc0d40050f300c1d50d00c130003400410400040f3c004c000c0004001000003000c040440000c3044000014d30001034041000040033f01000c01f00013000000400000100100c000400103c00f0400000140c04f1c0cc3300307f40f3c00303000000000000050140000c0f050c00004311400c0401010c04000000110310000001dd01f40000004000f03ff010004000010000000704000003d00000004c0c0000f100033cd00004c0100000000c00000c100007011c0c0000c003300413407340040004030c0c04004d44001f0044c141343c3c04f010000030300c0c00cc0003000001c031c000c4004c000001c000010030c330411000c0301d00000c0300040c001c30cdc3c4353f44c40c030440c03c000310f4370414570c00d031300cc000014c000000140004c05c00fc30c00000c30f070c3110d030004c340d000515003403d00000000000000c0000000101fc0c0041c03c13101c04f000dc003d00000000000004130004c000d0350400040cc1010c40000000304300003544043c0030001c00c03c140404c7000ccc0314040c4c0000cd100014543014d04300000c0500000ccf0144330300000010c0f004cd00cd40000400403c300410300414130000d00710010000107400cc1350040100c0000d1f30004003000000430030010141031400000030000000000103000014c440c7100f400400000007130c3141c0000000dd540000700000003035000c0700f11300001d300c4574c07d33033c0040c000c400700c00050f0c03000040000700400000400000000514550505c0400000d530c0000003f4300400100c00f4037000f001d40c001c0075f0003504c075340400c40000000001500fcc04c000303103130000000c34c0010050c0040cf0000400040000c0040c300c0c010d43004000005c1100f040000f001000300c30400400c0030c10000410044015433000cc040400dc3003141000004c01c04007350400f004400c10000c000000c00c000003000004d0004014441c03310c0003000c134430700000cc040ccc0000000040000003300740c00c0000000fd45400000007070c0011003300c100100004fc0c0c00400010001100d04c10c000100c0404030000004530741000011c0414004cf130300001c733130c7000c01015370c01c430f300c04003000c00c30d0000004d41004030f40d400d001007101000007c4c400c00c03c0100c000003c3c0000340400c4c4000c00404153074000000000c030000d0fc00005c0c403143107030d010043030030000f001410000d000c130010114c00030004c030cc000040;
rom_uints[375] = 8192'hc300c43017c0701003c00030f4001c00d0fc3c400cdc3c00001c04400c0000003000743c0ccd000004407033443c3007c04c000443d0c00c300c1410f0004c0c00000fcdc03c003c3000341c4000c010300c0cc44f0473005c3c0c0403130c040014cc7c340073045440330c40400c00c000000c30d33004003003f01cf010f03ccc10040004004c03cc00c0c00011c000c04030004030c0f43000303000d50c0450c40017cc040cc0dccc40c330307c0001c3c0000c00400470d030345c0030c0104c00c000f00c0000000c1d00d0400070c3d03000c0cc4c040340c34c3c0c700330401400100000f10034400c1cc0c4c0cc40704400003004040c3000c003f0003c00703430d0c31c301c400c00cc5411c47c11d000300440c0cc00c00c4c40cc3c00d5100c30c00c0c107040cc40cc1100503cf400043c30c0000c100cf0034ff0107404c3105000001c400cd0f010cdc0001000100c0c30701000cccc3314fc4017f0741d0c4017f0ccd40c303c00440430400c0cc0000300d00000140470100c000740500000fc040f403c04307100310300000400f0c00c00cc0001003ffc00334c0040c0cc000010c700003fd704401017c411040f3003c44334d000000cc00d001070d4f030c3004c0000f4ccc01c1c04400d3c401c10cc0c400073f03700000044c51c044c000000dc04fc004004c03400c40010300434c7c0404034007034d0c014d000c30c01c4f743d010c110011c00144030d00403003c500000f0ccd03040000000cc0000304c443cc0f0000040403000000c00cc0000305010c4c0cc1c41c030d40740d0700cc01001d0c0cc00c410c0040c001c000d070c1cc0000010d00004730f01c3041c000000040c0c04c4c00c0d000010d3cc0400c0c01003004004000003775c1000070004401410007400500c174000fc0043d10cd010cc0400d40054405d4c4130003040101150044040000c00ccc0ccd000000400c3cc0400f0004c403c40d00031105004d03710000c3cc40d30df04c001300f00000003ccc0c030170cc400100005f040c030c13c34004c145c0030f30000010f0f0040dc00430004cc0c00040cc30dc41400003cd00400cf00d03004c4100dc010d4040fc0c000400030c0001004500014740c373704c01000300033713040740c0003004310c070c710cc300d0070105030300c00040117040000c000034cc70c4c700070f05c41d00c04100cf00044f3f00040d0c00440004000d1f0c0d34c000c3c007c40c0340c03c00cc4030440303c14c4df0c413cc040533c40c4c410c000c0000dc1cc000c1044c4c41000dcc0f3000c040c00c40400c00cd00d00405004cc05fc00001000f0c40000d000331400300000444000001030c77c30040c0000f00c043c0c1cc05050f010003c3000404cc000d00033d05000443030;
rom_uints[376] = 8192'hc0130000000050015001c1c1cc00c017303100400c4c5340030103314cf000040014000d107440330c0000c1c30040d330c7370730003c0df401c400cf030400400c14000404c010100003c0000030c3d001004cf0005103000fd0c003003500000f01c003105c4301000c105c030d3d0d100004440f500d0010500051f00cc3f10f0303100c003400000000300040133034c0d00003cd003c00c3030100c040f14040030c0c41d0400c30c5071f0c3701f4000000000c401010001c5f0400f405313100013044000c000c14031305071030730000000dc01005cc30f114000004040000100300300c5c00c300144dff0c00c13000400400031c50f4130000045310c0f0000f34443310c0f30c5d10300c017113114001c3c41c0c134000003101430c001510010334303013f4c135f00d000c4335d3c00000f0d1f330470c047301c401c33c3310100cf14f000c001341f00030531013301df3f03000101d001007c0f151000103700100110400c40300005300fc50503fc5cc350ccc0000c0c3d41100103404340701341003001503c30010c03c00314344050103c0540f13041110133cc40030001c00304fc470c30070307cc0f503405c41003034d37d71040c0c44400100400c45000000c00cd333340c013005043d0003c00d0000cfdc070c0f1cc000013003c33f13045f00010f0cc03010fc3404050f0340033c1051f4133c43000c0004010070000433104f00c7c3430cf01034001007f0cd0d00f70cc3350c0f4410140007c403f1310540fc77cf5c00007d00f41c11c331001c3d304c03f0d14003c000c30100033000f70010c04310c313000cd70101c50c4c40500c30c05c400c1347d000dcc3003c001300034470d354001310f414405303c10003c0c440c10301033347c45114d00000f7c4010007c0f104533d07cd00c000411c400004034000c403000c3474c3dc413035d0033050030500301050000030100403000f000c000040303c5050001041430d07000110300303330c4000c0000300f0c35000fdc0ccc0000c104000c30131c1c1cd050001c10070fc43c07354000000c050c0000c0300000104401c700534000f45000c00407303743040d35c00df5000cc30c0c3003000033c0050035c3ff000004cc0d30c143014c4cc34c000fcc00c13004430000c000fc3040000f3c113c0000c0303f500c0100cc1c4d0004c431c10140cd3f000f0000f00f30c00043f3004105010733000c4c0033c300d0413043400130343100c3303cddc030005f3534000730030c000307f0f4000dfcc31c0000003d740000410ccc30300c00dcf300c00c7c0301ccc000003cc10017d01d301d00c0331cc07cc3400404c04030c00005103c403000107c0033134c33f00301000004130f43001153f1f401405011550c033005000c3c10301c000;
rom_uints[377] = 8192'h373030003f045c0c07400c0d3443113f000001f00001f1c4044344053040c1c00c37743017530d1000c3c44c00030d3c0003070dc30030f1f000030373c101c000040540d30000344003031500001cf3030401300f14f0001df30c0007100030dc04700c03003df44101df7d00c0135f3d10001f03303f110d3c15dd03735003c4cfc7f3400107000000f3c000004c4000000000013fc00cc030003c0030d47d07337c000700031740d43007000f17500111f330035dfcf3004703c40001c0010450c004f004730c41c1f340301dcc030053cf030dd400c133f7130751c103df000030f3103c013041400df5cf00f30dfcff33701c000103400f0f10007000043cc03c00f3cfc1fdcc0030df1400f0c0f3c0f303713c370000000330730cc000c300c00cf0c1400c013cc0401004c00cc0044334030300030300103740104013050c04000403100dc0c0cf43401330300033303f31c14c0c44040751ccc510dd3000371f137133400d04503f00c013fc0001cc4003000001010003413cc1010f13017f3303570030c1040043100fc35fc00d000dfdc3411033c340c50d4c3c0035fd03c0c35f000003f73407400c3034010c0c0f1c040c7cc010c11c0f41c0131d04004000c001c3011f1ffdf113500c4cc0010c101000cc0c4450cc10c30cfc504430c0d311d30fc34d00030d030100000c00401cccdcf110c0c003043c440053f4c31170d341030cc43cd11c3ccc0d130d43704fc3133373ccc0f0c5001d3103014003030003f0c00f0434404c03344f1c0033104013030400c001130d03030c3df704cc0c30000c3503c543c1c00c30700300cdfcc3c0c1d01100103c054cc5fd333130001c0c00433ccc04000fcd70103c103311073c0f00dc1f300304000403140007000013c07c01c1c0030001f5cd014301330010cf0140cdc4371300c3c03c700fd3c40353040fd70dc1f3cccd54403100cdf0cdccc50000010744c7000dc4404000c310407407110303510003003001717070d550c3014007c01074300331004c3113c33551cd1c31400c0151000004037030047c10c30304370dcf010c0040fcc533d0000003c0004c103fcc1c0040017311003cffc440cd03010cc3003d0100100030c0f001030c010c407c103310c3f00001c30c043030f3d300c0c00031c00c0101330cc0030cdf1f00013c0313c400003d1104730700f0c4c03440ffc0c7100c04070fdd0f400700400c03dcc000130cc30f300710070f413143cdcc0401141cf40301fc3304000cc40003c1c3cc3d3cc34407f100fc0347100011103040cd330300c3130400cc10c0075310373000dc0100110000f04c1c3c034dcf004c0ff3f3001d33003cc70450c003c10030330fc3c44130430f01000c0310000f00c0133000000311170c40f4403541c01300c0317c7307500000030;
rom_uints[378] = 8192'h30c3c0000f1030cd000000000000c0c1030300104cf3f334030fc0300033100413c0ff40c00c000330044110100004040f00003cd701003033fcc00414003300c03041d1000f000000000033000c04c1c0740f03c347c54040034c04000cf53c1544301c0410003133c0f0100000c0500100010c0dcf040430140300c0544403cccfc0c0300c000c0c000030c0f00000300d00410010c00013000300cccc30010cc3400044400d7001c40c4003303731300f0c00004000134d000c014d0004c0000010010003fc544c7000111d40c5c10031400cc4f0030300d1000cf0d0c0f01c0000000044400003d0040334dc330344001dd513011000400000c0c00c0000cf4400d041c0ccc00c14c0330050c40044f0340401330c1cc0000c431fc7c04304010300c1c3c054013c04001c0004fd0ff03c010110050050330c304cfc010130044c101434000330000cc44f4040003cf3f00c0000003f00d070031405f04033c30c004143074c113c510d40304004100000000400c3040100f00040000c03430010103151003003040113c003300d03000c0033003c004d0117350cc300005c1101000c01010000c10ff0f41000f0c7007f3440300000c35000c3130cc303c000000403c0413034fcc300d00050033ccc3440003c40030014300030c34c004c3010071d5c1004c040c300000c40000400030100000c0c3f430040010ff0c37c000000003c0d305000c00cf30c403030403f0013341031013c0f430000303000100447540d000000c177501c003c04c4100dc000f4300c0f3c00103300301337003f011c45134c4c004300f30c043c41000d30030051d00c3010030c3070c030000c0040014c40304330043310000404400005f0444103104cf1c3f100ff300033431007134300f03c000030105341070df44c40ff100f00c041003f04104d7030000003010c113c0cc0f00cc70c43003f03c05010c440c101cf1f011c110fd00000000000134000c4030000104cc000c13004410000c0c0001cf4141c004430000400d310c03c00f135000d000000303c0c0c33000c1003403030334000304c00004cc00110333000c0c40013000043c34f370500c00c00c404030c0307c1340c001030001003000c04100050510000000c0c000000f0435cc33140000cd010100f4f0c10f4010740c7c40c10003fc0f131034414c0000140001003c03c701700cc03d04f00034300000340000054f3d003c10031155105013001003c0f0cf000000030004c004351c0c73c0001430f0f07c330c1c700ccc1c130c00713040140000d5007c44001c0004443c0f03000154450c7003004404c3000340300000011cc31107130c004001d00100000000010300000c1001d4010c07f010000341c00040000f05ccf00041c00c1035f031713c0c040030533c404010f00501500;
rom_uints[379] = 8192'hf400004735300400c700c7c10c000d00440cc0cfc34f3d0cc0003004d00f110301000011fd40130113041410d004c307317034140040307000300d3c5403400c003710c00c0001c014001c1100400000410041010004300004011040330c7000c7500003c10cf30c040100400c0330041c40101c03cc0040011fcd011007c400cc71303f0430004000000044000300473043001100cc04003d4fc3114c4304410030100c001c30110c01000114100000443c0d10001d3f4cc4000000400c03007c0c1c3000c304130c4c03110fd00333c0300d43cc3044300041010cf074301100c0000cd1d410104c4c000cc0000c03c00c4c0d0034030404c4713cf1c0001400100000c0014c31430cf40c04100001c373c4300733cd14000f7c4fc4c703c500c707007c1d07c0004c410c000c0000410d3dc34045c40010045703503041040003040f00c1010300430d030705001c070111005001400005001400101c0010403033301c100d04c40c100305c05000047004c001c3ccd513313c03000f00010fc54340c050c03d030f000031007cd00c3000c00c003000d0010400000d1103500001000d000013001c0300f7100330330c0407d031000f4000001403144f03014c01040c0c11450041300f3dc0100c0d300401410fc77d0000300301031d4f14c1cd10c0310400c0c4070c000104000100031c0700410405000100c14170fc010010c03050c73f000c0cc4714114043400004411040000010c35014d10414c040101f0400300c30003140404030c0407350000400c0f0730004c103400010f400340010140c1033713c4000c0fc37c4730000c4c0f100144f51003033037cc34005c031303370104040103c0000d031c33ff441fc00140444d140000430dc00004c5041400c404c10730343310d4c5100c030003d10000000c340000c3140530cc0f0c4d10000c310c0003400d00170071fc00140c0c1400037fc1000300040c0100000300000543cf30c40005033d0041c454003c4000fd0003c70000440440000c0f3c00704000040c404007017303301c05c000400540c040d331d4ff040d04cfc7cc110111040000474001400141000447030c04000c0c100c00000d30cc443373c4100df00d030300001103c70c01fc0101000405303037310c00c4d30ccc15010003f0000cc44dc7d40dc00c004c1c17c0370110000d501cc0fc4d100c0cc3130c10030144c4400cc44c400000c4c0405000030033f10344c035354c40030c5c0003103c30100f53074141510cf400fcc004430340000f304f0700c35015cc0510f30cc5303311c0070d307130c51c140100000d13010c00300dc0f14c07f40cd7440c3c400404001dc4dc033c0cc050000f030c111c03c500c000030f11130c4501040300c44f000114317070040f0f000fdc03033c43011f001300;
rom_uints[380] = 8192'h7000400000000040c4003404001c0300d0c340ccc03000400c7f0001400c10400030111c70f4c0004431001034004310c4c0c0c0430400c00040c10c4d00c154fd443c30403110c000001310c5c43100c100c0d0cd315c00415c0c1140dc404030f01001140010401071340040c11dc0470cd310c0001050410f400300c5000dc4c3c00111d00033100000d77c0003cc001000c500313343c00003100f13000010074413010c011c10f01f1133030040300c01130000350c00040003f0400140403d5073000033d000000034f0c04040003c70000044f130c030c000c1fcc0130007004c041330501030003f41f001134000c33040300001c4010003d04000f40133134f07000c1c10c0013073cd31c5f14f7745c0373110530073f03c31c1c000c03300001cc03c0001400040004043c00031300000c000000010000440300404fd00d0c0c04c00000d00f04000c401430d10c4c0305034000f0f0007c000340100c30003400100040000431f30c034f0d0c714400003000040cc0c000040000754c003c50403007c0c10033300cf73c00000111000043040c000000c03c0000134100044cc00001014000430df0c0c3c0401c734c073007000000030d01c1d4c00313313100005501c0000000033035fc000d3040d001301c000000c00d4fdd100000fc4c00000504000014fd00001f1310044c0300000df0044c050000f700d00530400000030104040430404010030f47014000043401400c730700d700030c0f003d441005400000c3053cc0040c0341301007401d0700703c33000037000c400141f3010000ffc4c403c0f101000c11003003000004d30001c4003f05c3c1f131300f300300400ddfc0100004f013000dc1010300cf037c4700c03400030dd37005000000014c3700f7c0d34c00f71df0c0d1045401d301170504d00f70037703030c7f00f4003c3c40f0500300df0400c00504100c000430301c40140c030305000000c10cd330c1000013300cd00c0c0014030430fcdff001cc0f300c00030703f0770d3300040303000cc03001004105d00c03043304400f131004410f34040d000c0f0100000f0f01310441000c0003f07044c404404300330d00031030070337430cf34310f00c0d03030c000d0cc04d14011f0cf04f5040000000cd3d0330c00401330c0301c1c0050044074130100f0300010fc3d00035313c10c000030430300070cc04031d140f01cc30404040410c07cf41400c00c4043f00170c410110044f0d40100f5c11007300001d1fc4cc3fdc044000740c000000c50003104344347c0c000101000400351c000c00d0c0044f0d00100000100101130c000c5d4d41070cd0033cf000000c0300000310101101c4070000d0014017c00f0305f1330c1400c030541300501041c000040000304f10400d05cc0003000;
rom_uints[381] = 8192'h47400010707c01c100417cc05c310f11c30c0400c0440c00000c00c341001103000c0040410d10401000c0000c00453440000370f3000c0c00c000c0c700030000440dcdc0c03c400000000c0f00cc0c0003c37003c05403000f40c434330c04c04c40410070030c1c004c000334333050000cf00c33d07404004044cc00004351d070c000000c3000040040040010c0c014cc010000403c34004070cf30d04003510d00c01001000d004003c3f40045c00f40c100c0c001c74c00104500c030c07d0d0c403000c3707100700000df04007430f3005000c0041000000030000c4040000010cc00c000410034103500c434cf0040f41000cc000c50310401c0dc330c001070c0013fccf3754030400040c1dc1c0f00100004301040c0c040cd00001000005114f3c0010003c00c0cfcc4405141003400dc00cc00c040c04473040500004c00740400c04400cf00031010d054400f001c443f4c04334000d1cc0007c1f3030c3d1cf000400d01400100330000c07030c000cc1030133400000c00f0c0ccc04451f0003c4400700304d075c00010c0000037000500c1c304147003c10c104c0c4030c0000dfc0004f4cc0330c000dc0d7341300074401cc007c0c0dd3040ccc0c0c00c307440000c00d1c0057cc0c040c300500333000033f4d030403370c0d0f014000013001044d004c000001001000140cf1001000330400170740cc53140df00103d3141004044cccf400d331451fc0c000c500c50d070010000711c00300540c4007504c00f0c43c030710c3040c0304404001cf0ff0070300110c0003030c00000c030f0fccccd0000f0000c00010c1004430010d000100440c000000cc0100444003100c00000c0003000c0c03000000033c144c3007c3c430003301c0c0000010f0407530cc4000401d744c0000010100034c04cf04010001c100c7c1d103401470131307000051070ccc00c101cccdcc0cd4cdd040000104000000400004000ccc00000000440400c43d44c10d0053040003fd00030c0300000d0f000000c0070cc7c00cc4c0440031313300040003f0014004f00043010433004dc0c0100000cf0cc00c01f7304450cc7d010d400000c0ccf4fd04000cc370000f000000000010300404cd0c00040143cc07300530070101730114410c0f413c310004000c0343030fc143c13d0fc0cf030f000d3ccc3300004c073000170d0c0d01c00c401f00010f3000c04000c404101c0df40c01000040744740030001d00c00040cc00c00cc0c000001dc010c014101007c0c000c44003c004000fdc0040c300d113c00000c0c300c043c0cc3c04c300001d0c001100c0c0101400c45170d00110000004c07030c00300010300c101d0c00710003000cc3303c1c100cc004c0000fc3001f0c03000100004c0d000c00c1000d070c00c00030c00;
rom_uints[382] = 8192'hc4c0c0003c007dc3c030000034c43010dc00c004c004c070001003000c03c0000001cccc71f5003c15000c0113000104f34cccd443c30040041c0dccd033040000015c714f3503130d00f101f330410003f004f430dc000003333df74ff1400010c471cc0c00d073fc30c11100c433131003cc45c4444014000dc43014070c401f03c0f3000c0050c000c030c00171d00c050000000003470130330cc015104035c150c0000c0500410c0333c0130cfd00333c300001f3040100341c00003000304173f4000051010f05003d3f0054400041035003073cc00303ccc40f0704c000c1004f101f1340000003f30c350011c0c4c00043040043cc1344030c000011cc3c7040c1c4043011cc0ccc03d100ccc3311f0f0f013d0c470c00040133140dc3d1d00003c03007c004c3103c0070c301000c0c1704d000000c3073000f11100373c33cd33dc005010343d07cc0451300300005c0047f003c0001c03153011cc4f300000031110c11710100303c33dcd007df33134d001c01cdc031430c001311d53500c5c040040cc00000030030c010000000470000431cf741cc003407d344f145047c330457010130310007c400f0d0053301c4407c4010cc0114cd100d417000c000cc107010703cc33c40010011c00003cc340c750415100000040f40c0c03054c0fd330107003f000c1d700413300c010073c4100401073000f3047034004fcf13c10007d1003100000047c010cf33403c1c0c0043c4c5c1030104041434000c000307000f00000c01c0004c10fc3f0010700d04133c00c0c400c13f40c30400010c0134c0000ccc33c44003cc00c13000031010c040740040130c3d0cd00041c10d00c00010cc1013003133040c000530df003110100435000d0010c04001cc5d0c43433103c7c3f3c0d00d7003c110303f0c50003c3c0330743033301ff400340301000030fcd4301c015c37003000507400d014c000f31001013003317f41030010000c77000000100d040041c0140345c70c34003c50f001134c10000c40ff004d10000003c4004000143d0731f3703504003000700143510c5131003fc3c5c3740f0c000c10f0000c347c0710cc00301c74100ddcc0f111040743dc004737c400000d03c400010504dfc00cf30f0c1010000cc0313c00fc004013001140f007310701c713d000004047dff04fdf301315c3313000000000300000c015400030c01000cc013003300001c030cf0414401d31d43c0300c3c301000110c30d01310103004100c34333c03f0ff3140cfc11c3000000c434c41c00000305001c1c0001000dc1011d13c30c3c00100f100100370000100000104f303c000c13f0013f0c7f040004010c100c0d0304040340c400070c31d1310533704f14cf4f4011001cf1c00f3303000000017d0175c007571c1c400001710300c403;
rom_uints[383] = 8192'h1400010003d053430300407df3030c0c1f00305c1310dcc10c73cfc33003c4103c0cc3715c4cc00110513d400d00031c000544c0c003000c1c1000101401c40030d03300c00c000d4c003c103400c10c50c1015040410d07443030f007f10c3511033010c30d0000c4313f500313ff1004c0400d0f0cc5c0000c4ccc4044c0007700c3d30100c00c0c300c07370040c00405000c000c0f335733303cc31cc070f41044010430c30000007004cd0c00300071030400010003050000005540cc4c30330cdf00007f3d4c3000100100c7c0c0f3c4c113c33000001f30fc70d00c3100033300cc4c300c0cc0501430010ccc10c0031c4374c00c1ccc3c00100000fc103c3050303131070ccc37f034f31c4dc01f113140051f0d044407cc130fc77004000f000c0000773c000c030f00401040c10f1700001f000c300f740cc10000cc40f007101334000300400030471000c0d001d010f001000c30f1f050c00c0c00c1000c070c3004c0c30c05c7c71cc0004050c00c301300107c30173007040c4f04530cc0700c30100d3000c400cc303000c0000c00340103cf400000c000c0745c003030d4110c00f10300f77cc0cf07030d143d0070040f0007c01c04043103710400cc0c4cf43c403fcc3c307100c44c01435c33f3403070d30d31c0c1403003030dc01004f3c5cd0004040007314030c01d4c4c000d3104c41cd430000414313000f00ccf0010c0f414f0310c0035d304044f0dc4c43030d3100334fcd371304c4107c3405400f0d0040000040cd0100400401c00040034000104004cc3d4d4c00d004c1c071307000403d30cf0070000c03400000117441010310c1014141000c003003010001ccc4cc00001ff53441ccfc0000000c30d1104dccc0c0003f401c3c00c40c0c000c411141c4c30c01510431c31330c04c03c00c1130d4400c107030c0c00fc0733300c0330c04cd74404c07c04c4101c403414c40140c4000cf030700000030c0300c0c30f300c000f0c1c00c03c17100700dd1330f301000003000c000f00000330030013040030001dc430314033000cf1f00c3c1134070c07d5311c0304f033ccdf00700c0c10301cc0cc5c410443c0c030c0503030cfd0000c140c0303d3473d00000040000c000475001c0cc40000400dc0c7351d404c0134304010c0000d0300514cf0010000c0f5105000040104000cc00fc00df030dcccc0fd000c30cd5300000c03010400f00400035ccdc3c00003150057144350fc03300041031005070400303c013004c010c70cc00001000001fc010000037d700c4300d4c40300f1043133c0c300513130540000004001f000dc303000400037fd0d04f340000113030c000d010440f050303c00fc0cf0500040300cc030000c04300f31440404d00041107000fd0c00000c00c1001c05fc01c0000300;
rom_uints[384] = 8192'h500001001000307000045f0055f530000474473c1500001d04f10c00c100403334c5d04500504c00c030300000f000341ccc7c0c030005010330d00011044350c0000c000cc30000c153c100430c30300004300d431f030cc4c040114c000c10fcc00400f1cc1c534c4cc000c003041f4f104c5033c3f03d00c4c0040c031117400503c304403000000f41c0703d0000001000f0d0000004d010c0543400cf1001000c007701033c404014f053f0400f0304005031c00734000c0fc033150413033000d0c1c1103004d4000130f0034015c037111047f0c041c3131700511345c03010303430003001f1001000f0cc013fcc115500f000c00c07000100fcd1100413c0f54550c301545c410307003350303c044701d4d00d41001f037f00c100f0001404007000101c504300330000440c3f34340300cd000030000f3c015c003d04030301343c1c040d0110400441f451c000311cf30300f51d007340003000011c1c013050704330000131c504000135041050410cc447153c001c000c0c0733f0473d0c043c0010c001004003f0003000c0003c070534c0c0040000003513070030c000c000300c00040c3d041001744c570c000d0c004f0c0401c53014c0c53000000403c000004007004c30c047141040100c0f5033cc001f30003014c500f010f00c00171043cc10c000340003c031031000001414140000055c1c0f0000c1d34000f000c33cd0001434f01c034337c00051330030313035000700705500fc130400100050c401c40030c00053cc0000034034037c30040400010440330400003000140f310c005c500f040030d410047070000c1c1300131474c3470030f1fd00c0100304d003c00d005435400f3040c3f1040000330c00015c03543000130c00f0c3003530c053100533c5c377c330f004050100c0101000d307fc70000f0000373c47f3337c0004d373453c300014400010373000f0fcc0c413fc50300000000403030f00000030400700377131003c345330c0003c30303c003c00cc300100074c00343000005350500c5000530000300c10501c00441730004150001333003303c100144313c0140c034100c4000010013c300c3cd501040c34c500000030d030cc01cc3407000040c0114331cc5000000f0d03040434531cfc000530434f0000c0c4100c00004410000cdcc4c404c110437c00c040140f130000300430c10030d0f01003fc0c01101c1c17500104300c4331500031131043f150171c00004d3003c03c70000007c03043cd443c0c0030300cf01030f0c00cc00003d0f01430504cf007c03c0c3d1c0c34c3051f0010f004004000441103c0333311c03453c310071057301000100c044c0000c03c0000c41dc3003010c3004040c40040003030014000100cc0f030c0f014f00400cf3cf000703304300000;
rom_uints[385] = 8192'h1d00c000715c1c44334034030f040f70d040000000c401c000d4730000c47d3000d0473c103f0330333f3d40ff0334f541c04404c010c0f0c4000cc04040c3031c404cd400dc441c00004c103300100c54d40370d5cff00130cf70374504d0c00337c4d40330043170d17f001104140103100c03cf1003071c0070010f440411cf7403301134c31f00d40c401301500343000000000c30c0001fc33003103340040000c00c7d0740d00c1000cc4c33d1034d7f0000cc01400003403071c4cc13040014dc30001001f41500303001d40c301104d300301d0000f10c3510cddc7c003004c0c03c4cc0c40100f3cc150fc00410300f4034031c0cdc0d40004c00cf000454713430051310fc43034001c0f0fd3c00fc00f01c03340c10011d40c3403300c000310140000040000c0001dd0001d700cc0cc034003fc00c00df3c000344100504f43070003c0300104400043c010cc0c0003fccd4c104c7331fc1014013f3c310370f115dfc305f10007045733c07cf7c010c5c0030701000dc0c01003005d100334cc0005d100000334003430c00030000000d1c033cd70c700470c07cc034c3145000100c050cc341353300510304301ccf500014f03f74c335405400d0d00000c0001407d100c33c131f00c5303c040c45cc44000d4004133c03f3030000fcf03001c0333d40cf070c00d01fccf010cf0f00cf00773f000000f45d7731c477070c1f00374ccc74047000101070c40400c10040cf000c3c40d04505354f3c00011f10040004cc00470040ccc43403c1c00f01000c0507001104ccf43034001304ccf41000f000ccd0140301c000070041f04017001c444005f07f4130330c005f305030c000c03cc34000040040dd0f07014000c0d1030000301c1000dd10c00000304101443cf33001dc30f000c701dc340c0c054c1c0fffcc3430cccf00ccc343d4310f401c05570030cc400410001f330f0cfdc0c1300f00c40430d00c0d14000c050510c443000c10300113d10710c3c3044040314000f0013050001004cc30c03300570c0cd1d0dc070cf40307c0140c00070000c000030c50f0c440c1c4d031073040c0cc0c73100c047700c4c7c00c533d7c0c1104100c00ffff0003314040000f0001073015311401030c0440c301404c470fc004304430d1301001300c0004c0c0d037000c030730040344111c0053d30c040c00003400f003c03f304c0030d7c430f04000100007400704c05100c5143c40115d04c00011007f00f00c4c003003000113053033300c00fcc00710c01011ff043ccf07011010d0c31333470d0cf00101403c007c00d0c3400d307700cc1c0400cc014cccd000f734014704330010003f3070004c0c0ff0c015c1053cc4c0d01dc10f101ccccc3c00fcc01d10144c03440c114c00f0031f00000d3c104c40330105000030;
rom_uints[386] = 8192'h110c0300050011c410df0c1330004f01050f00c3000c1c3010347f1000f3c110031c1c0cd3c304007c0c000044030d0730c355010103007c01010000f00441d0034d030c13d100550000400f00004103141c4005d004110003c37404c41004344d007c00700100700c3470f00003c0d04031000043d400f0003c04113c13014014000d0010370c0300c430f300001c35003c130700000c07041c04140cd0d30c330c0000c4010353413030001c03031045cc04000000077d00070c3500043310013d30103d004000040303d01c1103010000034033101c5005011f0441c30c001005043001401c33c001c040014d3543f44407c40c00000fc00040004003300013400300450541003c03d10331400001430f4f0d3000c0041447004000cd40c3014c33003503001c410001011c0c5100030330df0d540c104c0001031cd100510130d4000d3013030333030004cc3f0300d0cf01007cf0cd7f103c0430300c70041f04ccc4170d00010c4c0d4700c030040f0d0414c1000041c75f000c033104330c0f03cc4075cd44040c0d404004c007000fc13c00c4000117001010304300031c4f033c300073014d07c3d1047d031300cd7c0cf40f0f340d5f030005f7001f34040d041400441010430f3c007c00541c0c0300000c0300c3000c0030c003d003004301300531f41d0c0c130301003f0c433d0f0f41000c030004c0c1c15c0000300003130c3000c10300cc041304431007c00f050f1c0c4c44cc00c10c3105c07cc041dc5d100001d000df10070031f01400000c040000cd1310753004cc0df0c5100310300000f130100f0343030c0011100033004400100c3cc00353fc0f3403174f4343c401c01301c33333000307f031133c11c3001040000c40077c1034c500001f10dc01cf141013031400c4010f03001000f4000304000713c00040350fc00c0c330733130c01ccc5311c7cff104f0c30301c4c4c13000c0cc01d0fc3000000000000100c030c003017100cf13003c0c04f00cc3037f03010704cfc001000130c03000c0fd3c703300d04d504004c040003ccd00c4c40dc0007000c51000d4c0f0030050003cf1003f0c40005300c404004300cc3430c54000c030001000000300c0043f0450100017330440000303c444400f0140f000d101010041413101f000c00431430040041c0001c0c33430c0000000cccc3040c0f1f4c0010c013535d00033c044305f4033c0c33003c3100013f003cd0001d101cf040750d0c00100054000304c0cd1cd30007070f07c00c07f13310010403314314040400c41033030c50310c0d0700c40400007f00000400c40f0000f40000144300000c4df00f400f100040c03403400c00dc0070000041341d50d40d000d04131c00143c1011fc000c0c30040407403f00000c03150d0040310004303c03100000;
rom_uints[387] = 8192'h400004f003303f0300004f140000041d14407c11f43000ff003000dc47000000000500c303f05014fdc440103c5d001cc0f44000c141130003500f0c3c04c004cdc444c400340c00c0313000404c1c1d4c1351304c0c00c0045c00c41f0c00441c3070c4df413330c034310c3001304c34c4c0300043003037d50df0344033d4100003cc0304001c004000103730c004c000000441000f33000730030fc13c0d003004115fd0f04d1c50003004dcc051030000c1000cc035105311013045d0c04010100010c1c40031003cd0401034dc010001333330f0cfc0c0d03d453000c3003c40107d013505100341c3000000c335507110005000000c0c00000010f4000401c4c00473000c03c05cc40304003c407c0cc0fc34530330f00f00f03301d00d0031003130c00430c50011470c0c33003305110003ff4510353000c0dc5541d00003d10300700d0ccc0344003c307fc100cc0d3000400fd0f300403c1030100001f4003c431c003334dfc310053c4c1134003304d01f34c7000000c3103c3041f0d11301073c10c1340f107cdc01000433100cc430d3001101c100c10003301f0331000c0d0434000341015010101000443130c00cc11070c3301f00c0f14fc4100c740051011fcc103d00300cc0d043400c110c35000f1005300f00f4041000001f100c0c0f73334000f11101c73000070c0000031000000003c0f170d01f3c0c100c101117030f3c10f45cccfc01100cf13500353430705000044100530c5c0000c4c43300cf5300301033101034f70104334ffcc3f511010300fd7d010c004035311f03d0f00034c00040030000c30000400103000401001f7f0535400000fc371cc00f740703010c104c0003010010304003300c0c030001f40001001f0004143140013410014c7f001cc000c0713144c0343d0c00c0001c440104307700000030cd05c00dc0001030000370dd4f51cc0330c31000754334010004cdd30401000005030401100031100c4300301303131000d45c0c3d0c13303000c100740004c40107014d3000fcc0c0dc0c5c051f0001c400343d0d1f0140c1c0f304743f301c00d45300c105000c0010000f00c3c005c100300cc00d140003017c130030171074103c4c010300510c05f1c1ccc33414440040df100fd733300d300c030433c303003030050303000f010000043003000c404c31dc00f070410703043c3d71c4001dd043c104d003c000c334c004f40040c50c3000d40c0301c0f7003030cc0030300300c0000000c03c0003c00d00d3100cf5351c03dc010014310c0c005c4000000000c4c00c000c00004300031000130400010f00400ff0034040cfc4c30f30d001000c04401c0030f400150403c403cc30d0c34c350c3c100d004010cf0031310070031000030151c3000001050173105400df30030c0c00;
rom_uints[388] = 8192'hccc10003cc104003f30000000000c0503f1500c00c00d030004005330f400f31014131105343000073734c10c3007c10cd731071f00034300c001cc00c00c00c00400040c0f050170c000110cd1000100000000df0c707d0f4c30df000000d01c030c04000470d0314c47100c033c0c373510c4333cc0d00c0c0005f3400c00003c5d0033c100033010d003f3c0050f1c000004000001c3010000044c0741000030043000d71c00040d004c0c443003430d0f4d00010c043304000c3300400004041003130007000000c04431000ccdf00c0c4f70c0100c004110010f5d300004140000300303000004030f00f53f00400c0f40c0034303000400300c0c3000f00001110000c431000dc103c700c001d315c030001000d04d440ccd0331000f400d3000014f041f401403c30000040df0f4300311030f0004ff31331430c0cfc0df3d3010000d5004f01443430c00414441cf0730074c00d1300c01400113c3c04300430d140330c441d700f33d3dd7c11000cc0044cd100100113c040001dc033c440001dc000007f000014000030c0f000c10c1f00dc011c0c300003c00300030c00413c1303f500100103d030050dc0303c3041140dc4000074703000047c5403c003430003c030007031400043c007004c30001f5030c0303011414010f04001d130d0f00c0f010c000000c700c033300c70000c0030d00000044d1010d10d31d34c3000350001c0cc0303413130fc03c303403004301c1000c10fc0010cccd03310430100144045f400000000303c70d0000151315303100100c103000d000f0d4000003000f0f3f470344470000cc13040c3c100003c0c03000000010510014043f03300ff4140d05530011cc03000340f11f0d003007300c0f14000301000004c0f04300c4040c0cfcf01f0000ccc5d003004d07000010403033000dc035c000c3d1c3304010004340340104301f1000041403030300000c0000003d3cc0011003000010000003400003d10ccc000f0330330c405c033103030c30040000001007070c03000c00003c3f3010113cc5300300004c0f00d43735550000010c3c3c103704101cfc1003000c37070304d00cc0000c4003001f33d03000004330300004d4000c004ff001040c01000000011c000c30c000000301f00000040000340030c4c415400753030410f4037c340c00c44c40f0005f1c40050000050f1310003305000f0c7d003d000004c30c001143100c17041f4d401000030c4c033011147c04073004000c0d300c30f0000c045dcc1700d001401c4c100c300030473c0407c5c11dc505300c0fc0cc00c0003003f00003cf000f40400735cc5c3700f104c40cd0c35c044c7311003407c0001340000d0004040c0c300501000cc01c7403053c4000401d0440334f00300c14301004050370050c401f000740300;
rom_uints[389] = 8192'hc3000040034001c30000110440040413ff10c0300100c004000d00041d40f40c00d04153c403000fc3000f440000000cf4000c04303040310400000d70000004cc014d0400c430c4c00000cf37000c30000150cc304c03004444c00140000cc001c0c10cc1c00d1044075c0cc7f330dc030c70130700c40c010344fc04010d0c47cc434501000c43000000300140070c0100000300c30cc4c10300044007014443003300004c300c1041010cc134400d0001010000c74ffc03030d3001070104010c00000000ccc000c3070043c0c0c0c0d514c1c000d00cc54001c011cfc30f00d30040c03c030400d0004700d70010000143c14f0100010103c0c30144000c04030c00f3c70f0f010103404dc30003cc744c144043c000453401c7d33103c003cd100043f700c40004031c5c41c3c00f030105c00041c0410c04c4003c00c0cccc040fcc00c4004c0cd07400d30c0c74000400c55c0c00004541033c0f0c0c0000c40d13030000003d0cc400445c3340cc0345443704040c34000cc04c00310cc0c1073f0f00c303c100c003054c11fc00cd3d1000f4f43045040c00d7500df13700000f50cc5d03cf04000070400101000f4d7c34001705c03300c3440340c300070345340c00000d104cc3c00f010d71007c400c1d0f0cf041c3010144cc4f41c00fc17c0c040d4d330041f3030004c00d04310c00c301000404314410017d0c0f4415100100400cc1430334404d7101c540cc0f04cc04cf00c000c0100c0f100d1dc033c4040074c50004c034010d0c0700c30c700000c44500010044734031d340f343040c0101513005430f041070cdc3004c00030cc00003c5414c070f31010f1c4c0f0043c300003003c100c4404f0cc30145000fc00f00cc0340c30400c5c70000000cc31405007003f00ff0dc4f35cc04004f03c004034f00c040434f30314d1cd3340403057c0c7c003f5c4c140c043003c70003040100c0cd05400c450d0000c0000c000511c00c0341c040340cc4c00f4c0500050000c004011100c0c0c403007304453003c0c4104d0300471d0300000c00410f1f000c340f040003d0cf500cd04d00070c01cc44074f4d7c004f0003cc0077010014cf00000004000030301001140c0000d0c4cc000c0c11c4037130000cc40dcf03301c00c4040f050304414403034d013c000c531403070000c4cf414f3c45004fc000c3000d44c30307040cd1400c0c054014cf0c410c40031001df330441c1c04101cccf700000000c0f043cc0c3401000070c35c143c0014c0c00c4c744407c0f0031550000040d0c0dfc00cc0c0c050100300c1f0cc4c3007100ccc04c000c30cf00c0000dc00f7d01c50000f341f3cf00c0c000011c000001cc03f3cc0cc0350c0140000005f070c307470410000300c0047100003313000c00d3c17d4000000003;
rom_uints[390] = 8192'h370140000040c31c0000c3000000350140400000003c000140d030010c0c0d10101cf0004310003003c401cc01000c003c0000300111040000004c003740f3000130055d0003c003030010303c0411000001000f3cc00001f04dc1d030c0400c00000f333c1030003040040370f030cc14100030100030000044c1c034470000313030c00c03c0500001000c00000054000403000033c0000000040003011540500fc011000001335100000000100cc3005c350000047000100000d010c0140cc400400010004000005101330030100cfc0c33013000004c047c0000f0f00c0103300500cc1010000c4000d10030f1400000410f0f0430100000000d007000040c3f30400c0d000000dc0110c0001000d011040000440d30430d305400cf00dc30100c0051010c00000330003c301d001001d0d100110000114c3070000310c140000f010003330015000044d0cd1001053d0000301340401c003c4330010003300f031004441c00d10c100500f330010000c43030c104000400700011c03c30041003414d000000400d3000003010344700c00000004040131433075040704030031c00003c10c000314c110300dcc1001043031c037000000c5030cc3031010dc1350000400030303c04000c0000107000040c000011033003030c00054041103303001400dcd1300010007030340110000101113001000c0300433c3050034cd00c70340100030000500d0000d000c404403c40f003003d40410040003001c01010403cf4401000c0f0c43c0c0000c7304000dc0101c000301cc43d007c40f40011c04cc3110010043c40cf110330c1040100c0101311c0000c301cc100430d1100010414003f30c33d030400113cdc7451c100c030300037f0404c40304330ccf03000000001013c70f03010f410c10c107dd000143d0050330300003c3c403c4010104c400004c0404001305040000033001030c00011405c33100000000300101c00000c0c300000c0000034111000f0d40103c47f0f000c3001001000000010d40d000051000c04c0101030000030003c3cc045003314300470447004dc30401000d40003cc400704004000333d4000301030443000d100cf3310d100c0c000400f00074107d3010300334003730007c330730000100040300004040050401170103cc34000030000140030003c0403c000c04434031c1000304c0cc00c10d114d0040001f3c030401010310000000f0017040500c3000000343c0f04410c14000d000f10c0045034001c44100000330f1000dc000f7c1000dc00000040c000040d0d104011c030041010c0d1001100303000301c007000001110444c001df0100cf051440130300000f30004030017c4000400c30c07c0034f500014000410000dd43004c0d03c0070f0403101050030304011c35033103c10000000;
rom_uints[391] = 8192'h514cf310d300f30170c3000313010f001f00100c40000c0333710400f34310000341c03430000000410c00403300000d130d131070033c0c430003d000030100c300003dc30c0000cf00073f0113c330c33004033f7033114040d00017c0301001c331730000013310c01041004130317051c3000c000310c03343043c3704007fc0d0c0034000710030c0c1010140d01014c03000f3300cd04330033040f0c5dc003003031013c07c0101030130330043d000c30000d0400300004111000c030dd0330d0030fc73003c004353140c00004041c300d070150047d03401300030c10c03334300010f0043400f4f033d030044400001d4000f11037003c0070000c0f77000130340d040375574d131034330cc3003d01013030740047f30c07f43000d4d0000cc01035301031d1001cf004313f13011034d33000010c00fd04104c03004053c3010001c307003c05d0f000c03f1f0001dc0fc70cdc107ff5cf301000130317400330041d30000000404110450dc005310d0f0c313f3c40311d704d0000c0314c0301003c3004005c04cd03c00000000100303d3713041301c401004007001c303300c001f000c10c105f01000ccc0f303d0f3c0c01cc100114003303f3030000c03cf30f1330030000300c00400c100010043007340c303010330130000300403004d04c0030c043f0133510000cf4733530cc010000013110013d13f00c71d4dc1017110030001000100000000033300100c100f1013c433f3104011c1004c0000110011f00433001300411c04c040cf4441d11070030740c3c55011ccf0303c00c001017c4d3340c10301330000001f4c0000d515cc41031104430d0c30fc40731003400310330100370d1301c0c330d7f0310cf310f01300f043d0cc33c000734051051335010c004430400d004cc0110333c331003d3000c343330c0cc0130041d0c07141f1c3503c00d100c100000c4c3c40730343734013100300c300000001030040c00034530301011c01c1f03311035000304103070001000001c3034c0100000f300f00010113001041033051000303c003410043400303d300333c30c10110005c000040000010300130714310cf7130c0f40003500ff03000003010030300410300c01030000004cf5040430341000003d3df43004303f3011c40100003f00100f01010c033d0001700c000c143c3100c00f300cf33030033ccc7004ccd44000c41c3103c50100010ccc01d000f5000c1131311504000510333003040c1070010413330030010c1103045057000c1101041f3000dd0c300403fc400130000d37010000c00007f13030140134330030000c00f034300400103c310f0d000030c03030000030100f13000000031f010503175370300101011000c33100f110343440cd033c0f7c0003073447c30030031f300000000;
rom_uints[392] = 8192'h33300c000013030fd10110cfd0000754f0034170000110000d000004c004f050404c7314170000c3c1300003c153c013f040340040f11cf0030311c13300304503c414450001050040007011300f07000033333141d0100f7013040003c3100000d10103000c07403030c00074f303f0c0c40044000c007030001c35353c0005005d0c0c43f0011000301700005f4dc140c0050000c000130401c0c0010d140000040103031f005447c10340017f3070403310c0010f00300370043731700173f000001d010c53c0c0f0dc000f3004004c4c54034355f44040f0043c70f3001d0c0000300430144030f001710700c4c000773400410c0407cc0404470000c0013010d10043001c0fd0f3c01001c00735cdc0c0340c040700430c0f01c1f30dc0503000033f440dc330c1c0c030407344c30c0157c041f00134f7c144c104c1434003f30c01f750043cc30d0c3001c05c003150d70010f0d30c717330070d301001700c01514031300f13c30f00430003df013005410f311001dc43c0300c11337003074407d000fc433300f4411cc131c00103130004340d4151410f07c101c4f40c4c4c33070d10c301300f305f0d3c11003f0400307c04030430000003d00014f4c10c007c0f0d000001100c010103314000c0330033c0453707001c001d0030004d000130c1c04d3c3300440d00c000c0430c00c300d04000050333f43fc0110f03d14c0040071433f30cc7315ddd010d0030000cc37cf4d1c0f034334ff0d311cc00004c000000c1350c40000c01cd0143303000073007014143f400007035cd043001007400cfcc304c3d3440000010c003c000000307403cf41d3000f001134000c40000030000c1d10c130075013301c4c530f030dd3c4403d304c370400d0410c1003004014170310075043c030000000040c000304c400c0074430c3315070310130c0f000550cd0307040f500d7041500001d030c1301004c10cc7000307330007000c0000300c00014350c300c43404f5015c14c030100030010010017700330d370000114c00c0cd04000f700c000004c4010d00130510c071c3300cc5330100001dc0310cc00c00400d3f00c30510450dd031d011010000c70c443003540000c00400c37c01000311c0cc10101007c40303d100c310417c0010013c3105134c00100143c10c133030113003130d01f0013c00cd000700017050f00111304000011d14f000003037cf00cc3013f7300fc00c040001440000c000c1475000300c40c01001cc35000107503c7c5cc004c010c07344fc04003004c4000000070c40104c030c5031140ccc000471c40330130000037000000f441f01c30000d304c701540fc070c0440c0cc150011107f40004d04c70f010147c010d01047c031d0331301137430c00770000410cc4000000310344c4d010010c301;
rom_uints[393] = 8192'h33030000010000050f01cc0cc3c013700c130411030000c000f01001731704030c34f40cd51d00334c400c014c0000c4c30f30c740cc0c1404c000c41000410400000105033043c3040000004dfc3c0c3001d540f17c00c40340c15c00dc3107004300cc03003f433303d0c00071c3000105010d0d01303000d1dfc0401cf0005100f41003000c01c0700301500c010734010141000c000c0011030c304d10cc3c0443070105400c04500433500f034340c3c0c0001100010403005d0300c00cc3c0ccc0c000c3110f0004c103014c001303c10343005001f7f010c0001d430030c0000c4c404c43cd300153414371df0041000d03f00c0000034444370c001c0f110c073f7004333101c40d410030c4fdc407400c34c300f0c3c1d311d15c00000ccc00c3474310f00440c0c7037500c3300cc301140100130c04c0c033013cfc7301c103cf1c00344c013d30070307104c401cc00103c501c00c3c0441010c0c0c3100330f04415000000f0001f10100414000400040d00013fc054040c4030100d403c0cd41c0444107d005000ccf4000004000003c00f0c030f3c0f0d40011330400030000030300d00c03c04dc401000cf1103c003007100304401140433041000c0033003c3cc30f0c400d500337f0040f00c014c1004c0000005741730ccf704034300050004050407f4401404d0000c7104c044cd301440cc4c507c344c003f30c0c0c3151c41300c1074d3cf3c3f004c73c0103030437f1c10f0f04400130c71003cfc40000df40cc11000cc0c0f0003cf07d0001040c0c4000ccc44515f40f001f03000110703500540cc30001c300043c0f034d73c5d0c04c00cf0cd7004030000003030f43140001c0cc4000d14c00c3f00110004c00c100103f0543113007303c3c403df03c3f3011cf50310007ccc30010001cc3000c0000d4774503c4cf00c30330dff040c10f04101cf1000050740011100007c3040000c1100c4400000013c3c300030003c5000c43c0c05dd03141f03300130300000030f0000001100c4031000c01010450041f4c7043d10c03c0040d103c0cc05cc0001740010770cc03c54d04401000040330c000000f100040c0430f3000cd4100501710003000c0c4d0005d00c0d45015100710c004071d400304110c0307030450007330450f4cc00c0003cf0ccf041c4d0400034f00c300033c00d0000147f31c100050d300c00037f00c00c44000f0033d30d30401c1ff00033400f0403000c40100350040007d00f00c0f0130c0c313030000300c1d300030f05c0100431033f300000c43033330104003000df000040010d3017300010044004000cc0417370c03f3130434d3c0000043dff30c000c0710c010000100400c0140003143001000030000f00f00000141104d0100c300000000017444430f041c110cd7003000;
rom_uints[394] = 8192'hc000750307370c0cc03c30101f003454030400130410d00000370050005c50c0c3431c414fc140ccc01300500000d114f340c07070cc3c43500014301d1350001ffc004ffc0300c4000030041440c0c000300c07174dc40cc3537c010c340f3100f000ccc3000431d100034f10141c350c54cc3cc0300c5c00100031440cf0001001f3cc14c130031c71034c01007343040d010000d00500011c1c10100314050000050004f000070c303000f00103c10c3c00f10004c0500300f001f10c0343554c3cc70c0f7330c05cd0f0c4f047d0c03417ccfcc1d11cccc53c010dc50c4c77431000c1c000004034401d4001c47040d70330fc70001330d3fc3f0301314f1300140011c003c0303070df355c0043571304ff03c030c100c0000444013cc010f53000331f00130340100c3cf04c01cc003104d01000000f0d3100f0fd30c000010403115d1400cc50c041fc010fc5531c040c33110c17037011f1cc070300005c01c3031c30cc500047c107105377001707f003c1cc5113ccd3031000f101f047c33f30300d430c01033050c55301c4000040010001000d1441014000434f10c31403c3330400305c030c31c00503300c4074ccc500143440df704437400dc10c131070c0141c3010f340cf1000f1001013c0031cf34c415404403003c4d37d30040ddc034044000f4310d103c3530300041f3f00c00013c30434403c34c47400000d10410100501d3ff3403d404dc10004f00c3d0ccc0f0003101d100040c5f0373510000010c0001100001140004073001030030cc04043331004303140c041500000c0c0010400303f4f5f00d70001013c5f40334c051330005403fc00c1140f0dc03007c00f441c3410173c0011c043331000053c44ff0000347f130f107134100d3f101c4c00dc14f5c447f010cc534003df03100cf403300c0ff1000c1710cf001003010cc0107f3400005310451f0400001c10330053d030c400d01410000c0f00100050cc0001001f30c4134cf30c07001010f10030754430f3d0400040500f00100fc0041cc03040404530000f10100113000334c03c50430d1133130f100c044000f1400403500c03171f004c414c0f05c50400c07311113054f140000304334c0401c5c0001033c341f00401340f541040740403d750c3c3000c014314d4303c110000f04104001c0000001030c0c10cfdd333401300001307014c701003cf001757f1045300c007003430f4130030377070ddc030c0c100400c0014c043301c0000f00c3c1000c0000f0d041500010d00fc00c500013000010c71010f003053c7730c3c01550001c0300340500d41034310f14300303004000c3f010f3033300740351434d30570f1000034100c1d30c0037370000d00c0f000c400030701c03c04f1031dc0013303cd0040000000000143043003c1100041;
rom_uints[395] = 8192'h431041000f000431c00000c400c3040000414400cd0043400c0c0cc4c0c000574057c5c10f010004c710c40010000300cc4fcc330c304dc00cc1c400c0c00400c1033f400c444c440003ccc101040004c3c00510111d00f04f43c05c0cc13c00c1dc0c0040040c000f4d0000010c40c70dc01303cd0041010300c00c0f5700055340c0c0000c0c000c4400cc0303400cc10c00000d03c0003f0004cfc04d014c00c0000104c10c1f40c0010000c40f30000d30c0000104000041043dc0000001fd030043000c400ccc004f00cc0c4fc0400340000c470c007000cdddcff00700c3d00f00cc40000004030fc00c310300300f43044d000047040043000f05c00f3c03430f04004033c0cccc00f000030d0fc0130101fccc0f07c0c344030035004cc7000c0051fd4301430104700540c0cd403141030c10040340c04401c0cf0040cc0d05c3dc000d00c30340454430040000540303304104730c3c50c0c1c0d04c3cc10f4341f007fd010d0c407dc4c30500034744cc731103c40f000005c05dccc0500cccc00100cc0c030040013cff0000c0c0c00d0f00d443405ccf3fc0c1c44d0c400003c04030404c3c4f14f4cc304001f3cd0c0fcc000540ccc4c14dc0c03000c4c041c04f4cc0dc0000f00c4c0cc4c000110f400c300c010d00000000000037c03400f14c30f1cc0cc434000c0d00c013c30c010000730050f033007cc503330c054c73f0cd0c03004c434000c04f01f040037440404710d1cd0c1c000c31f1c40d400470ccc4c00cc0c1100ccc1df0400c0c0c3c0d33430100c30c00c5c4434003c5040df4c04030c0574fd0c0010303cd370011cc004cc00cc100c0410c0701570041130f0c04c30d04cf05434407cfc7c0c330c0030030c707544000c1c0040c4c41400f0c71c04cc1c000ccf010740c4d0440c0400044033f30c1c440000000034000410443ccc04cc4300d010c444d1c044013c0004dc00040730f4c4f00000000f0c0000000440040004301c00107300f4c3df33c0000f30403000301f000c1404f0d00300000030c0c007405430370410f03cd0005443300000ccc430050040d10c0411c300300440043c0000c174441040470004c00000d30c3f14000d00010c4c0cc000cc344101003dd0cc110034041fc0000d00030f03440ccc040440c00004400134ddcc04000c0f14cc100d30040304cc70cc3f3701000c34300001000cc40000c14c0ccc0fcc00c0cc03074c3c1f300003f0003014ccc0c400fc007c101344c003c0cc71040c04d40004cd0cf0c1c0cc071c04040c031cdf3030cc30dd04d0c04cd4403c110c00c10c0d00dc100004cf004000c10044404c3c0cdcfc31347cc37c551d0010040c5000c00410d034d04c0004040030cc000000c54f03fc00c000cf103004540f00000040000c1301000c00000c4040;
rom_uints[396] = 8192'h100001030d40030400c30c41c0037dd104000c3050037703c4c00057c73c030710100007040030300f0003ff0300030100100c434000f305000c00c0000303500043001000001030004110131000dc00100d0113141c001731fc33040c0100304c00c73f001330034351004040333f40400cd03041000d301000100cc000031334f3f0310030d000f0001c7f00010c3004400c00100000f03313dc0403004140703dc03c4170c000c0cd0c50f30300304700300010400030030433705330135004401100c33034030000070400000c0c0034f1c3300340400d01000007400113000044c0413043003100374f0011f40c00f01000000000c00000373700001d070000c31300115030f000543140300c033541f004014d0014f00030c00430501310c000304f00c300c043000000100fc10400030cf30000010430340d0003030540700010030c000303134037003170043350000c530d5170cd1c000171c51d00141c01cc1010000130c01010430c04301341c0c7314000f10f53c043004d00f00004f1104c3c04f300000310101330c000300f01000c433113cf1c07740010f15d01c000f303f10031c7070741f33300015433031c130331c000030c0c000403fd03003403033003400030000011f1305f3c370450d0003000400141f3310cf0f3000000007050c0c0000730400040130407100040f10c5070331000311111c00140c37050304300040000d0000000001045c5030030101341d001cc0140003d300101c3dcc50003f01003030000c003cd0300d0c10c130301001333000c13301c11000300334331cc4740c43301000433351000301300c050034f51030c044005030d53001003300c3034134014030f1035301cc040030001c0003300f05d50f1010c03d00003000cc7030300c0341c104c03c007000300c053d01053000cc011505010117533701c51f0140001004340d110007c4010300457c341f50cd3cc00033001000110040007034c011000430000f0300d30c01300c7000fccc4c34400d031c30043c040751043004030000311017c7003c400c000400101cc30103c1000004d317001c701013033c7100d300400f00d000040010354030c403301ccc34330d01101003cfc10010100400000100ccc003c30304dc0304dc5010000c40f3d01403c3055330001003c031030075011c3c03cc00c5c30f3005040d30c300043001010030400c01001c001011011010df0344100c53c1c0010c114c0317c3c5c03c300dc003130430f0400cf05031f014003fd4000c00d30013c07c007c13c37c004101070303000000030313c00004000c110d0300000000041317403c113433000c3433133c11cfcdc431300070001100330034310f3dd0000f1401303000003c3f3501301c30c0000c51330f3c0500001440301300c301304003030;
rom_uints[397] = 8192'hd1100040300000c0c0000313003341c0030000cf40c00001c33300c343d000410000c0000001c0044310100000004d00c040031030c01f000030015000100000005003033000c0000070f3d140c0510c33c001ddc05100c0000043400c410000d300033000c0013330400001000400017000401011c00031d030440fc4001cd070000003000041000c0140430410f43c030033000dc0c04cc3c0000303030003134503404141c000c3000cc3000041014c433000c001001370334c510c000003c00300000003c0000311001410130101c0c01000470000111100400310c00001140003c0d000000000000cc343f1c000f01d010033015000001040c1300003c033434400d1014c4000c741400001c0303041c344c3c0004011001d0000f000010030001101000003c300434040114000c303f00010000030c043003304104400c0f0330034500000c0000000300171c0c000c10f00430c71034300004000001133303040303313034c3000003c1030000c10010351300003000000100070004c434313434011c04103300300000313c1003000c000440007001c1103f400004443000340c3000f0cd0c0f300370300f0003040034000c0400000410010d143c311c100001000cd000333003300c0400010030010d030400033504033301ffc00c0c0c0071043c300c300c003dcc0c000c003704003000003000001000040fc03004007100c0303c0c73c00c34100003000030503d0c040ff0dc100c3c300c000f071030000435000c04000000310030003031100cf10f000c00c033000c3070340c1000000000003c01d000dc34003d003c00000035c00003001f371100310c0cd3000f44000410001f0010100010011d003c373cc1030f03c73003300010000410c10100c0003c030110001c30c40c3404301d1000000000100001400c343c31dc30303433033033c0000c301010300003000030311c00300300100013030400000014000030000030000003110400000c0c000000003f003034130c0d000c000cc03ccc010000030100000000000c0000040000301003303033001031100033005410003f1000000000300100050010000037000103000410141c0000100401031001040c00000c70130c3005000110043d0300010c104000040c3000070c100330113000000011000000370400001c30300033400404003c0c000c0cff30c0000034c000010c34000c30300c3000300c00300c000304340c00000101000c100001000000dc037040010c3101101f0cc01d103400000730003c04c0000c0104f301030000010000000000303000000405040500003330000430000000000034300c1401703030c03103000410000000003c0c011c0414000c0c0010300501310030030c3c0dc03c003033c400011c3030f51000140015101430313033000;
rom_uints[398] = 8192'hc340c4000c1c3c0000f04000c030c30330010030334440300030140007c440c000130c53f03000300003004000040f041cc40c500000c413004000040400d030000c30307003c340c300704cc300c000c0d03c10c44334c0f47040133c43040c300107000304c30000c4405c04500fc004cc0013140030000001101030c034c0770c004c33f4005000300010d0c07cc0c00000700004700100000034005c313030404c0410c0000400040dc3104330c341310d3000040c1330c30c10c4c40c00c301001d1c00704c047000c3c413c0330c004133c00004d004f000f50f300c30004001004054400c004300cc07440034f0434413c01000000000433c014000c0c3000031c33040d0000000471040300005f0000000000f07030c1f1710dc4dd4c044000005c0c014101303500131d10000000400033000300001c400070030001300c050375410c000f0013c330c0d0431f0043400031311c50ccf07004000010300c000f34001c4031000001c00dc5c00040400050050003c14471f43f00c0403040c00d4100730c0c000000303c00334004f30030030004300007000104104040f01000fc0000c000000000f40100c4100c0000004c0300110c030d3df07304033410c30344001030351c00000001003c004c0013030003000310000313441d400400134cccc13c037d100037c00404005447c3033010000030004d00cc0530301001cc40c0001000000fc13c4500000f41130035014cc0430400013403c00051c4100443c00c4001040404f00c03c1000000343dc0c40c04cd00f000004101010000000c004c001d101c0433000040f05f300370130ccf04cc0003d331c44030100c0333000c343403004340000c3c0c000100c00440c0010c10011400000c30051000000000c100000d313331034dcc0c3311034c15000c40400000d003040040f031c0cf040103cc14d3c430071101000003003034730004140000300cc30031cc400005c00730c007000cc4400000c50f050dc73101c0004040030750c010030140f1000440c004f40005041c003c40cc0007000004f0500501100000004101cc007c00000030007100cf00301fc0000000000400c001c30c0000010d0400000001041c000744ccc34000404050001400000040410c001017300c00c01043300000300400030005300343c0000000003430000030cd4d407014300003743000330331004300003000540004100c000401010c00c403c00000c00105000d030430403031c00c1f443000f30c4c0c4c00cd4c0d01000435000001c3407000000d5c43c0413d0100040c0c000000f004000301c000c01000000001000f4c0400300130000c0c00001cd1104f4400100100104404700fccc00c0c1403001400004f030744000045c300c0000033cc07cc00cc000c0c4100004000c04c40030;
rom_uints[399] = 8192'h130dc13030c00030404c0000cc00c305c414005000041c0f00330040c04c001000c140030535100030011030000004104101d0134304c7030d0310fc3c00007000c014f005040403040010c14c000114100430100c3cd43473f0034c000010500450c010100c40034100c40050cc001330010014c45f044c40c33c0030c53d3cfcc01003d14140c400fcc07c5c000370011051000040503c0f1c4c1104345d04010700300007110530d7033030d1411000700044000f0f3c100300405434fc0c401040f10000c40003cc101c1410c0003450300740401f0154504750330f40005031400f0000c0003f4cc0033cd73f000c4401cf435003300031c0003c1040011c1010341400300c741f04c5f30110c03c1310d054541c40c073c010c3301c300007c000403c10d0c43cdf034034ccc0003d030cc434000003c0d431c500c017c50f4000000cc030c000c0003f0030004f0dcc0dccc4003d144c541007c7100410314df0d50d30303010c4d3c04d4004403fc40c3033003014540100303054003310c1c55404104c1740000c33070004300010cd000010041405f030c0f105c133150011133004170c04030757004c4000001dfc5c151401700df400dd0c4f10cc034701030f0400c4d0c400030003333041100c3c50c30c000004c01043040cf013c014144040f341cd4c000430004cf410c3f740c000f1013f07107004cfc41110134004f0144c303003043010c00050f0410005c03701c305f0c3740c073c3034c70fdfd0101000c71c0000704c3030c0d04cc0d31cf035c400c15c074c4cc0730cc33033401004307f300f1f3400015014c4c001d70343c0307001030413c00430f04705c70c01fdcd170c00c400010c0f303031000fc00301311007fc3000c0cf1cf0c00f1330014341dc0133150d010170304140cc0300000030003057d0cffcf401110040d41001fc4340153f11700101003340c004043dc000000cc1c4c100c00300c04c4c000c10001403500c04300300f0c0c01040013071c03f00c000cc30dcc300310014c1000c3c030d0c1003730f0f04410c1c34033ccf1370fd41301001c0c1740f0000003074c0fc73513c00f0c41344d0f300c35030001053cc000100c40000c40310003c00c400070c4103040d00cc070000141d0c4404001cd0c0c5100101131c4000d0340c007075000010170330153c010c3031c1d500c00010d4050330705033cc40f033c0304005300010c3d0d30000071440c073030404c00f00c0000c1033c0001000cd7c7c431ccdf00000c004001d3000400000030cc4f4103c1cc30fc00140fc030000f7100cf3005d0400001400cc03407c0050404df5450cc4ccc000401100c0400101c4c040000d4c134040c1301550434003c0003043430fc3130f404070000c5104c0010444f03fc00144dfd0070000;
rom_uints[400] = 8192'h340000004341c00300f1000c3700001141c40cc004030010300d30003c04700400100c1ccf000004f331c000c7300cf44000030c004c00c400300101ff00000c0c04c30f001f000d00003c30700004f400c00c34c00400300040030000000000074413c000000000400c0c4300fc0fc0400003cc300c0033001031dc0c51700043303f0000003133f000003c3d1000c00000000c0000050f0350011ccc04015f0303440034300c000337f003c40000100004fc00001044c0104c00340743000cc00030c000001f4000044000d014f01704700c010140c7000117c3001c0440101d4f0c110004000030d30044f3dff01d00404030c3000c3001c1010cf10c000c0330001043030c00000400ff353c310000c40414000703013d003110f7000337400f0000410100000c0304030430cd330c000c010f35cd03000033443f000000f000000303c1000000001dc03004400400000c500cc03000c4f5034c0d34003c410c03f0431037000311cf04053c0cc30c00007110c1010c00054c007004340033fcc0004c0030000300000c433c100cf500310c30004100005dcc0000040000010f4c011030000c0c001c0f00ccf001343304f4010300c30c003c01c0007100dc04030f0c01034510001000d3003c31751c0c30050f3c4f3cc73c000d3500f10000cc340000c00f313030000c000000300404014d103030c400004c340c0030c0c0004f1c0c4d030c0300040d0c0c0030300301100df30f0c14c5c4c04c00043430f00000430003c04fc040000000c0040f0c4003c0443c0440010034000d1c3433c0cc031cc00c333f3c300fc03f4c3430005cc004d31c0731f03040440400044c0c4dcc1c1c340430100d310000100f0cd0030c300c0cc7013303cc0f740c00c4c0007000000300014100f400f1170f331431011030010cc15c00000035000475703c0100c00c04074c00cc0d3cc14cc30fcc0003400cc1c00030030000001070050001000c3040c0000000000001030c010c3f0300003c3300000c4344000f000334c0030070c00f000300030444000003044c101c044c01000045f030c371000047400c0030c00100c000000c0c100d000c000c4400040c03c04003c14305c30107341c303300f01c0c0000c400c00c00100040004137c0c000300000c3d0040d3000100043000c41001c040c0c05003037f4100c0c30c013300c300c0013013cc4300c0c310007000000007c0f33310f300c0cc710c300000c003c0030330c4013cc00033030140003400d0540f0014c00701d0300034730003f100c0070c0301000c40c050c04010400300330000314cd430330ff400005000104140140034cc100000c0103000c0d1cd000104c140c0340410404d40300000041c00134000c00003c001f3c0400c30cf01031041c3000100033c7000d010040100000;
rom_uints[401] = 8192'hc001c100d5c4000300013300c0001110f01000013040550c00400d01f3f00700c0c4c0404f0c370d34f0010cc0c374c010337340000000f0100000c03d1ff103f001ffc30074004504004011cd00c10400401155c1c003fcc3c0f43d0c40174100c30c0c00000d001001dd0431405040340010000400c443000d0073cd00500cd00cc700044100000d04c0c0000053000d014030000000c04103d0cc3d001040c00003004003c4d53f0004000d0d0c7000030f45000ccc400003c0341000c034744043c0c500c07004cd04431f51c131ffc04c030cd1001c40cc014003704010000000400301dcc0030700fc734303c1000300330c0304c001030000030000c33053100c400c1304c0050f10c40f0300c0c00dc000034400530000014341c003c00f00001417404100c1c304c03300031403c003ccf10c30c0f030030011ccc0cd404304000041010d0c00003301010003c7c00c13f101133431c0411000700000000047ffc5c3ccc304d000c00c111040f4000403c4053305010d00000010c50013d50405d10cc0305401401d0cf0c0dd0001c30000100100c4000151401500014004c0030f000400000003c0113130031000c0074dd0045703c00030c10c401004f003000301f13000c0331374004045510500c04c07c001cc001040c40cf00c0350c030cc3f43c3f704c35f3c3300f330c011070d00c051440c000f0000440ff000101030c07cc30df3d330f1c10d3f14034030f711c0f00cd1d04d3450100071f040cf00500000c07100c14000f000c50f0000c30770037ccc3d5f031000403010000c00044014c0f3c3f0c0c3100307413001c3f10cc030000040000143301c0333dc3000103003c444c000c00ffc0c17c140305001cc00d3031c04c10113c44007c0c037400301030cc00000107113f40ff31310c100cf0000cdf0f04310c03333444c0031c0015cc4400f30c0cd0015c31c333cc0c50030550011000313000c30c00000034440003c00104c1430c4d14f1430ddf055000c1c0301cd000f00c005c310f3c030d0015004430030773004c0c00300000010030000c33c001500100710c4c0c030001100010c00f4cf331c001000c00403c0404c10010500c4fc00cc0cd1d110003443404044c04003c033c000f400001340c0041c070000cc0005f3cc04055c00c00440c1c0000000c0010c4031003103f704003dc3f3d041000f0c0c41c0c10043105100d03040d3c740c4c070c004f000003c305011110103cdcdf170030000c131ccf01310004004001fc100c103c0007003013c0331004043c004001010004005f110ccf10100cc0c033d0000c340000300c1c411130303f000c1c3c1ccc0000004c000c00100fc00c103730047410031c340d74005c01cc0430703f00c0000c40000cc330040000401430fcf37d00000c000030000;
rom_uints[402] = 8192'h500003c0c1d00000701dc000000c1400000010401340c00f000040f30c70000d1040cc75f0300d0d1c40000f300f35130013400401c1c3cc0030c100003c4c001c304443440c0700011f147000cc004100c3ccc70c03011cf00130000010ccd1417004700c1133300d03547140404c0c54dc5413747440cc30cf300110000040334100031007d000300cc30c0303ccd0c040c0000f10c0f003c10f41004330f340f000cc54f0003cccc01d3f0404cf0c30f1c000000143107000c41d101100137101c003010000d0f440400001f0400051307470c00c040c1070507d3000f041003010400001040c5034fc40310033c4070d00400010051010000034c00dc341c1fc01100c003030000004c440100c0f3fdcc41010014d303fd74c41cdf4c130f0c000c043330000001340301cfc00d3040c001001100d040010c10041f0011300c4cc0170f00c730c05003c00130c040030c40d30004c130040411f0330c401701fd35710040cc0140330fc304f7330fc30011f503001171140c31c1c00c7dc5103c4c4c0dc7cc4cc00cc030d140010033d7cc00001c111000c0cc0001101f01f103c0c50f03130f400f03034d3300001c30300d10ff41c00133103f4343f00f45c14300c37044000f00c1c0c34cc01500cc01c0401d00010d0300330000407000310001c10000f0c30c040501000430ffc01f000c00c70000000c0005040000c34c3703403010030ffc1c03c704c017d10cf503010010f01041141f040130331cc4430433c00000d750c10034c00000c0401110430000f4000000100dd000104404001d310c0d403c0c37c00000000c13000040c43400c4c1030c3c0dc05100000f04ccc401700000000c0c03000c313c0000000c00c1c0cc00cc103010110f30c000c00000c07c54f5c0301f01101101000030c353004300001f0110c07c70044100c40030c00d00301040030c533d0400c03f471401d00f1fc74d04140010030330007fc004003304010545000050410c0cd0050011c00f430704030fc400000010000431c105c0040400300d4f0100f01c0500001404f003333f43000010c000014c00c03300c5d000330011040c000010034100cc00000f0d0cc00c400300010d1005000033550cc01dc00004303430f0100304c1c0fcf0730334cc4c0c00330c100404007070035f00400fc733344731140c00ddc075005ffc0100304003d0c01704000340c1f0440043004000074c7d70c1c0d0c001044751411007c1c70c1700d0140070030f730304d000007030007d004044310f00c303045040f0c00443c30030030013cf4000403f001300dc03004c0004004d000c43f40000c40f411f4147d4030c014c11100300c4111d0403304001d0000403f07001100000c400137070d43fc3410cfc43f1003300f41400f110ff070c00000005004c;
rom_uints[403] = 8192'h3c000c500c00c00c103c00000d00301543150001d0c4003430030303f004cc000010f174d0100c040f01c0471004401c0f553003f41300d144f31c0c03c13104fc4f10c000c01d0c430004100c100ccc113030013004030300c407dc000340001fcc740000d004c0013075cc0c0c3ccc0c4053001cccf10d003000c571001030cc310004c0100314c000003c40010c00005c0104003000301170f5000030c0101110001000104cd0c11314c00004303071c0c10000c0f00c103400c3d30304040145304d0410c437d33c305001c10d1f07370c303100040d040d0704370cf0c1110000001cc00000003000c1c3030c00c001400f10300c010304011430300300c3003110f1000ccc1403031c3400004313c1c014541c3c0410043000df334cdfc0070300c0c13c0050330fc0f40440dc3010033303000c04003cc7ccd40010d4003300301f040000c40cc4543c3c00003171df030c4d044c13044430135700043030cd104c4700f7004040c430c00dc0f00f0000c004c1c750437133f4041011130f4054045f533c7700003010000c00c400340033000c01001101d0403007d001037001c3cc0313301004303010f004ccfc5003100fc0301031d3044c00f04f10fcf0040110070104c4400004000d10340100d00043011d001f574304f10001c004cc01140c3301c1c7cd4c01f101343300c040004000700410d00c0000c10c000037c0040d44301c3cf0730c045411c05400005401030000040d4070371d700f0304000c0c43d3001001004000d00134cc0c0043474000103344103003140414d031110003d0404700f41f000d0000300104c001143d005cc303f17c30030330140004011444fc000300143530100703145000000c003c000010c00331d0700d370c10f10000ccf47435c0cf104c14cd1c11304c0000cd00000410c5f0040071cf0c1000044303004010303001347035434017c000cc10000004000c130f015c0c0000000077003c0c34c300004300cc0040c330000710003004131003f0053c0003103410cd1c005c000f00fd44300cc1004130c0140f0310d071010030340c000101015704d43040101c0d14c0f00101d7000f3701f000cdd04301c0003d0133000cc30d0030d33c30d00100130010c1043f333cf00c00705400303004500000540c144c404f3100000cd501010031043003d1fc000070df53c1d001570130440cc0145100c437070400100033300c00d4c1134c0f753ccf40034000c300ff07c5033000c000101c00f5007000f000cc010d0f54403003031000004400f04313cc4340041014cc0c01c103cf0010005f003134000c00c1c104000c110430000ff5400400fd04c005330101d004701410040c3000133c0050ccc01004005510cc00003c110d1430f00310047f033100400c1304311c310000147311000500;
rom_uints[404] = 8192'hf145303cd1d40d031dc00300f35040dcc340d51150040100000000003f4cc004103034003c4d0c30dc01c03015c0001d3f7304f000044344f303fdc0733c300300103543133411c10100c10c5004000101000411105001044007dc10d03030c0000f403cf7300530030075033441f41014013040310004300030c1c41715013c0033c0043131007d0303003c74043c00000c0003000001cf10c03003c01ccc3430015cf4dc0543fd00d33c1000f10f05500f3c0000000300010400513573334301003cf0170004c0303f0000711503c30331043000c0100435350431341d30003000033010c0c4003f0310330fc00400c0175c0f33d400c0c030f4c3011000c03c1010110041101c1cd50c0c100f1133000c1cd0004030001107007100c01f1030150c0040c1ccd101041074000003403c03f70ff400001001070513040000c40310100001d7cc0003400c0140504444733f0001c014f3004145300cf01c410743033044f40f1c1007c0f4333010d000101307141330140040333c110003310cf0007c000730014f003c47d4c430703030011001c00000f004341347510c31000d3d0030c33c1c7700c700701030d33014c00c50fc5300173100000cf030073c0c0c4fc1000f004004f070000c0030c004f3304c0f303cfc30dcf1033c0cdd1fc37c11010c053100004d30430031303005cc3003cf1c0037001511011000010030313007f43f00cd00301c0f00fcc30000300c50f1034070034033333003000f530430c0c07504cc00003450c0000c1013f00301007350003c0030031f003c01140c03040d00111c41c010707050c0001c010c04010000000c770c00cc11047000350cdc0450044d00c0f0000c0040d43c00fc301c00c4035c0000c001f00c070350fc010f00c0c31440100c1c710c053f0fc1d030f0100310c4c40043033c3013400c3c04d33400307034107c0100fcc33000400331343001030fd00410401cc1f0d0000300c0f073cf000341004001100c34d0030f01f000000cdc00405f05070003303330000311cd0070307c00cc4f00373dcfccc400c0c4c010c13400071c03d34400300501d13005d3c00407fff30cf000cf300110004400333010150401c000133130004c005004100310001004d07d0f304317c001dd0dc00c3f03cc0014cc0c300000000f3143003000c0000073003f41d50304013c70310573333111c000110000000cf01001fc333043033cc334c3004400133330003100303c301330350c47000f0071d55013074004c00000174dc0dcc040333431fc0011004f34100c04031300057710c0473c00100c0043100030000c000f0400000040313c0000007000700331000c00003731c3000000313ccc30007104440c310100ccc00040f0003c4000c34410f0000033050041c40c0004003c035c10000c0f044000;
rom_uints[405] = 8192'hff1f0f00414400cccc1000f0370c4004c0000000500113000c30150d305f0c404007ddfdf3503100300f0c3d4350cc43071000c150540733044c4333f130500c3c44330700000400000041c01500f3c0000c45000f03400000033cf4c01107c04000d10013000c0310143300c0cd110c0cc35005534003cc000c401dc4c10100cf300701405c033411c3c301dc00c30d0004010000c103c4c0c113c0010014d1043d41c04134030043070700001c1f310150330100c0030d00040c4d4d000303113004c304000330cc000f010f4037300013f5040141cc013034101540ccc40050410000030f00c40d03005101114fd0014dff00c174000300004cd0430100f11101004141cc3000305dc000443d00000353040344051000057c0d5c3315000015431300331003510030047403000301cc01101700413000040c4c1754d00c4c37dd0d11c0fc010043000c350cccc03c47030040500700f70300c1051073c733301415177c030303000400c01001c503107d3007c37f04c040cc0544034005cc0c00030c050500f0001103507d0043370f000103000003c04107030051c000003d5040041c04001700001310f3c4410c000000430000c450c04f037c40000011f00dcd0c33134c3300100000c300f0044d0103100301d31f000f403c0404314301001cc00010c00034034c0f00fcc00430c04cf00330000000c0c0c0c0cd31031107500d4000000130f0c33cd40404f00715c40cdccc3153f37cc3304130f500434d53c40c43444300030110c04101cc0031c400c0174040c03143c37400c10043c030c3c0400c1104000c130c444001300c1d0c014730040000c0100c4444ddd400044ccc4f00cc00000004100103700d33c04014cd10dd4300530044c00310300c01c30c1000c003c1040100dc0d4f3404570c0f10c03310401000f303c5440373034303c07c11c010d503d00003cc1401c71310401c00504153c400010cc400c3d0030000041c1df3001003f0007c0037d0d040010c35d30c5040cc40c300c300034d100000500015033c1d0037c40030105103d0000ccc0301010400c0301000000050170c7540000000f04107c3503000007043c01540073d0441c1100307c000004300300113514444c1404f0c0140c45d0c4f0c04c311034500100001c000c0f010f370500ccf37c0174cc0c50000140c50cf00f10713dc000c03d0c0017c150150111003114031004104c70000030534400007c0044000dc3001cc4cf300431c5d003340134003f000100cfc100005005300000304f11cc4345c00301045c000c314c4700430cc40d13f740c00f3003df30c04030100770033433d43c01c700010031444cf030001c4c001c0c00407c4000c4d03017000073300c0cc04c1c0300cc300c30500c011300c000f10c00c400040030c0f404417104000cc;
rom_uints[406] = 8192'hccc700c0303cc404fc00f04c00000300c0c0f0730340fc00c0c31004d43403fcf01d04c4f40000304d300033c7fc0d000cc000c430cc5410cc0030105000330030015c410dc400fc030051c044003f104004f03370111c33407d1f1040341d301cfc10ccc10004d700504c04303400f35c5c5d7c5c00c044000d0c040c4004003003000403c40010000400c0f01007f0041100c300c43340fc3cccc030043433410010f0301c0c33000fc003f0f334c4c004000300c0cc301cc0115c10500074d430f13c0330cc00005430f03c404c5100c07334f10c0040100003f504070400f503000f1350ff040403033000c13700007c4141c40f0140033000ccf43c0301374c0000501cc0c030cf000d1f04300000fc00cc130000303004303440c000f3044cf000c0f500fc5c3c1f00c5c44c50cc00100f553400000f07330c04fd531cdc44444010f300001cc3314cd4000003030000f3305ccd0c7cd7f5fd001c0ccc40f534045cc4404c0ccc0314fc0044030c00303c431f4d10d0fc710c7030f001f0f74dc0f11d100f70f0c1c040000100330cc00000c141401c7c10000540f00331350303c0c000c5f004501033075f330011300c330c1030c40000033700c7041005330010f100410035cd00310c0010040100c00015c471c4040000ccf30ff000f03f0351d00403c4c0334741c4c04070fc00f0001100000100033c030f0c53f00ff0005c51dc4c43003c3140cd0013f33007c0f1c00fddc000301d0004c00000001c33f41c00c0001f030430313011371c0d0000fc5f010104314034c03c300004c05134001cf100cc045054f33000400c0300341f5d00400553f40c0cc133f1103110c00d00fc0df00d1030f01010340c30103103cc301000140cf00341354c004cfcc03130d1330033353cf43c10315d1dc100000c0404ccccc1dc04c4c4c0cf01103401c0c4000d31cfc0c303f40cf044cd00c035300c5000f1c001005001400f4d00000101340cc4073cdc01300000c3d4dc00334cc103c4c30740030033004011f0330011000c3d40c1000d40cc1d35f00d070500453fcdc0cfd40450fc75ff0c35d00003c300400040f40d4cd0cc04c4140000000c0c104f7400335cf30c0041303ccc00c0f01100007c0110f40f04cc300510c0700c00f0003c340140ccc40c5d100d3000cccf000341c140f441c5073cccc0005d3c04f004f04d30c000573341310000f4170030040004c1f000f34f101f03530111001100f030300c100000c3005040304c00000400044c07c1f4fc31101f0000044f0f0cc400140400004041f00d301300fc5fc70000c1c01d4f345300000300001f000357c0f000f5f01330c0f04f40013033f100c0fc01005f400154c0d03f070033401140400003f440f007c03000c34d440114f03037c00000f0745143100c10f00003c0c3;
rom_uints[407] = 8192'h31c3010c04041010030000c0100c010ccc000c3014f0c0000410041051034d0700001f005405010300040000400003010030331100c0cd35000000300c00f00f0007c04c00100044d0000c103140010000000070c5c0c40030300d3000c4c00d33340004000003cc00f1f010c00100040000000047c501fd005304c0050c0400c507d700cc0300c740000030300340700c0c0000000040000340000c540101c303040030c03c03d110311c0c0400c4100f50004000010001301301300f0100d4400000c0c7041001c0cf01c030c7300c03330c1000c05040cc0c0400d40400c0c7c0003000310000c00c007f3100c1113c040c40037301040c030c030000000100070300034f100430444004000c00000140fc0d0d00d7c44031005d010400c30530c100710c0104000033143300c3f0430000310770000040101000f7c30cf4c0000404c03001003c0400f041000c40010c0400053400003004c711004ccfc0c034041500100d1300f000030104033000310004050104007c00040400304cc0000050fc0d000040c0300000040030c30700000000001c00400401310400000041d33c00007c001c000f0100040307000440004f0531004c1c0044004000c11000000100114103011030003444400140d03307000c0c11700c00f003030131c0000400c70000413134100000007d0100713050cc40000000f44030c0000030d70400f001cf010f000d500c5cc040001304010043cdcd04000c3c013041110f030700c00d5c00034c00000400c0303001c3c0410101030100001f04073430f00400010303000041400c01000c1077000003310c0040f403040004101100037010cf3d034000c70c4033000000300341007101403400000c1300030100043015d34ccc00300004400cddc03004c414c40304474331000d010500c1c300c44c14000ccd0100040c0c000c07000c0fc5cc4df4c010c40540c130340c3300cc0f00c7501400d00000030000000000313c0103011c3d00d00c0010004000d4010001171300104c47030100340f003c1d310534013073c000430c00c004c0000011cc0031000100431000011700c00040cc000c0037f0000d0f0d00003001c707003070101000000000410101d030454403c40001c3000d0ccc0cc070310c1c00000f4d01345f31030c07001cc0d00000000503130f311c000101000001dd00040100037300004307070000dc3405000100000c3000040cc047700c0c30000fc03000734304c300d000c3013340107cc000c00030000430c53cc30c0303300003000110df1c40031cc70340114c0003cc0000000050c00cc30030300000300000000d00000107c30cfc0c0300c000c434c0030000040cc040cc00cc00d1c0000101c0003401040011000103140100030dc03cc0000341010c4c04c4400030c430000000;
rom_uints[408] = 8192'h4340400300100030044010c00c0730c40100cd3d030c0300371ccf073000c40000034c10dff30c1c0c100000030303cc0d0003c00000c010c300c73cc104c003015374c03fc0370000030340c414400100c0000130140000130003cd0300c0000d13f0c0d001c003031040404033c0704700c0000d7003330dc1040343c100041f507cc101000f43c4f000c3400000010103040000c0c31043c0d70300434347704004300103c30031f001300c1000001073c000040dcc4000400001c01c0303000003000003c000034d0701004000303370c0333304c30004d0030f4340000000000c0140f3400004000cc030c000c00300004040001001c0030034000003cf0300010000004143013410700cc0c0c30d4504010053300ccd504f1c0c430530c1310000c7030144000350704003000004304001710100f1c4303f0f377004c50333c0c730400f003cd740d0340d00cc54f003030c4d0f0f3000d040050033000f03100307c471433370c10300d030010000040010504000cd430f100110700f3431c0c1c0c0c04f07c7c014040f40f0010c30c000000313c011100f3430c003cc043f0300003dd700c00331433f3c3c0cc04301104c100003000030000f0cc7400c0300041000400f011cc00300000c1c4401300f07004304000100d0c001010f000cf4c040cc410130400300400340403000000c0000f300400c0140404f73030c00dc004c074110333000000100f0000d000030044010cc001c0c430f0700000030c0d041c0f0000370f013003000330400000cc14f03000d0cd0c0004130300c00d00010030003c0110f40d0300c04c41c43010011cf34734343010050000dd305c400d041000cc000c0c3001c4dfd1403c30404033c0344c000001003400c3c0003040000303c0c3301030f30ccc3c4c313c3d000130cc410401cc340ccc0430c00043301c07f030d3f3000ccd0131c404303034750c00040000cd00c000000c0300000030f004304c34c0c00c3030fc3cf037cc01040c104031335110300070000004004010003001703404003033010001340d00fc043400d10000004730053300700cc1c30003300053303cd15d0ccc4c10c1300334400331c4100003ff0045c30100700137004004000c000075040f10dc0333d3401030400cc0cf0150430000c10000cc03d40c0d3000f00044040310000c0044040004d33700000104001000030010300f44401d00cc1003444c40d00300053143d001100c01000400413033301100d00c0700cc03070cc0373d070c41ccc005044c00000f00003c00330000000000003c0010307000f000004f3fd40000043000400030c00440c017405c305cf0004f00c00101c31000000401040003003330d000070443300044000000710d3041001031fc00c014000c4c031f00003034df0d01c400000050;
rom_uints[409] = 8192'h1000000000fc4010044001400000c00033c33340dcc00030041dc030431330004110000370730000dcc013011070174c03003003350031033030000343340073001153400140000000004f00010111cd303c3fcc111cd40030cc100014011c01d3000f00301374704c31f00033c303c4f3c00004d0010fc00c3f177000005014f07d73400330c170c00c0070003000d033d000000043140033031c0073000100040000f040010f000101003003503c40c03f70000030031c0c00000c50d00004103050c000404100130040500000c0301d1c301c0c0703004000010030d0000140000300dc4d017000c003511c400010131000400dcc1c040000c0331000000c0040033c101001000010430430c0000444314dd140100c403040400053d0c0000170000c03000cc04150001340411044c70000301311f00031c013054df000013000400c503c04007400015004001004000cc01345003031c40c4cf011ddd1000d040701047714407d3dccdf3440400007c03000343c3441df4c3007437c103510cf000cf4000101cc40c0c77440c13c300040c470033c0d00f10070031330d41c5fdd00733041c00513003c70104010000d444341c0f000335430001043f0f33010410530cc010d3071000400c100040c40c4003140300000c04f31733303f0301ffc130c50000cf3c0300d0303000000c05c043334357d000000130000fcfc3010337d313c0030f73000030c4c05300ddf03cf31d0c130033cc33130314f0017050304001cc011400d3110404c4c000000700c007044c0004f00c00000443004003c030003300003057040d300100300c10c00100110410d70300c03411403c074c0c041dc4cdc01d0340130010c714040c430c0507340c111103071c1cd3301c403c00c030c74037d3d7d0010500300c113075c3c40c10d304c00c407101c00000370c000000cf53034103d0c3030403dd0cc0350014000070c00401000701010014c0000331d70400030c14c7c0030c0c710300c403ff01330404c13c401000510cf04c0040000710747030030d00c3013703c0c00000c0c010470c10004c030330001d000030030c0f0030c40107c3030301001c00041f0403c4f44cc0000500c1310304004c0000303c0401000c11cd110c4c10c3003400c13030043c01fc1c00cd11dc3700000010114c130334f1d010701103c4103f3501700303d1f0033374010c03030c0c0c0050c070000010704d0540510d1d700300001305fd5004303c00001d40730430000303740001c0031c0000140004010010433300415c150010c3c004030340011100431003000001030000c0103000070010003f330030f30d000003c4f0003f03c01d10100400031004010d0d010500310fcfc31c000c100040101300005c0c30d003f43071000f000704710cfdc401f00d00300c;
rom_uints[410] = 8192'h4cc00000ccc3c1010dc000000340d1d0d543c03070043c0300000d0c4034c00c000dcc10d0d30007400c10d14543013077c301c04000147c301000314dccfc00004cd3dc010c407dc000dc101000410c50101401040100f0cc4f11315f3400d30cc0c10433001c00c0d3dc4003f5f4c000cc0cd444504d0500cd7f00c0404c41c0434ccc0c070c50c01300c10040f00c007400100030304c0500370004d4ff0000001c74003c0d40c00c3040003f00f000003c0000104c40cf10d0013c030000d4d30430000000d3410400310f3300040c10dc74000400c000dcd03410c30030005000c343004c4000d00370d00704304450f4300f00000c30044500f11010300040750c1041573c0000cc107c7c0001f0cf0300c000cc1011d005d5314f0c301c31070003040740043103ccf00334f034000040000000c0cf00ffcc053c04454c41000004100500f0c3004435c000c0d130030030cc0003c1701f10000c043ff040344415df0400c0001c40c03cd4f04c051c4011c00f004450100040f00f00c4054c04d3030cc3050401000040dc700000300440c045c0404c400c050413304cc0dc0033010470041440c00c4c3c300300cc7110c000007105cc003401dc04107500c01140104110545130dc101040411013f3001401f70041035414cf034330050c7c4003d0c00371303001dc01d4347031c00cd00430103010004f0010410300131c40cc00001000cd10c3131c5000000c001c0010000cdcc4cc1044170430103c1031dc540f0004cc404545005c400c1c1414c7030400df5570d100c41cc000d03c43cc4c013000403c3003305cf0413400f50341c03411c00111fc4d10c013450c1130104c00010003c3000013071c31f0044cccc03035301000d000001001c14000100104d0105cc00c0405cf0100cf7341130cd0044cc00c0d00471d44110001001fc00310304d3c001cc4cc0cc700403fc3f00c30c103410034f01000414f00c0001304401c001f04cc104cd0c4030c00f300435000f34c41305f5d1c00c00070cc00c4004c103435d000c004dc00040c07d000001300101c04100534354f01c04000440cc000ccf003007cc4004010030d1340000c000044c300305ff00040701c01100071d0050735004007501f0400144100c3cf0cc0073c001c30317510c0443c10c0301400107c1000f000c11f4003003cdc430c00dc1534f33100cc333c0040034303100c50400ccc00cf4f4044100d14700d0c0c0c4c45303400fff3c10005040c0cc40ccc05040cc33000dc00f0440451410c04010700cc401010000000001cd0f000710f0c00f1004d00010d0000001031000041c4d30574410014043cc003c041c71000f31c100c40c3f304457107cc00c470101014500c1040043144101f0c4f0d0405311c01f330cc0010103041c045c3174300304c;
rom_uints[411] = 8192'h30410040034000c4d04c03034f007cc15cc070c4f01c3f0000c0001000d3c0330041300000c0dccc403400000000351370f430c0005c0005c01040000cc0f00013c0c000c040003043003043c0403301000f005173f000fc000030c0c00f100cc0134000c1340ffc0c003c04101470c40cd140fc4c1000c0100310300c340000d4300cc03fd000100000001cd00054000004103300300040c0340040c010d0500000f04400f0117f10c74000c1c3cc5000d50c4000400cc30433001dc0f00073700c0c3f400040400010100cf0c04340000cfc7001c004dd01c10c410cf41030c00000c000c4000c001000c300fc003000041030f41d00000000400440000030cc000004310303104000004cfd000500c150c3f7c0d03000313c40441f3d0010f0403c00d0510c0001c0f05c101000cc00c030cc04c04000c3030010300100c0cdc10c000c13cc000034040c040000c01cc1031334300c135c333033001110c03c34c050317010c0000003144c00c14000000000c00c1040103c743010f01d004450440001110011dc0c4040cc00cff4c000014030c01000303040c04001d000c0c10c0c3c01007340c000030040ccc3000c00c0141c4110c0c0f000cc00dc5c370f50c0304143103011000c4100100050c000400000c34000cc03040cc0d40c30c37cf0040001c3c03010c0c010001c40d0c00c040000c04044cc00f000c00f300cc0300033001000c10001504cc000103fdc0014000c0010c3cc710040c0c0c00050c030f000fcc000cc0000d10c700c3cd11c40401c031cc4703710004cc010c0dd3400c0407d00031c0c73c001443000343070d0703400d0440c0000001435f01004d104100d30340d113010000000f05000f005c04030473015003c0c03c14cc34040030010005400c00f77c000fcc1f013003400c4400c10c0f00043d000c30c44030110500c443c00400cc0c0001f7333000fccf3100c0000300543005440cc004000c0003040c04c4070c0fc104c0cc30400c0f07000c0cc403040c03300331500301000c07000d3001000cc00cc00dc500100104313000030353c007040c1007140000130004000c004404ccdc0d0007000c3400330005f00007c1cc000c0c13c4c0030c00740c0c0001000004c0c0c005c00000c01100c300000300400704c017cf0c070004f0070000000040c100440c0304041504040005d0070c0040cc0304040c000407cd100c040000c0f334000dd400070fc0030c00000115000c00340000030003040c300400c3031dc30003c00c100344400c0ccc400c0040c053031f730c000cc4000000000c00044c40000c0c0100000c1000f4000510340c0f04101cc3cc300c40007cc000c000103c0001d4401c0c0f07c10301cc0c4c0c000134313c003c330c11031d40c00c400c0c0c0404c143ccc7c30c000c0;
rom_uints[412] = 8192'hcc00000d0d10c343d0407150d300c000dc100c4030f3400001c3c0f1c34cc000053c3503030303113140030f033070c3170cc0c0d30030700041010101043000f0430500400030d000000100405000710c301f110c0103c00405cd700c00005001d1d3130000c50d31347004001033d0040100007345000007c0033043c1000ff4000c010000000d1dc003103000001310000000000344c0030001130d4100300340c013d10001c400cd0d0103000d300c03000004f3101c0c0000404110000f004000011305f1f330c001030303c470054040000000f00c003c0033f3530003c000c0000340000040f30470050c030404c33d007040000003c50301030000c03030c030411001430d5cc001773f400310330d0300510400011300304c100c0700400000710107043110044450000030c37303d40c000001000143c3004547cc300cf0d11040c0311000403d0cd10303c1c000010573d4c37c01c0c00410c0700300013c70c0100430010000f0330040c4044010304104cd0051c0c00f004c0c41c001c03304101504c000c330340070c00330c0000c040c4740000000c000104c31cc00300301c1c5c3fc030010330000c0c3404cc3400040404c000c00c0c31003000000c4403305c00f03c0050041c0304c70c100c00000d000d040c1030000000401030310c001cc43c03d040007730000000300000133003f3040030000c104073031c0033037c0c011c1c344704f701013c1c0c000003c1010d00304d0435044d1c040d130013d0c7d137000030c7000000c0c41000040030000030fc15344d03003cd40001000000c04c30003031d1001005031000c013c03c0035ff43100c007c000c3130100d44f0001034c3000003004033d301103c000d40d01cc3d0c00151c000f34c4100c3d3c030005047073700505c1410000c34710c0000114000000c00000107004c0705131c474c030dff030013ddd3010104000c011040df001000003c053740031000cc0c34000004334cdc00331431003010d00c4300001c010334030c30041000140d040f110317d3000f0004c00103003043130011103000101500403300037100c00004304c00037003c01400030cc01c331130040000003430300100c41111300100300c30400073003010110c0010110100043f00100017000033003c040110043c00040000c300300c011f00000c01004cc011310004030000400cc33041030000010000031004370c1c3c030000000000014030330311005f30f1013075000d704c01cf0c04dc1c3330c700df0043cc00003003304c01043fcd0000105d030010c1000d4000700000030000030030110f1000c0334314040d001c030401700000c0300000000003110001c1041cf0d51070f43034c110c400000f30003300031c0fd0100400747011301440d31f30730100;
rom_uints[413] = 8192'hc0c5c0004c0441000c040343030c03003000040fc1003043c0704c00c001300400001ddc400000001040c0ccc400d03c310c05010c4404004fc40f33100cd400c30300c00044334040000503000cc0010cf04400f3003140cd70c0c3cd3000c004034c0000c0c0044dc37cc0000c0305c07c0c041030074c40d1fc41041ccc03cf5c3f00000c40144007000100030c000f134c0000c03c3fc4c34c30100c5c0c40304000014110c00c00440300c10c10003d4101000cdd014c014c000d03c0c0033c104000030c0433c4410c0d04c7c0003f5c47c0ccc34c34cc4000c0f0c310cccf000f3340000004c0040fc505304000001c000400000c000307000fc10043340013d00400444d00c40c0c440c300c304040f01043f043c130c5c0c0050f00c031c3000c04c0c4005f4734000034cc500f00c0c000000040cc303c45d00cc144c101030c0c03c101c03c00000000400cc304d0cdc00c037c0444304030345003c40cf4c0c0010df300430430c500c0cc0340011c30050047cf0cc40d0c0f00517f0013d0407043f4c704040c00c01300005133d000001f000c07c4011c1c0c1501cf004cc00044c013031000cd0403c50c050d333c00004d340044004077001334040cc3f00034c00fc300000300001fcf400dd030c001000f00034000000fc00310000dcd0d40cd004c0313003fcc11004043000300044c5d400c0c35c044c044c0dc10f3400c0f5fc71c3dc04c00c0040001cfc04050030c700700c34c0041407100f1cc04110000000503000300c0c0c130007c00050dc40503c040f0cc400000400c000c0041040d40c40c00004c3043c0c400d14043f705f0cd4100cdcf4c0043141d0c3d1c3c0f0c0f0c00c001dc00d444f3c10000044300f0034c000c75733000000000004fd5c0c537001ccc0000c0000c4c000400cc03c7c000013073004d0400ccc0003400c000cc4003cd0c03340c00010300010d700310c00d004c0c0014000300c0c0034c00004003c0007c130c041c0cc5010c0c30050d0c1000c7400703000000400000340c430ff3cd415f0f001c00030cccc34040340001010cc1074401430440000140cc333f0cdc400303004c01443540043c00334d014000113c0040c00004f403c0044100000c0d41000f0043710d00c440040c0c00cc470f50c703cc010c040131000f100041034d3000143d00f7300c00003040050cc01c0541004140f000044301400c0d000cc50cd0031cc400000c40c04f01f4000c01cdc0c4000d00c0c013f4c41c31cd0cc0c05cc0005503c003c51000004404305c70c4c140003003004c30007300404cc300010d00000c0000c40ccc0344c00cc433ddc0d304443cc0c0000000030c4000000cc0c00c0c07400000c0c00c4c00003d3340530030430c70440cc04c403fc507000034410c004f0100cc00;
rom_uints[414] = 8192'hdc000007c40003cc101000004c03004004f0040c30c00c14303c000050c4104000401d0417f00000334c500c0030c3001f1c0f0fc1504c0050c0400000000000400d10040040003440010014c0040000d0f00710400c3c3001c0d330030d00000010f3c37c4c1d000010000440000c0c0c000c3c0000341010033d1000d004003000c00c7cd00c100c7000040000433000004c400000040400043c04001000d44000cc403cc113300cc0300000070100001000000010c0105c40000c5030031441c0c07404400f1c00101014404c43330144300401307474100000300cc4000c000000c03c400003044003dc0c000000c0c00031c130040c00000c1010c000c00000000030c0001ccc003010c0004000000c0001044c03133011045303f40d0c30c000000440030c000f30000c1c30000010003d04300000100c04c00dc00c0773f0003034c3170100031c000100cc14143c0100113c1003703000fc0c100d00070004700d0010103c153cc04000000004c0040c50070030347470300030000c00144c1c01000100104400000c00c00010040c4000000000344f300c00141003dc40307dd03c0034000400101cf7c000c44057cc1c0df43c000c5c0440001c101c10d01010701410030c0330c4041004447c503111c430c0100c4c00400c10303000f7003c0c0003005300000314c01c0000c0140c0007301cc00010c0101f00704c011c54003000040100d000103300c003300c10031100401404044410000300100000000cc0000cf73c0314000300fc30c0100c0000000010770000001f010fc040003c004000043c30300000340003504000043030000003070c0010040054500001110010440314300030c000000010000007004000104510040c004440033400001030c4100000140040400037f030000440c4c41014440c00000f001010000c10703010340c3300c0c4000000300433410c3004004000c0d4304cc4000170f0cc0000000303000cd0574010701c0c0c0004300330c1000c000c30c000c000303303000c0c0037000c000034000041000c010010c3305d1c300030c00cc004000c004007c0040040000cc0000014051030c01054000cc00c0400003000071004030370000d4000d403300c0030100400013000101100f040304540dcc04c000403030130000040003c73401c00055ccc104cc000c100c15400170030400000001c003004dc3c304000140dcc0cf00c310011404c413d040c000c100000c01c3c030001440c0c501c1003000004070077500070c00c00303443fcc00000f007c0500c0030500000400cf003c5000000130cc0044c04045c00001c00000c0041007c10000f30000404c04ccc000003c000c000000c4c10140140000014030010031d3000100000c403000cc0141100033303000030001300407c3003040;
rom_uints[415] = 8192'hd50c01000010d0030301030103104c00310f1134d0030c00c15004001113d04000001004f0000034c04100103c03d03c3370d10744033d373f000000dd30d1010c05043c301004c7d1000414d0003c00043d3fdf3c0d0c003c0c10f1c50331310030ccc0703070c1004d35740100335c3000c514cc10f03d100007c03d0130003537004434c3000c040c0003100010000101013500c1000cd01034003c0d40003d13f00004040cc400100004c000000400430c1d000001cc740000c0c00170013c50303c7000cc14073f0400033c3dd11034774c014cc3fd01f007001015010030000000003cc031004000dc001c3c0400173010030d00310003300033140001c013d1001cf077c0031014001407733c300f30101054d000453010cccd44fcc000d0f300400100d003303f4044003f1033501c3c333533c00030d0c010330d0c3410d3001031c1000c334fc10314f1005cff0c3c1cf5030f0c0030d7033300f300c10307dc340fc0c1033454f114733300d30d550c10500011700550c0004400df301f075000d34c0c533510f0000d0130000100c030143015413101101000c1d5cc00000333003433010f1c14f700045c3c03c354cf0100070c000c0d033c400303fc401140003dff333c303f0c30c1043140c04c3000f0000003004003d070131310c717007f1c4c00d330f0070c31300c330454300031011000cf14100c1c03313c540001140f410c1f3c7c0f350c0101f0100740c0300303313df3ccc04cc00dfd44c03145300310f130cd0013314003140040c4c10d0c543c311d00d7400c0c0c00400c300c0c030c3110c300151d0c11c31074f1310000040c000c041003310401fc3100c407c3c3c000330c00ff340f00c07314000f1003000000c501000c0c44000003300c05053c4314010dfdcc30037c31173d000d4300fc3c000fcc00301c73143c070c10304f0c400011040fd43c04030d00300140c5c1d00111cf0754040300d300fc0c0075003000441c10c040001cc3030d1f033333d000303000f003d3304c0000040dfc3c3f03041f4cf0303c0c030c11400300350001cc17dd0410307000301000c03c000300303053cc303c30000c00fd000c1000443d7fc10c0030330d0103001000001c34c41033dc7f00300405303c0fdc00407410f310000100c017030033770534d04c03f13c01330315c0017cc01f001c3f3cd4114015f0c000000c00410003433000003f04c057000d34143f0f04000133c300fc303c13d10cf33037001c0001fc3cf40510c40f317003331007dc33cc00000030c0400d00003007d00c00f1330d003300cd000cc1c043ff000173004c140f33077f117307773d3031004c44f0cf34000104300d00cf07f100510043004c0c5405d0303111400ccc0351000300c03300173000c0d040f01fc00014d400000330;
rom_uints[416] = 8192'h1d400c01034100c1434000000300000c77030000030c5c0c00070f00440045400000c031ccc000cfc13003fcc0cc4f0d1ff300c0031433f3c3000c433003730c3000303300c30004010000005303c430c003401033034133003330400d0d00c0333f00010f00034c3100070d4c4c0f01074030c0003100000c00cf403700050333cf4000000000000c4343440100c104cf0301c1000c0dfc400d00700045074cf00c11400d07d14c01070100440cc333c300170100c1d040c043c031d103c7000c00c04307004f05c0070440c354f30c0d1f00440c4000c10c5103dd0c0c0c0c100004c001070433c50d43c30440c3300c41c3430cd000c3000440c0000d00030f41011117330f0055410000430c1c070330c040c0001d04c107400f41d3304143000300c0ccc0410300c3300101404c000c000703c04300344401cc0f0c03001300003040c00c00040c01d30001030c30037c40f4330c133000470c03d0001400003c00cd3000004407c731030014401041301044417dc310c13410010011c03440030000040401304cc0007300331333000003c3001cc000c3014005001003500301043ccc4c0330ff0300010043cc11175404d41fc031004407050073c103c1413000100f03d0c04c03c3000030017007411303c344c301cc1c34101d07c0c000030101d0d1730340400f0df134314703c3451703033304cf4c000f43c04c000340c4d0030400c0fc43f1000f04c30d07c03000430c034f00f35704714c500d0400c3733c000c007c4cc035101c00c4d10d0000003144c070d303c0001d4000040304c000010010340033010c400f001003314c330007004d01c01c0cd531c0d3f001070400c11340fc00030144001fc340040001100103500010010c3334040443000704400c40cc010f0101750340c00c113003403000130c00130001310101430400c5000c0c4cccc300030f3403103c0fc1c37040f030cf0d3cc004440144cc0001000040300c04c003500013000407c4031000d050140c010f00070410004001000000331cd30740400c110f704010c4c0c3000030030c34004400004040c00d001510c433100cc00ccd0000c01314c04000c44030440013000003f0c47010c00000401400710300004003c00003cd0f00330103d043030d0f400c01c00d0100c3301050000003000c000400010030f4cc010445f7400000c00dc30040004000007700130f000010c4030001070cc30c030c73f0c37cd04331430010070f3f30400044c303010704c3430037c001001c0003c33305310d100703100c030510033440c3004440c300c443030c00370405f500d7000000c7001100c0c3010010c7f0c3fc3f40004d0030cf0004cc00c00c04000c4c0300400300170cc04701000033c0014000f001003f04010070070040400037c3013034c003040001;
rom_uints[417] = 8192'h1100034f00d0d40cc700d33414c30315c0010d003cc33000504001d4c0700005d340d1d0040130700003c0004c700c707c47cc34c5413400004040003d40030000401004d30003c00c031c300c0000f0100305dc013031417710c47f0143030700400f40c00004c1003410004f333c0ffc3040c3010ff003c00030430000fc344730300cf004c0c0c00030300c1034030400000c03040c33000fc330cc4c3500344f3001c700300f04d031dc04c4000c15003003f53f7005130f7f31c105d00300c04400041c34d4000c4dc1044004445743011f0000000f4000041c401c3040f00c003030010413104c4000cf37c0c003c000c170000000c000cc0040000cc04010cd70f3c04c4c400f3070c3c0c14c015d07003000030d0340c7dc3074010c44c00c30c4c043f0d00411000100c0c300f0700033dc0c30c3004c4d530c0110c0c3cd0004cc0c0030c400c4c00c3c0130000c1c330033c4053c40c7c03c0c31c0040c00410c4c0404c044403007100c3c4c010f00c00c04d00f0010030140c00403cc30c4000100007004f011354c70004f3c0c0f700341451cd30303f00c4710010c000004c0cf17f3047c430fc37c3c4f00cc0f00331c0c04014030f300100000001cfc343003c0010c0000c043014c00c00ccd0dd0404000c00d74c404d7c0c3003fc43f313cc0000100300c00007d0f0cf00c01104c30700100700c100440037700c5c030034c30f440c4000131405044c103c100d00c4000045011004405000000101d0c030d504c1000c0c0000c0000040000f03417c00c500fc0034f0001c0d100c00003000004dc340f00400c0c3c010000c0311710030c3400dd0330003c303003f0301cf301040000c0c404d3f040cf300473cc4c0003d0f4c1040f00c0c500031313304d0070005c001c0114301d300cc000000c0cf110010d4f0005c4110300040047037434013c140405c0000d0c00000301dc5040001047c0307cc71000104104c000300013cc03000070004f30c4404101004000c33003f001d334df00c0c004313417cc0004703103dcf0c0c00007d00370004d00fc0c3000404dd4c000fc00000073ccc00440347004d0d4c00001413c43730cf0c07d700004001010000f43410c0c03000400c044fc00c00001300cc41dd40041400cc334d04170043000c404c04003f4300450000040304c000d3040c0f300c1c0cc30cc3c3d0040040040031407c4cf30c030cc3300000000153100f44040403003030c403f4001cc0140030c70301fc0004dc07c0040400004571ff40f3cf0c00730000004011410300c0000003c0c3340c050341cd00d34000000300041c300c7d0cc7ffcc0335550000c7301c0700c0000c40c001cf004007c4c003ccd3010303f30010c34c000f4004000c40040c03000000d1cdc0d3c4040c400cd0000000;
rom_uints[418] = 8192'h14c00000c30130d004c0030030c330df1400131c3c0041410d4040d0410cc00037410d31c0000cc0c030301044c0151705053000301030f03d5300fd003c3030cc000c70003040010030c050003ff00c3c33010f5f30030517013000033030d51400374c30000c7300030030103000c0000030c04d400000000d34df073c40004c1d004f30003c000c00300001000300c0400c00001015300014003003301c3c0c403010f107103c00405c03300c700c31300300cc00000d01000c41c00000700030d0101000c0fcc00c034700fc3c04411c3c4c001000710d30703101c00044c000000c340f1c0c00103f010c5c00300100f000100000c00c00300c0000c73010403cd403f013c40dc1010d3c0c3011030000013f14007c1c01505f431f1000c00c003c400310303033d031000031f0c000000c0003000040f0003c3000303f4030cc010f3100cd140403410003440c7403c03310c000f35055cc3c0cdc03004443103c0fd00000c030c050057ccc101d100f00fc0030303f003010000f04c30c0330f43130f0000c00c37000f000440040000304f130fc30c070c0300004007cc000fc70000c0003003301101d4100c4003cf0cd0c000300040403017c00f4100c0330003033000cc4c0f7c0dc4c5c0440000470300400103001034d031000310011053030413cf10014003f0dcccc003c03000404cf30000c010030301031005401343f30c10003c0001100c003400000303c00ff34300013c4f0c37c0110c3173c003c01440c0d0000014001101c0ff400c0030c0c34fccc001c3030c00c3c33030c003f0000df40000043c00104003c003fccc00001cc30003510c034330030cc33050000014000105f5d30304004c10003003070d03cc0000c041004044100003f001c30d005414333000c04c3f1c70d1c74d41f001c55000710140fcd330c30fc3330000104001c000c0c0f11101404d00f0c030034033070c0003400101030000000347400404cc030007c110004001030000c10f0401000c3000004000cc0330300c010000403fc04000004303f73033c00c0300000c010004c03000030003c00003c00000cd0303000143f000c3c033c00001007301331100c1000cd00c10c3317c4001c30f0300103104010000733c0134d00473003ccc0433c00003c00c400000000403c0010000c004400f00cc014000004c0d5003c173443003000331f0000005530c0300f0c11030c301c3ccd301000c000003110700cc014c0c00450c000000c0000000c04300040705100ccd00ccc41010130cc3740403c30c405c0003f3c0000103000000000000704701430310000003c003c00307c0c3f11300cc17c1c0c0c1c1fc300000000001014c03c004404100c4df03d00000d0c000000000c035d00043d004030400c000000000700000105010044001040;
rom_uints[419] = 8192'hf0d30c0cc0d010470331044c4004d0741c03c000c303f040c0d00cc00400003cc0100c17cf03c301cf04c0340103013fc4003c337100010c4010c03c43373dc00c40f050f0dc00c314004c4c3100403fc04044c3c3014001f0f01341fd00000000c010c3cf000000c3017c104d3003774171c03f0110c004003137cc013044d0c1ccc170033300f100c300350000104000000c00000d331c00330001704c3d015cf30000c331400340003431303fc3dd100100000011347071cf0300300370101fc10000c410130c345000007c3c470100513f31c334007f01400040d44000c0400713310705c000c41c043103fd00c400c05005303c000130c03001c01c00c0cc0000403c300041cc400c3005f30400003c010041001cc0714005d0c0cf47c03c40070007c010f14300300040400000000000c0157dcc130c1044c1cc300031ccd0ccc003d504c01ff0040c0013003001c000c0c00c44001c700c0f105410040c0f00c13dc001414c0cc41334cc414fc0351df00131f00043173fd00100340cd3c013503c04c0030133c4f07c013d00c100f1330030c440f03c030cf3403001331f700cd1c33cdcd010f700c07c3030cc0fc10410400c01c70431000c37f0c14d04055c30c30001033403000c00d071df3c03440570040f05d047130c3c00c70004c3133f4c73c030470c000001000d001030430000303f3dfdf000d1004c0f1c0001c30c000000003010304d3003404530014010130c400071011044140c10070031c0d4c1000f0003345014030033143530001cc041300310047c4030d1cc4c00c0301401c04c0007117d103304001107700300c10c4130dc74c041350010307100000d00003f0113f3ff33c0000300cd1470c014400454f100051c0f03d10f100133c0c0c0037101313f0c0c073cf03f3c040f31300000f4030030d003d330f50c07c0fc3d0313c0cc0034c04000cc00534f01f30d534c0c40c400cfc00c040030151000c400d0cf00c0003100070000141f100d410cc0130400cfc31434cd00d313c30350100030c00cc0c00000004d44c0000d000000c4c0530134011000000c041c40053347010c00033401003000c1134054010100000c0c3c50031f314400410000c00000040003030c0350c140370143f70441f0334033000001430000d0c13c0c004000c3d0c30f01c1c0034f0313cc0303004d130400c0dc440300340c000c3cc0754c014003c000d340ccc1c31410c0d05c037d3000d400140054513c44dc00000c31c1c40cc10435f37c0fc333c040d00000104340000000f3501c1341143c003d00030300c00d0003004701c410003344c301010034007cc000c0355703310dc30300fcc7d703001ffc01004000c0033c311000d440334d7001310c010317c1dcc3f00c034fc7310110000033c0000f1107003c0300000000;
rom_uints[420] = 8192'hc0044000043010c3c000c704f4004104103000cc130544030010000300c110040c4c1f0030c0000c01c0404004c00137400c000001040344c330050fc400044c0c0c30000c070400500c1d4c003110373f33040050103034340c5d300010040004c010f1c030d415004003114ccc000011040c0031000dc003c00030330130001130c0c040c00033c1400000c00000cc07000000000034f4cc30f304c3c10104030454300000d04000040300300400104134300004035f3111004040304007440130f044000f13130045101101011f004414040104c00104004c00000dc0c301c0c30c00051004030000040c0c3f44c0cc00034c000c00001000014100c003c010c700030000000300c0cd000f0d03010541000110c0001330400140c730c4c0ddf300044d0000c003000100317040033400413c0100cc00d010043030000001434c0005070000000530300044005050300040001107c451410c00000d414f000070110f43100d10010f030103c110040c0414770c0004c017315000000147c3100101130cdc000000040001c401041000050003c0100103053000cf33000000c5115c00ff00001310d0000f0d03f10433010ff00cc3031c400130cd00c153c037000cd00400055300c000c300001533110004000f13034701cd0c0c0c0050330cc400d0300c30100df1c033011c004cc0c0c314c10000c150c1c00310004300014407c4004111000000030500300005c53503c1141d0340c1171f00c001440041f13143dc0c01c001c0c00300003033c7033100404c1cc4fc0001000c04000c0007431d0c01701003c0c1340014c00004041c0f014c001f03c1017c453f00004010000310c0d000001c01010d0000cc045313cf0015041100000101c004170040f1310000030331001450f50d510003ff01710c5143c0500370c00000003c00d1510c003c0c15353301c40c30014cc5000301401f01001d000507c10010403c0310fc40000c000100310311000c1140300000d3ff00d3053000cd3ccc04cc30300000430031100004400344310c0010440001340f43c3c3c103300003004005d0f0004304443ccc300007c100c4030070c0c0c3000010004441014003c5704530c00f0c004307000c333003003dc000100f03c337f4000043000c1015035c3c150017010cc1041014c137014134c005c730030003d300c040c0000004444c00c04000f00c4004000001000cc005000000c01033c1401f4fc3c0400f0703c00340010005500c004400100cc0040000000530c14104000c0000400c00000000440c00300f5001011000000050c50305c0005000c34000010330000001105111030301f00004c03530003cd3341003100134c5d00001001c0000411110301300050040030401301311c3c470304c01d51c0011500d004d0c4c07c100500000c00;
rom_uints[421] = 8192'h1c3100000f0f03040410cc0007070f31c0000c00100c0030301301314c4c51000333030030030143000001004d0031130f3fc0f0400f307000103c110104c001101cc1341c3f001c000003300543f000330c10003c010000c044c30c00ff031c50053433003c10c0cf0f3000c1d7c3c101003733703f1033000403f311070333511f3f000c5300fc0c00000cd0331011cf3100fc00001133cc04c0c0c001033370c1c1c0c007f03c001000cc1d150033015f4f1c0010041101300f1d5f0cc00005300f3030c0f0300c0104030000c1101f5033f0003c030040300000cc50000107000041c5013d0c0300045c133d1dc003037013c00400101000043444010000333c3f34300030cc44110c33dc370034005d5101f310033c1055c370531cf10103410f0007c0cc01031c35f34ff0cccc003c0013301100010000d000ff0f440030003343305400100010cd04030100151104c0001fc400300000f00c13100c000030cfc3f300000d013c300c004c343030c0011c3115cc04c44d33cc43401f404313337cff0300001000030df0c01403450000d000001311c333cf013301045445ffc003f3030cf30030330011fccf501c010cc37f01000343033010513010310d0d0174070000c0c1034330f000300c1003000000770f3f00d3133c401ccd4101003d351003300440c301307035030d740c1010401430003c5000335cc0011dff00044ff0c00f0f0101d1410fdc3cd404333310f00141f0f003141400403f01013f0c100403f30fc030d001130030c050c30c000c0f04330ff07f0053000fc3f001d43c30301100c0304c3000c13003010005c431ccc0041000301cc0d4130303c00f3040f003030040003341ff003040030000cc070000040cfc300c03033c43010100000c040c301f000c13cc1c03300c304010730101004c330013c0f3cf1115031033003fc500333ff70c04c17030c300f01c003055c111035c004033c0340050cc4000330f3300001c103030000133c000070005330c005053371040133700000040fc003300cc017030150315010c333f00300700001c4100fc0f1d3100010010330f7c07dc00300101000043001004c0f0000530000c07030300001411f1304000c3314005cd0003003c00113000500037140d00c0050033f10f30c141ccf0043373f00cc0f000103303030c003333f1c011001107f0c700c05cf3435c04017400fc0015f31000c4f010c00c301c330043cc4030301c10f000cf030f04c03f01f100340c3300c00130330300f01f33100c013000330c1103f00d00c1c30100f1130ccc40cc000f153c41100000d004300500030000301000d00c034f0c0310030c3303cf3000500cf31100004f00c3d53003030c310301c731033c1030c10f101001000ff01103031301330000fc1045000031d0100f103f03007011;
rom_uints[422] = 8192'h300407000400343310f0411c040430c40cf000070000007d30145f17343000f0310ffcd00c0101400310fd030f140d00305000000d031070303c100000141003f0001c03001c000cf005400dc004f1c000f711307f1dc030001c0000c10c3c710003f00d330c0740f03003400134300000c10100003c00c30030404033070c0300000c000f4004004c100000c1f00070003000304cf30f10300c054040c01010f5713c33d410013304c00c304c33005f1130030c035173d0140df1300100ffc310040c0d70f1c300010d000140100f0f371c03000dc00ccc001f1c100f3c0c0c004cf00030000c300d115004044030f314140030c040014440017c3100313cc3f001f0ffc0000c000dc74c714c1c141cf1310104000333000f1350f040300044400c04331f00c71300035050c0d440000c405d00003004001030f05d0c0c0540000003471000307001c4040433740431503d1cf44f34ff11cfc1030000f43d000310340c10170133c4f030ffd000345104413407f30300dcf130500130005774d440f310030300c7033f100543c0000350400c03000c3f34140031c0000c5114c0000cc00400007cc0003c0c035030c03f40050030344014100153177430044451150743333000004301c000f3403dc00310131401040c3300040040c3401c17013c11fc31001130f3034003001c0c001000440430300c303430040c373cc000133c04fc3f1000010313d0c0110c53000c04713fc03c0c05c0c00050c010000130070030001003f140000000340c00f00030c170030000305d0100000d30005010c040f43000340010071401403140700030fc4d000c15041333504d300100cc0000310001001470f0034c340f0451015014114010cc3701f00d30040510f4140c04000400c4014c0d03300311350dc11310710400740f30c005441c1cf5143341040d313040011c33701030031cfc0701c1070444305031003c00300c07540f30030003031010c01070410f0430000530d140cc0cf43003533044100050000770410c00334005000c040047fc540c011f17030000030330004301070004300d303031100c310001fd03100000ff1011cc1444003430140c00cdfc040d3c0c500c0000031c004430301413040000003c370007300441003000c41f035003130740011004df1350d70001705130001cd001713ff0c0003100503070000c0f30343c5c040004000400000000070300041007c0003c310c131000403c0001c710ccc4105001304100000ff04010003103cf01045cccf0431f1403100350107400000434f1f31d343100310030003310000c0c1340001050000340000500c007000040010c501333033f1005030041000100015f003407300c04000003003c50403000044f00f1f03c3cc11037c1004100100400301747c0700c000370ccc00;
rom_uints[423] = 8192'h31c3004000330c40cdf014c13404df03f3c0000340c4c133c03030d0f100503cc077ccf107300000073013c10c00303cf343001137300c37031503301d000c0cc0043004100000f10300f7d30c00414f405c10c7f0cd43300030f01c00107004040d030301c43c3003ccc305005cfc00f0403c0f0701f00100fc34c0f0c011c4fc30cc400cc000f0003f00000001140d30701300000033300c00f50c005f03cc30333074045400003c1000041d3100005f05010700cc1000031c00433f004004431000300404303cf00cf04ccf0000003410d0135c10cd50f013cc13cd5c0cf01c3000c3400cd030c00430001c074cfc0c33f0441f5c40300cf4010370000400c00c0143430f0043050301cc51c17000153fff0c5013030c404f01ff0414301c0000c000c733000144011f010417fc133c13c145000030c01fcd7104341d0403c00100cd43d110000c013700413c00303103370030c303037700df1c05747f10001407010fcf1cdc5c37c53573c017540c400c05c040d51044d5c300000c47fc737730333404310cc0000010133003cc3c0010330000050054c0040d3000f7000c037304030000ccc03300c0050350f004d1c414144f3407700000c0400c30101301311f3430c03030cdc00044400c543c333f10c11ccc0730700304cc41d030c100c53d4400530f40705c013f3f40001c5030c314cf00c0d0f400f070c01cd11c400ccc0300031031003c1500f5d00341d304303c0c3007c00f0c031004d30041003f10003005300330dc0004030c0575cd0400757f40cf3400c0345c00ff0c4400cfccf00c3003dcccc030c00000000c044c013c444000043100075f7015d03f003430fc33cf001134f35c341040c074cc343003c411c00c3c0004043000cc33005147000330000cf0000c003f103f5c47070030f441ff00c0ff0c3d10340030010470d10f334000013334d0c13c14c0c3c3f3d000443c43c03004100f04c037304444c0000000cc10030000030cf0c01473541c43433fc4000c040040c034c3000c40c110400c3013c0004c3000470c0f04073c3430001035c0c00f513cfc7f110c05f370340150000c00c4000c770031c4004430030433000f0000d574001011337410c00c140011405540043d15000d300100f104071017431347001f433cc333003000550cfc0cc1000f00c0c01300001c0301cc0c4340c000000cf0ff10c50c0f04d3003cc40310450000c0000f051044350f040450000001c1cc317400403c10ff00cc01cf0f0ccf0c0dfc301004dc3c34700c00d10107101cfc003c40144c0c3000004f150c0c0317004010003c1000f0001440100c74000130133fcc1505c43730c03c3c0000c1f300000dfc440f00007040031f310c0f54130c15570c103430c1c0fc1f11031030dd03f0334303011c0337443300703f301c0c40;
rom_uints[424] = 8192'hf3c71100f3070005c00404414c0fd04cf3f700cd1000c04700c00f0400d00311c0d04034c0f4c30040cc0134000173cc43f0007510f01cf15f4730dc3c070004303334f040c31c3f0c0070c54000dd0c04150010cc000dcd043133400c4c00003c75c000003044700401010434003c03701c3d000044d4400c3c33c030005500f045dc0f4004003f4c0010c000041c00c004400000300040c0c30c0044d300f040134331004170cc370cccc0111004400315c003000004f37504c04f33c0c001dc0040d007007c00c400010dc1c0c1400017034c0034fc34ff005404d3f0413004300014403cc15104c400110073d34dcc000c5c04000c00000000011440404c03300000013000f1001c013c53c0000cd313cc0c00043c401533333703c30030053c0400444d34030c034fd741003c01cc0400d3330040304d03dc1c304c303c00cc000340044f00c1040040c0c000001f011c7001310fd0dddc45d00c004c3430115cc0443cdc31f0c1f034c30541d0c0cfcc0c00430440c044051c34c070100000fc440030340303c130dc71001000700c00000c00f03331c50040010440000fcd400040000c010045cf30013d4711170c0003150c000fc0c00100000c0407d03ff3c1110000d00400000cc0000001d4410cd03044dc110c304034000d50f041c013cd0130c4f0010dfc4f40111f04dc0c10700d04004d017400040c4c14c73100007f30d0c13f04c03c740040cd000d01d0c00d10c3100f103c0c300141c001fcf10d1c050030c03f53300444040403700703cf303704c3c40111050073d1c0430040f43000c0c0cc10ccc75d41310f03010cc1043d40004104071f40c0c4d141003f0c0d0400030f0c0041f0cc04cc0c000003507c0d0007fc30d44c1c010100400014c100400447404d0130ccf150c10d0cd14103c100c0f04c04004005304300cf0451c41013053d433c4500c3c0c0d00d010401c01030c04007000445340053000400c04040531007c0c11070040003cc0c0c0104c0f00c00d0100000c00000c3dc0414000c1dc10034c0044c0c1d3d500cf03c0d041443c3140c0030c1154f0404c3f1c01131000000cd01cc70003401735010c33fc0c0c3770030c4555c0d30c41d4f003033d0010403300c1300433400050005c500c07c000c404c0010010f310303100c4404140c01d13040000170d0cf304f1dcc7c03030ccc415c301c040dc10040c000d1005701c7c3f44041000307cc00533f00f0507033f0374535003700fc14c00cf40013000030157400dc117304c0370c4303070000003040303c3c1d01100407300d3410000300f15c37330000c003103c00d0d0100c0c04704030f00407041c00740d034030450dd01030f300404d07d0f013c113500d1005140c0c0035c053fc41000c10c01c00d30c00d331cf00030001c130c000;
rom_uints[425] = 8192'h4110400c1100130001100400400c30044c700030417c03c00c5000c4c000700001c110ff0100000033c00c30000543c4c0c00cc331001cc3334001301400c00dc01c70c041000f1100004c05c00d0443c4001cc0fdc04f40cc0077104011000030f0030100c0d300143050344033ff30005c0f01c1404c71071000c30c040130071f10001010c1031410030003fc7010100010000400043003f013131333d050037074001c7c31c03030000cc1cc05ccd7030310030030700dc40574070c0000103300005005c1f0c50001c00003300d000440113007340504c0070df0f100c0d000070cd0cd04003070c7f4000d771dc0144301300001000000000000540f11c0000004f007404040cd414f70c00000c04cf030317000d30c404033700770300473f00570d04c0c004c40000c0001404430000cf003005004c000c4041073c110c0c0c0d00dc00c000005130010c07070c344c44c00040c3c30d00c707030354100df3df4d03003c10c70f0d0c4d33330343304004d001c10011101c010501c007104000c31301174f01003d111411cc0001f1300c04000001400d1f440005f0010c0d4030003000400cc510f1031cd00040f70c40100134033403c0cc37000300030c40000043300000c00f00340055410c30030040014d0c0c00000004ccd30f30cf0000300c01cc040000000350470c4104303c400001000440010444151c00030c1100d013370c00c400010140010100d40d4000003c0011000110114004c0c3041f44000500c40d000400c7000c14301040c0c70c04073c3140040310c0c543010000000034f00cc4c73300411007010c0103d001035307101d00004754050070030000c413000c40dd00434c0c401430011c000003d3f3500c4f001444ccc30000cd307c4c1054011500fc0c3310100c0c41c50010170000000fc1f01d0751040030400114cdcd30041004731300c5000000540d0c40c001d0140041c001040013000c3d41c00c01145c71011c04cc0000c10f10c1047c0000c0770040000c00cc0010100400d00c4f0300c4404000017cc0400c00c0100c01f11400300104044c0430c47c000030010000303103004c303300100c0300034103100007010017ff00c10007f40c030103c301400300130344401007013cc000004000103d01c010c304401017170110c101000d00040030000000000fd30c0cf031c11110743000c1000c010f0000cd0047033000f1c30000f300c7340000445104000300c13010100c7cf07003c434000c300101c04c41300c00d40003173c0d040044cc4034f310d07d070000d0cc0130c107fc3133030010000000c00000c3004103000ccf01c04d303d0c03c045030c30d1010104401000450cc0001013005300017c005405000000c000d00d030000535c3c340040031c030f00c4c030c30c00;
rom_uints[426] = 8192'h33c0330343000030c700c03500cc0c001000037100007000003d0c01f01010c0053003004000040fcc43130100c0c0704c100c10f111c30004c100330000000030d0c0010f044cc0000d4c00040c1340440340c734c7030003d3c0030c3010000000f00c04000303c34050c31c334030cd401100c1034033007000004400d03303c000015000040010c00c0c3c307f000fd000100300430fc3d000003001500010cc3030015cc0513043c0401c113400000f1300004000011000000330003430000c03c010c030c40410130c40101030f10c51003050c0030440014c3c30044000300c103150100030f00030303001d44c00f00001c0000150000d010000041303d3c034000530440003f03d4000300103700001505000114407cf30307d01110030300100340fd0400000c10003cc050c3031040c00040013c07c005045010103f3130000f3430340000714c0040c40000034c1000001103c0d17104040070001f0400000c001000d4054d1033050c001004c70000030015003400010004140df530c01504010d0f0000000130130400030010300000c141144370703c15403dc50c11001010dc000c00c0cc04c0f003000cc0d10417001700c101c0c51f001c0c0310330300300fc71000333041d00304c1d00004004401103001141001003c0003c0c0c0005dd71c0c3c04c1000c430c011710300c030533c031d500d430113110100f00d0cc00f000000d100c0c00140130c1003110000101400500353000cd0001034001c4c01c01001100000c0050333040c14dd3037ccf00f30000c30010051c0c100000d3000cc003f3c10401030d0730d14013017f430000c0400331100000030001f70013041400040003d330c004c01c0400000c01c014470403353001100000003010f40c3c34f101c0c04703000300000000040000401fc014001c0c1400310cccc34ddc100c30c1403c30070300003c3010001f0400110c0007000400400000110f030c03034141070314100100131050c33cc00303c3031330004c303c000f01f415340040c007c103c304c100130500001400411005003117303703001400c0fd10001000c10300301f11001040010001000c0300001013d00d0340c014034040cc0004cf3c1433035107430003c05103303c51110010f00103c400004000010000c3030110000c0c000000303c00f304dcc0043007c0453d000001003104c0300403040505cf00c400d003000010700cc40001300104000cc0041000004000c10100070000304500c0c0f310014700d03ccc0410cc0000d0010f01554700f5030000010500c005005311313300d5c00001d1001000cc340000c11040d000000c00c7c107035ccc00d011f0000fc0c4010000144cd43310d035110340c031130003f1003cd101003141000010433c04070000c0c0010100;
rom_uints[427] = 8192'h30c100300311103c0030103c010c40d30c300f3714df4040030d510001000030045003c00343c40c0fcccfc000001dc7c13000004f400c30c00cd1dc0001c007440d315c005fc330000111430000103c450c17c0c11dc0304cdc10cc10470c3ccf4107ccc04ccd00013c00010333003035df43c040434f0040f030703c000000704510f013c0014001cc00000c0001431040000003ccc043030c30f40401d04130100040c1d330404d3c40010c003140117003000300c000000015d155010000f000cd000034500374730400104171cc050c1400000f31007c1100cdc1f04c40c30c0001f01f003c70c00040c4450c33030cf11001000000004341000030300010003005c0041d4c05fd004dc300030dccf0d104533713fc3530030003d01331c5334000007003001401044101f701c404044000403fc00c30c5300c10414d01c00c0040000c704dfc0c74c0070043103741334f110074dcfd0f0f73401400f0f03f005cd3004001d303400040051510140c1304c41c101137c00004410c00cc4300d304007350f43340000dd434c130c40001000030737c0000c0c4000000130cd5f54d473000000f0d034cc001cc30dd1510c003300033100170313d03101c34430001c330c30110c3410010040d30444010f4c0c10d300cc4c3000f300fc07440010d3400f0c0c1f0343003433441c0c537d00cc034000c0c0300011710001000c30c40303133004c7101c070d0013d00000331000133c3101301c30c54001c51f0d00c17400030103000f3c00cf0d04400000044300000100c0100030dc510c0dc30c50003350004f1504111033000f1c0004cfc00410705440d000013c010d3714d0d770400d433c01103101c000301500f00d00100c770f100030c10000d04740300000c041f41f1f0c0003000f1c11000cd4041f0403330f130fc030430d0337f03d30c300c0f50110001303c031f3d301111433441cc7300400351c4d4030101400300cc30c000c003d73c031c5040c30570c0dc003030d315c030f1d000317140400070c0530743730011f041f044f3c0400000c0000c301003000744001003114c1410000003c0030c0004c01000c0d117341f0d00141011c345fc013c00c00f14000c03c000d01300c0d00143c0400000c0411007c3d3cc410d31f00071cd700cc0d0000340d00d00030d153c31d300c00035f54c40310d4533d400051c3d00000c5331c030c0000340004173d300701157d30070014c31c30017310c113100054000033040cc100300cd30330c000d0410c1400033f1d10c1cd314147143013c4345044000001dc01c000cc00c033000c5fc3001f00411130703000031003c074500c400ff033cf00353000111c000c44d0101700144030000fc030cc03c0f334ccf55c300c03007407d000c01d0d701fcdcd31131fc0000000;
rom_uints[428] = 8192'h44c30d700003170500003f103071cf01030c031df000dc0013d0dc004cff00d30313c7c5044c004430dd000100c0c0153ccd0400ccccc30f0c000c11310000000010030030c030430300045fc1043f0c00c0010050c400c0043000000c0cc103310003471300f410d350fc014c51f001f7c00005c4ccc3c3014040c400330000c33033c050310000000000003100c300407c0000000004030033cf304001dc300d0c034c00000f1c00013003103c43d300f4cf30000340110c1000c534040003303f301c000013c0000d00d700030dc403030f000310030c41c0010030450040430c400cc010d30100044dcdc1140000013130c500730041010004c04c000000d04307c01407400cc035300c0100110111d3d0c4c140d3303f033003014f705c10f5fc00fc0300ccf400f003f33040d0441c70030540100033103100105035c413100100f00001c0013c30f0c4050c13c30c0cc0c0034c0fc30c5f001001d0c300000003c3000c00f0c33c54cc143004003d114300040c100d0c530c01003333305d103c33000c5114c07700c010c03c0c0040400000310010c310c4400000c0100510330000c430c0400c004340cdc0300040404301340300c0000f117c330140c03311001350cf003400c01000401c40735c0000f7c3c0004d04414730010f300c50c140340504c0ddf003f043c0103100fc40000c434003030cf00040335d131c0c340ff003c10155dc73cc3011c303c00c40f0c0451700dc10cd0c05c0010041031c1303400000c40d00330007d000330100011c3cc0000010031000000000cc0d300100c300f000100437cc014c051075fc0301c00003153403003d13450c00003003c407030050400000f0c5f3c10301000c40010001c730000c143050f00000100300010300cc03c0c31300c31001d0f001d34453000f0000100c0ff000cc1cf01f03070130cf0f300303740454cc401000c0c0000044cc130c430000c01000c000000104004330410c00001f4000dc4d0c3101031f10300c04cd00d00300004d100cc343000070d0000130c1d0c0c037003004c0001c04c0331130034c101000531cc04001030c4000f4300330000c03d1c5030300cf470cf4410c01ff0100c1d0400100d1f005110c00d0c0c00cf04014710000010dc0100c10744000030c3c1000d0c0cf000f40500103c03301003113440004f04dd0c00010001cc17c31f3c050000c03c1031df101fc04cc334f3141000141f0100c05413071104013d3030300174040334c403730c30340033300000004000431c1cd017000777d0040307513cc4303011030c30c00ff001d017344000c010033000001c3ff0000010fcd40354f0c003c400c5f140000030cc34100cc4c01034045dcf0c00c030003d300c3cf33030005f4000070f000c0000c500035c0c30030c01c00c00300;
rom_uints[429] = 8192'h401044010000c301c00c0c00000000c0f040013000c1001040d40004000fc4c0c7300017303000c000000fc00001004004700000c1073010c0c0c00fc00000004003004000003d40000071101040000000cf0411c30000c0430f40404031300000fcc000c000c00c000c00310c40044f03000c433d3403000c400c7c000300003c400004fc4004c004c030c00040100001c000c0010c0041d03070000c04c00c000004c30c0dc100400300000000c10003000000000000003400033f400300400c40c0440040043000d031c00c4030c0414c0331c000000040104c00c1400c0d00500100000400c00050043000c3007001004400d000000004c4030000700000300041030300c400003000333004c0007c0000000c0c0c000c103143dc1030000004f000444000030c003130330c033315c53703005c000000000c000c0000000340f01030310c00000040c4031d003010c400003c70013030000d43003c030040f1004070c0f00f40c000040c000c00000000404c013030000d30001003003704c1030dccc0c1c3c0c0001c40000010404004f000000040c4401010000000004cfcf4003cc0300703000130000000000f0103d4cdc03003700010d00050000047000c0014000c0000c0d0000c0c040c0030005000005c000430c000c0cc303000c103403c40cc00044003104c005100d0330f3c004004c100430140303c0c0104010c505c0400000004c3000105300014043170000d00c003000c1f30c0f300043f00071330000003dc0013000100070c130044c100c0003f040040000c414003c07c400007000000c00004c0004003000000000030000c00c0c0c3f40c004000300000004c000d04c03341300000c04c440d010333404035c00003cc03040c04dc10c0004000303c303704c0000c44d335c0403500031000cd400c13007c03d3c0c00430fc4041404073c40c4000010000d00c3c004003c0003c00005403300cc01004000000c030c0c0000c0d40c40001c7030000000000c044c3c044c01330000004c30140100430c1c4dc000034000f00dc007300003000010c0010c014c3004003040000c4000c7c304c0000000d0303c40fcf7007000000c03004c3000f7040c0133010030430000c010c00403c0540d0143040cf040c0c143000c030c070c03000c1103040403004c3300c00f044c4c0c00000c13400430000407400000300301c400000003c4307d0040000004c33000c10cc000c40037c000053ccd0c34000000000c3c04400c004001370004c4104c107c0040f0375070c0000c300000c4004c50030000c040004000f000c00300c1c0030c000400003041c40c004000030c0c3cc340f0030000c400000400000000c0003700100040001c0030000400c0400003444c4d0130c000c0031000c000f0c1300cd00303dc40000040;
rom_uints[430] = 8192'h10d000cc03100000703300400c04000f00111111df30430011340004307c1403510403cd00f3c0011cd31100d0140c1370300305400400103c0307003f30cc0411f040314000415400000c5500037dc0710100cd413c10f03307cfcc0017c4c000704511c7d1300013304c01c0033c030c000000d040300100f05030c31f0441cc033043511000300cc10003700cc0334404000300c01007014c0340f1300307c4cc0111040c4710fcc104410d13710000c0301300000dc05f0000c0c300000100f100140110330011330003007000cd14017300003000cc301300d0fd1301c3414f00030c0d0301d1cf0001c004f0100441d4cd33d10010011400c740000017003d111301c0077530104033304050f0d3fccd00007000104c00c01cc1030131cfc40000005c410000000d3c5014000f044000c4c11fc0030cc1c300fc04010030103000100d0d00300f00d00fc100100303c00c00cd0001c14131400040c0c3cc403105c34c0c7003c101040f3c33c0c013c05000c040cc035140c10730503c00540040030301c003010000c30407700c000050000005040044003f053303f0d3001f0c030000170030c10000143003c40000cd5004007544010330c40d30c000c0c0007c053c31cc310300c00117d4343140013030c030c0100001751300010f30041f001310034c0f3d000050000300c13c00033f04d4410300000c00400404500033c0710033000ff300f0c0003c7104c0000f00cc00c11303cc031140000000f030c31c1341003000000d013c0c31c300c0cc4030cd43030140f000c1cff0c33c40140c0001c400300031100c4500d4300003411003c0c103400000c301f4000000f040000c30540fc74004c03014700303005003f300c307c0c4fc40040cc000043c010000f070034c03134010cc145310444f7cc00001fc003c001000c00c00c10104d014fc15470107401403ccf030100310000310f00443100c0c00d04040000c00c1100d04700c00dc005000307c1f07fcd003011041c503cf34000400c0c405c304c400440dc000d0c0000031c114000004c0c140004cc0d3000c57c00000404100503c0d0000000004f00c70c03fd3f14000053300c03100501170100004cc0003c100c140304c010c00c4c013031030c04000070010c33043105041403150cc00031041713057000100c00004d3c0d13330310d0100c01545501000c3dc1000004c37df000304013004000c404cc0ccc4c0c40440170135cd11f000c3300c00c0004500003d3c11fc105340000d00303010c0c1d334ff30003030000cc10150704000c0400043c07c3c01fd0c00310070c1c0017000001c130000d1707d00740c0f00051351010f010037fc0400010040101f74c570c330c7001f0f003010544130050000d0f04010c453000104c0c310c00c30c3554c000000;
rom_uints[431] = 8192'hc5014000c011c300300441404c400113010401c00c0c007300d0c54003000c131314173107f700000c03300001000c10c00d0000010100000031030cfc030400001c301d00130c404000041447404cc04f0000dd0d0114c0430040f30100c4c0014c11c714400cc00707005d143003cc0c1300030cc34010c0c300c300410c007144000c00c30040371100ccc04000cdc30403440013c440dc0f0000c30300c000f031c0cc400c01c1cccc00f40040c441104301000000f00354030d0cc30004c0044704410014f34f1000c3c3001d1000050f4c170700070ccf0c03cdf0100074040030013101400d11cd04ccd3300000070c01030500000000c31303040040cc030003c34c4f000cf00c014d5c0c030cc43c010003c407040000c0000dc000040d0d00c7140000df03014c030447c0c30000014300000000000c40304000001ccccf1300010cc031c0004c00c141c404500500d004c0cdc0c0c7c40c0c0031030403100700000c4d1444413007c34c01f33101030c0700014077c103c00c0dcc0110031c0cc004c4d00040c300c70c31000311c000041354431f730014040c33cfc0004003cc4cd07000000d1544001104c10310c304c0010133c0170c0100450d710c000130400403c00504400400c10300000003c004007c00000cc0c30d0300d13300c0d00000114d0037cf03400c011000c430c30c170000c31c0fdf04c1013703c10cc0df4c40c1300040044cc04000c10f01c3045c030fc00340c3003d0c3cccc4440313014f03011003cd000d37040c51c541c7000300001001c3c450cc013c0003cc14c1fcc300c1070c030011c305c35000410c0003d0004043c0174101040000030000041c0c00c4100344030ccf000c13c7013100d0cc003f15033d0c0000c43c73030004f0ccd40d00070317cc40534305c00103004000000c03cd10dc001300051103c70dc554103f57c0d1c5040044400303c001000041430007000cc000430000000000100fc0110010c13f3403c3431100c031000c0d0000000000000c5043000500040000001100d34743003303004040030030103100c504c000c41000700dcc034c40c000400350303c400030c4004130c14700c1c55d3c0040f00300010031c00300cf100c0c3004430373cd0301c04cc0034740000f30004440510013c304410101030700010300f1100000fcd4000000f0d4c304f0c4c1c34437004d040003033c03fd00cd04030140030d0d41070040000fc3000d0013c0d5d30400010131c300d01c00001037c7c0014cfc1040dd170010000cc10c1000cdc410cf00d010f105000d0f0001404ccd03cc0f000001000cc1c30f015c301c470c303300003471c4440000530c4f00000cc00044c00d01cc070f7c0cc00040d0010003c0c10303d0310303c3400040100004cd1c0c001400300c00;
rom_uints[432] = 8192'hc03741400c003c4400c0c0cc7f00d503cc00401c500014030034c0c074c74700c4c0c40dc14f10c0500304c150030044300004c400c500c10c0000030f304001344c10f500c00000030000175500300030031040100070400d0100f0ccdf000cc000300ccd04c000c0c0040c01d0f1030c44dc050c00400700cd4c40000c700045f0fc00cc3000000c410000ccf001001000c01d00c010cc7101000cc4014cc000044040c04044c3c5400300d01404d40004040000100504140104403004430007c300c03010c0135c340403f7c045cd00c0cc03c1c034d5c0c100c003d13103c300c00700010d00430500c74401400404c4043d4d3010005d4010c000c0405ff4c00c0f000404100003003c0fc030000714c4c31411f0c4034400340044110000000f0004010000c0010054d00034c00c30003430404c300771c41104cc00007d40c00010cc0c00c70403007040004740030c40003d0f034c0cc3d100503700010d3f00c10cf703300300041f0fc50040400401004700f0150dc500040000005c000110011c00000700c000f4c043c04003d4430000d5c00c051c0400d01000dcc140000f3c01c3130c0d0cccd343000010001040010003c330014300c34040005307044c000c4c3033f400c40010030dc0034400c077c300d00c00030fd4f00c0040c0c3010f000c40445440141c0711c043c400c70000d74000001fd01501cc0404c1c043c001005334033c000c70cc1003111130103cf054004cc401cd07430c5040003400040333000000000c003c7dc004c00c0304cfc103c70c00c1000740030000004304c31c4710c470400c044cc4040fc0000303c000103147113130000050f10404cf4003cc03403070f304c00000340cc13000441f010c000c30c50f0f03370004f040ccc1c3c3134f040300445440c70f00001d30007040d300f070050004d04c0c1d00cc30c30dc14105cc0c04100cc40c1300040c140003c301c3c33000000000f3cd7003000407300070ccdc0c0004c004050773d401c03cf0004000c403440d00cfc40044c4d1003400c1c0000000000c0040d43450530003100c0430c404c37300010c0047010f003344c04d0010001035c07cf0c003c57c030000c0300001000c00001000100d0073c30000404100030303410004f31301400300c0cc400000033440c3d3017004c400c04cdc0050c00cd00001440000d071401400d000000f3c10c40c00c0003ff0c341c1405f10000430c1ccf0040000003407040000300010000403f4001100c0c307004c0000c5c040c033544040c4534300014df0c340441c40c34043000034030f40000c40000c00004343170440c0f3000340340c410f100cc0331003c00c030c34000cdc07014400410100fc3c1c0000000013c00350d10001041700004c0001001340f001cdc01000c0c000;
rom_uints[433] = 8192'hc014033313010300f30c03c04d04303730000300301304cc03103104437000c7c3c101c3407f0011d31704033100c004413c00004100005f3030c000030010301013000c30000100340054031300000000040005110043c1031c040703010f03113d07470c04030003033f151013cc001040c10f0003010140c3140003f3030003c05313073100c1000000110000003030c0300000c1c1003100010004137401c0133101010003311301013103300330004c0f0000303017300700c007701303010300110000137c0001045000303dc0000303f530030300300001f1cc430000030000303c0104010013003d47040ccf713cc1101033000010c1c130000030000400030010ccfd700105031c0010c4000cc53103103007f0034000f4d340010c1000c000c10100c33043d00c00c010071133043173741001400c4040000c0100d303c0040110f1330033301304c00034070010cf030c110d130071c441450003c00d31010000400f00c73001000f3517404041000f130701cdc7034c0010310c0d44ccf1d37d0cfdddc00d4300f55f01000000100003f1c0033300d007000103430400300c00c031c00003340301cfd000730030c0f0c0310110103313003c70c03101c10c0c330cc3310010cc0003000dc0000100003f1101004301003740c413c300440310000f00c7003c333310034043310c04c011c5000000c0000100c03000000ff3000d30034c00401ff3031fc3044103301c10010300030c4010c001311f0c051d0c35300300d30000043500411343c000001c130343f40c430000175cc00103f00f14300104110c3011d04dd004040000c00100103dcc0333004044033c3103000f3fc71444c100343c0cc3100f1050f044300701c00000010f4cc1c37003000f003000133d070407c0c000003014c101354f430034c00000100001040c4000c4530c01303d011105c301f003003c00300d40d0d00c33f030010043041c3c0c0000000135000000011f00c403414f00431001130000303010040010c000000c0100100000303041c1500c003303003500030000004300c00003000001c043c0c13500503f4330c000010010411310441d100770041000000000040007030403011c000000c0000400100104c1004005310d7c00114007c3f015300035c0050000110704c000c100f500430c33050170f41fc34ccc0030000f010101c0035340004000034130000000c13cc1f0000c040303010511010000000cc0003d0004c33f00540105f0335c0135cd103703f147100010013031c700100c040145330430310733f00f0000003443400c00700003d104000300cc0000c030f13101001305f01333c00f0c1100d103034f0c000100400d30f10330dd44cc7000507400043cccc53c0330f003010d7d3cc004300c5010c00c4074000003c0070000;
rom_uints[434] = 8192'hc000c000d0f1434000c3003c0401f44cf07000501000400fc044c0c00c413010c0dc00f11000f000c01030001001ccc0c151375c030704114033340cf100f0000003f34c3013001310003cc33c0010c010007cd103cc00045c01f330f00c04005c043010301cc0f3cc30c3533000f03cc0000041103300f43001c010f031c0003dc3d003034000f330cf00030100003043c000c0000f0100300041c003701403340c34d3c440374400c04410dd4d0c03400034c000c030cc100010f1510f100c1044ccc40c00040110300110505c00ffd0c4c41f00df3140305c1c350300000004003040c30c0d030030004100303cd000c070cc03c400f050111c00100000311c00c000300043d0044cc003704000410031c0000000f030c0030000c403c0140004000070ccc011007050101043003000004004431010000100cc007cfc5050c33c037450c1f3003001c01700f01000011cf00010100c100053007c404004c13d40700403f04100300430c0d10c5f400430f1300003fc00f0c03cd3000050cc1dd3d10cf07000071000340d00c330c0000003c04000f0c03c100c401c0c0c30fd5f051c0f0f00d700f303c4303c113104c11c0c1c33033450010cf540f07c04f01c314f04cf00c0c03c00001104014400cf00014000c003001fc4c0040140104010f0103150000143dc053c3cc011cc400031503001000cf0003000d34000f3c010000030c400000003fc00f0f003004401d470c00f3cc03101c4cc40003340147315c3c10ccf0c0003cc00ff00d0c0040fc0000c0017703000c340f400401000c0cccf0010ccc434f41cd3004440341100400cd0000040c0c05fd0c741140011100cf0fcc50010f3133c500c15007c3c40d1c00c004f3f14cf343004c703330c0001d0cc0000f07c31300cdcd0d001f1335000104dccc10cf10000cc0033c050cf0fc0c03cc0400c001343503030d1d004f0f0045070c0510031f0c00d0cf000303c000000f100c0f00003000c30f0c0401040340c400433303004330c37000700c0343000100410033c411c1007430c0030c40c4f4000ff0010c117c100c0d0f037c05300501ff140304100000001530340cc70000c00f0c00003cf3310340101300011104004f0c400703c001cc40c0100403430300030050010000403c05005c304d01cf0300010c300050cc0f0c000f030140cf00010c3000040c7341040010371403c00c043fc00001000070000c3030450f314404433040c3003c14034000031ff00300014d1cc5f000001f100c0041c0f410400cff33500313c0070041100cc0100dc033000c047000c0cfc00fc1cfcf00000000c000000fcc501000c4dc71d0053ccd30cc104c0f0300300c01004000c3f10f100431c10104c00cc03030000c10100c3043000fc300000054000300c3c7470c0fcc4050040004103;
rom_uints[435] = 8192'hc3c4004c40000c4c03400cf3c30cd03000f30f00cfc0ffcc00c0c001ccc04f0704010045dcc30c4040000405c40047f010f140050010c000013f3cc0000004000c5133c100fd0000ff0053100400d0c434040c77f4c307c30fcf4d000371fc004005c043000500c04f00f301c3007c00030f0371040404700cc04044cc4300000f03430c000300c44000c0c07040fc50cf4c44300005cccc003c0300cc3c0304c13f4103301001043cc300c00703040001c40d4300d01300000410704300ccc440fc44d01500c3404101004300c41015cc30c041004c300300011000ccfc05d0770500dc01c0c0c0117100fc0304c00470030d00007040c014310000c003004cf07443004400010c035c3f00cf053c01ccdf40c3007c0c3057004f00ccc700100033f30001030c40c1cccf414000c5c0c05000c04500c40007050c030310c004750040043310c003cc00005fc0531f000cdf33f300c7ccf313c13743d0cc0c4010c440c0300000100f30c441d30f110d000c3133c30fc3070c514733c3c34f001fc033cc57113301c4f00000d0400cc4d30040c30003000c40c0300004c1c000033540000f43c3c30001cc03d35400c1030c0311304c100001000f100114f11150310140040040c004c0000003005044700700c10c40cf3000300005303cc005000d30d44c0f45cc34000cc0000004c0c000c0c0000f4c300743c3000f1c104003f5f043d514c30101cc0050000cc0d13014100303c05c00cd0f13135c0144c10440c0030470c4000000c74053003304d0403c0000cc400001010034f00000474c4f0003050f0003f41cc0c0c033f04700043c4400301400c0c444003013700d0fdc0001340303434c3fdf33c3040000000fc00000000f50504c304033c1c01540071f00c0040040cd40040403c3c34404c07100c1f3cf0733040300c7c10040c40c03c0050403c50307c4415403c03c371403c4033fc3303000c0030013404400000f1f00000100c500c0040c0f1330000510310440cc400403c0c000c104f4c400c54cc1113004004413c40c1f0c4110445140dc000000400300c040340c00130430c37401c4c0c100100dc0c0000c0c0030c04c001340000003c0740fc41c1031000000d00cc4c04744317044f00f0040cf1c11c47303c30700700131400000404d04334071010c0405040400070040f1c000034f000f100000d014c0c00070000cc3341003100440100d10c00001d4fc30cd0000d0017d300444c301000c1144f4cc000c41040400104c00c45003403030f4001141c051c1030103f00c04dc4000c4d33710000c00000007c310f3c0d017700d00010c0c000000c0c3cfcf0151301137c15410c00040c5370300040f03c0000000000403000cd0f00003130404f000c33004c310430101000ff30431000300330cc3000f333301000010c0;
rom_uints[436] = 8192'h14f400100030430f311f3041500001403150004c1000000c30cc0031c403000400c40307405c0010ccc00403c10004c3c314003f5cc040c001301301c100040110001414304000000f0050305400030053004000140504c135cd10c1103cd400c04c00300000f0000000100414c03c01c0c0c043303c00cc30334300c010c0300113400c000000300c0000000c10007d0000300c00003c0000073c000030401000501100ccdcc30300000c004433c00c0010c300003313000305c0fc5705cc040040104000000030f40000310400c00000300c00000000104407303c07400000003c401030f11d0c3004000f1007c0000013c00003440000c0010c00000000400003040004d05000100100100d300000f1003000c0c0c7305340004000700c001d010c00f30c3030003301111303d00004d333f33000c1000030134331310334130c30031030450031000004cd3000104c700403c11001000300007000c0000030043c0c4401c0d0c0170cc00310501c00f040300133400000f0400000c00c411d174100d7030300c10000700300f15d00000c030000033310030341c0c000cc5c10000401430440311403c00ccc330f0040000c3f3c100c1000cdd0047303c030c0000010c70c033c0140003000010c401410cc01403cdd00010014700c307300000f400000f0c40f0330003173401400000f004c0c004154df00040f0043c503c0504300700000144c43c000c000c00000001c337441d00f305c40000010000cc4000015c00103000705f330c0003030140700c113c00400744001d30c374dc001500514c5f3000070dccc03d011f004000030010004010c45c03030cc0154001000003d1000310c043c1f400c000c0330140404111000000c000030403d011400700cf000000034f044050530c0d3410cd4030010430dc03c33000014c3d0c5c3c000c5543c4c431003c10f40041c0000c50000100431fc04d13003003d1003000000000000c00400000dc07f40f0f014c30f3334fc540701c3c0c004cc00000005c14f0003c0104001f1003040dc0001030c03c0003c0003057010404f00c005300051c0033cf010300c10303040000c0c00d4007000000010c0130c03100d30004031500040040070001303130040303300d03c0100d17c0f443000c03000c01170d000f0310c30040d10003c00000d31f03040003dd50403301000d4033000004d0434000c40c03c003c00c031111433030303f007f375000345313400c000d0d000000500c300d0540044001f00003c04c400040c3404c300034c000140c3040000041473c0c1000d0d010cc3000d0000f40000000030c000c0003ff330f0f0c000cf041010403f40701cf07000cc300d00c3003c013c71143340d10c00300001cd30001c030d000c00cd3330300000010434c1005700c4d0c0013003;
rom_uints[437] = 8192'h130c0c0040440c53c0c0c1300f000071cf5400003c410103c4dc00c00f153010144c00d40c03300c14140404cc00347031c030fd5f031c1131043100070c004034c0f3300340c05001000700cc000003cc411000311c0c000110073000c3c000400dcccc0f51d00c0000034dc004f043c34133350304303410040001105013040fcc15000330004000710cffd0d0001c00c00000003041100434110005d001103341c0130c1cf300c004130c10d1f03d4144cf430003cd3400d003054000003c300c000c1000fc000c31003d3100f33030c7c34f00c137001030c104c7710000c1c000ccff0cd000303104004174001041430d3c1cd400771434700c00300000f1f40440f03f710c040010331404000100450c0c0070ff0330cc317d47000c5f0c1710003400003441d00000141030030030010f003010301030500d300f4003c0013c370300170c3dd0331d0f40103ddd4c0cc3f013103143031cc7507101d3030c0cd3f50000000010075c103c00451000400000011014c410000c301c4700030f3d03cfc700044f4031017313101331101030c000c340071c1d4003000110c43f07fcfc3c30dc0041c0f00700101101c0f0700530000043000f13f0140c0400703503c01000100300000c00000410030c305cc0f433cc00cc1300c1f40dc41403030c04345f01000c004f4c000430f4410004f3010100001cf0f04f100140fc3300c713d3400040000343ccd0d310d41030731c3d54cc337ddc4fd000430400005054f3300403001013400304370070f3f33000c0010c0040000c0000f1dc01000d0c300c4f3010070c0cf0c1c30c0c00f53c40c03400405c4137f00010003d0000cfc3030153c7003055c1007c701f0400000344c73000303f003d0000033001440303cc000001c4000fcdd043f0c07001004c3404cd000100001430c133317cfc000004301c11104030ccd7c034dc10400c003c0c03510100070c3000030300f104000017ccf00000070070c403c010035400f0043d504000100c001c17dc00300400403ddcd01ff731001700cf0c0073140001000030043cc7dc3770001f707d707ddc0011d43000d40000001c30c0001070500500000c0cf033010000c00400cd4300000033c0043401070c10000100f0401103005370103100fc3007011703c03c3dc7d0000c000fd347d00c043c0f3053500313303c330001030cc100040cc0030c1010d3303041500013133314005001340c51f03c000047000004710c101cf30070001f040cfc0103400cd0c01c000c000030f301d3c3510d3c1003034f03031d3003f3300301f00000fc0034c0045404f0433030c400cf0c00100430d33400c0fcddf000c0050c540001000cdd04000003ccf0334003513000040000d000c3110000013c0030007411000100043071514f717115c1c003000010;
rom_uints[438] = 8192'h30100c04c440f340303013430040cc00f1001000c1111c003c03000c30c00000000f033101011070001c001c003111303f00c3dd31100c1004c100430c17010404c03003010010000000c1d30053001cc5050100000000150ccf00007400f300103473013714c0300c00070154000031c0405035f141300150c014100400010f0c000ccc03000133010034074000130f3000000000301cf0430000543130010cc10c300c0330f330c0030c00df1004000d0100000c1005cc0c01301d30000054010c000000001c070c1100000c0cc03000010f003400d01c0040303d030100077400010f04f01c04030cd0010131030700c314f074000d3001000c3c10000301370c0c1c5004000c10400500013dc01c1000c3004005033fc304cd15054c0307f01000f0703010000107040031310100013010050f1000031c0d100107c40000010401c10ccf00000000c04130100c7d003705f00700d500300f03f0cd010000c4330070471cf0c0f0f0500004c44000040007003d0100003370040000c4033701311034f0310000f137100000034f1c001000c01000003341000005df003000f03003033c010c0003c041000304f101101107c100c00fc0013c03044cc400700c00100c305051300500040300003c03041000033404c70053110c54010c5c00010c0c0410400100040010000c450dc010c300043c03104d0010c0f310d005c00000130c4030cc04000d3005134010c4001c0000000034100c141000013d000c000cc034740c000000130000010000043400010030c40403000113d00435d440041173000001700007000c0171c100007110500050701300dc3005303f44c0000000c01430007540c000000c0cc040dc10d1317333c0443c01cc0cc4104347400c04000104000105c000001400443c10013dc03003100300c4040340003300733000f1043300100035c04430001c3c04014cc4c00011cc3110c0c004100f03350750cd00000c3403c00010000000c10033054010030c30f501c01031305f07100003010500c13000c00c04f43c010400c004300c0c11000005414c05040001ff044300cff100040300405d01c310304104000004004c000300100134100dd33343000000c044440704101f3030cf0310133300303300ccc1000c0c00440f00004000070c34301000000100f3300400031003300010d00003f404430001c0c01cc00011c010001c1f000000f0000c0034c0130c0040401f004300110c04040100f030303001131300011000430034003340000037301000330c0d40d413003fc000310f0c00c40c000004f034400000004f13411c00003000000000153c0d3000044134c130303c0d135000073310d4000403030031cc0c0000c000033301030f05000c30000110011000300300cc003c400001010053300c040400c0f01000;
rom_uints[439] = 8192'h400c0c050003001dc10c0c434001000d330004130dc030000d000000f00c404004c740c0d00000004000c1cc43c00041300040c1c103005001c1314f300400c0000000110300000f000305c0700c0c0400c0cf45f1040c30c0cfc0400101c17fd10107c4040c013407c1c501c700cd0d010c03c00c300d30000003400fd0c03530f040404040000100c001054cc0cc4100050300003f0c0344c30000c5014100410040014c0c05400c0000140000c300c4000c0000c3040004010d4c45c0040c00c3c701400cc00040c14f11c0cd0001440c13440414000004010000340000c4c40000000c40cd010110cf44c0c1cc00040d004000400400003c00c0400c0f403703cc070c40c100c303c00003000fc0400c03cd0d04034410000c300000c4144c00300c00c1f00c10ccc103c0c1f401d01035c0c01c0c03c00f4404c45c03cc43c0c4004140300100c40fc00d0c1d4543cc0305c03005c1c04704000d0cc3c030f0053303c1c0040400000544000c03054d43041c00c0000144040c00414040014103cd400431d003c10cf4c3c503401000010c00440007c100030cc31d00730030c04400000c40c303c0404017030040000d04c0010d4d430000c007013304cf310300c130c130f0c30040c100c044c1c100c04000c0c0010000c3044c00730373030300001d34400104000dcc410f100040cc43000f311c0044354c01d1374100c34c0001410c0c00c01000000cc50d400001dcc10d0001017c04373100c1000cccc004c300400003c010c4c000cc434c003000030001400040004c03050101410300000c43cd4c43cd0004c3404040c3033f010c0f000100cdc0c0004001cc000f014000c00441030d00010000c0c30fc0c1c00047c0c003040101c144000f0400304400404301704140400100000410404c00030500c3040c00ccc40000cd05cc010d0000014004c1cd130c40f401c405410000f430c000c000cc00044004005fc040000cc007c0c101c0c00000f04104101000c040730301fc0f00d400c000cc0031013fc00040cf10010000000303051003000000c101000300cc0c07d4000004cd00000f0001cfc000400c01c30d00000cc0cc404dfc41c4c00c01000f300c004000c3010c43030000c1cccc30c14741cf7c404dc0ccc000044750100f43c0304c04300c40c17ccd00c41007000103100c1c0c45c4014000010c0003300d00d000100000000c03cc4c0f000000430f03013d4fcd110104034011cd0dc0c000c00003c00c0340c04001000c00000434c40f00c000400c010500f40c014cc0cf5cc3d5ccccc3000c454c4c010c0dc303c100c14dc0030c00000c0dc1c440040000c073c0000f00007040c00cc4c44d3007c0c00044004031ccc04c004144c100c00c3001300150c440fc00cc33030100030cc40d011fcc05c30003000;
rom_uints[440] = 8192'hc01cc00001001300103500c00c0cc144403000330c7043400c31c3c00c3130101054d041505450c30c0000010cc0000030c40403437400cc170011c0c30c11000c4050400407c003000000c15301c017c0070301f1034103443300c3030044c0cf51fdf0500140030cc3c00c043303300c1004045343540c035f501040ffcc315c3c430310c1104400040003c0c001cff3400c000000c0c00d400c310300d300c01d0004dfc001d47070f03000c3300300f00f0000004f71d010315c430403c5103d0cc0f1c0004c00301f034001303401c103d005100cf0541110303dcf50000150c04c100fc3f00d0100df31074c03030c01040403000004105434540c0003100c00100003f000000cc33f03400040c3104c1453407000c34100104cc0000000300d00d0003110370fc041f0f031343300034371000f00c030d0c3f4070d003430cc010c0c43000003f113000000034cc4c041440f007411f1c0047405004c00c4303114c5033330540511000c070100030c30c4505000151c0101000c05fc31005500044444003300c10030000004c300c3c03300f50000d00050310c14033340c4030c3100004110350013cc03030d4071431c343403330000ccf30040f1c040403301c50c41110100c0f0f100dffc35c130005043f1003000400fc00f03033c0050d343304100d0c140005c07310f40cc3400fc3303c1cc5340000ff354f1c30143ccd150440d01340c3c37d00c30c4c30310011c010c1c333ccc003500307330f7005410550003f30c0100000103430050c0054c03003051c0f10000c1330c03c30c070cc03cc30013014100c05300c310c013101000053101f5405c0d514f0c005f705c00450c0004f0c041044000700033c017310c000100c304c0fd04c300c010c10003503154041405c0f0c03314d000d41cc00010c004c000c140404c004005c40d01d0f13000f154c3c00030f5c1004150c1030030005350c1c04000030100004003d0100f0140510354400475030300130730f03f4c40300f000000f0005000113000d71040044071f730040030c0030000c14d430d4f00470344c00c3141f5400c03c000d00040010004300c0c40301c0000401005010f1004100f0040cc3f3300c0310407f0005003400fc040cc030050ff003c4104c13000ccc00400cc00104003005c0cd000f040c1cf10cf100f030ff435051040f1f50100000c4d11100c0fc030c004f0400f0070440fc4445541cc003500c0c4f0000030001300f10007004c000003c03011c7c004cf5013c043033405fc04000c40c3131030c3300304f34000100ddfc0000000f103314c00047d0000c7004c10dc0000000fd430c34c1ff1033310c40c004000000f003051401100c000c50dc0f5c00300000004fc0c0030303000f5000c401df4c154400cfc005000130133c00000;
rom_uints[441] = 8192'h73100443cc04c5c03431c1100071103c0000df301cd0400074304343dc43c30010003f05010010000f3df1f000f4c0f30070404f003cdf0f70100c1440df000c05404410443040440031314f3d110c3040300040f10f00c15c3c40034d14cc00d447f4c30c00307c100104d0f0cc00c0dd00150003003500d3c0411f340100fc4c31733300000430403c00100304c0333304310000cc4040c30c33c4c3f0031d4cc000cfcdc03d44004403000c0d44004d13400035dfcc0f0400fc0cd013444751000f3f304700cf0f13c40f44ddc1400501050cc143dd03c301404504100d311d030031c0cc104403c0cf5c34fd04d040c3c401df010003033114444000c054f110003c4cc01fcc34cc113010030c40cf033c001003343c0000430070cdc00f344000cf00c000dcc0c0143d0c510d030004031030000000744d003001300cc041000000f0c5030f1c3037740400f000d3001c341c00c3d0407431c0c34d01d3033740f13411350cc0000ff00c0133cc003ff000f3103144cc01c313c0010030014700c03500004c1143501d40cc353c30cc00c0c010103c10c00c4cc5c0c0005fc4ccf0f10044303c0340037f0f1c70c0d0cccdc534c40400f3501fc00d4d01400350410f311033403d0fcf010500341d4c101135470c000400ccc00c00f0010074cc0df40cfc3f401c1f00d1301c0004000403c100c311703c00334cc105743c03044711041ccc1c50314ccfc111dd30d030c470050343fcc00f4c0301dc004003c003ff0c0c4c003f403730c14130cd001301474100301c331c1040cc3000031f40cc30fc1043f0400044f31034033c34007cd0fd004c5d3100f00fc343dc0003030c10c0c0cd04f0dc0c4040fd170053cc07404000f4440d11cf00004fc07035c00c440c703c37c751014430031c1cdfd03c03c0cc40300030dc007000fff00c1440313350c14053f074000040dc04543300011ccccfc31374c0103700f1440c440000dc7500304475c030c5c00000f0411413d33474104005001c10004300430c573f10300000d10100101400000110303047040c04c1c101045370c0c400c0000f470711700001311c000003f00c0000c044f1174fc3404101dc3c03130303100d053003c0734ccc00f43100000dd404300f7000cc3010430f1f30310c3c01c01f40d0100300000044cc0d3040d03075300003cfcd13540100400f4007c00cd00c7d04c14000c0d031007700300c31ccd0c17c400d3300700004c5130c0cdcc07f0301cf000700cff70003cc030c33110f0310cc34404fc51c0004717400001334dc05014013c13f414cc03c00000c334c000d0c0030c100cc44cd000730c0ff033cf0730c31d4fc33c131003cc00703000331cfc0041074cf401070cc301000cf7000c34430104c0074c0034703100c0000cf000f17033000101000;
rom_uints[442] = 8192'h313f0300c1f0000000c0310df104ccd4010d01704fc43c1031f00000030000510c504c0cc00300030340ccc1401c4030f300100170400f300f0fc0303003004f1310001100c135003000d0f004c040400001c13f7471c000c013d04000f011000c40041c40000c33cfd7dd0f344f3c100f10c000130c33c005c0000c01c0700f0c30c34c1100000001f003000f00c0430000c0d0010f0c0d330030004300300c0c304104041c5330c040c405003f401441f3c0c004003004d000c340d0c0000400c00c03300c0401c3044004c4cc0f01101315c05300330050d5cc1f0d0d0f70cc00000044400001c01000700df345c540011d1c50d0000000004dc045004530370071001000000001434fc0100c14045f330044100305cd30c3cd71ff34047040c0300f0100350013fc0fc1000043c00f01015000444045374000010f00c1071c70c003410d3030c000001571004030333d3c00010003304107d000305374100c400000d007740003010cd30704d350004001c140000400150300f01404d0303030010f15d00033700c0103c07375c070000000300c10dcc00c30c0c003c004f010030c000004300c1033f015c03c3c0003f3000010000010030cc040cf3c30c1000040cc4fc33c0300040c0404004c33d0003403c401c040430100c031c0410f307c44d540d40041330c1c1304cc0fc44075004400c034f030401440c4cf30c0c010cc17c3c30c030300c301000c3070c3f000f045ff1000c0f0c4cc03c7f040f003304f10001013c5c005c300c0000cc0d0010343d03cdf104d3f00000c730003010100114007c100701cf03000044345cc0003111100cf1004f3c0001c0304d04c0c3004c500103300517000000004c07cccc37000c051cc10030c0033001c040000013403034c000fc301c5f0d0041110003cc40d004010c0033044000330703010000001400ccc0344cc7057c047004c30040f10c0115d310f511100cc4500100c000030000c00000000d40c000cc33c40cc000f1d00303040c000710000013c10304c40000dc30300000003c03300c7c031400001c403f400054040010c0011c0001030340000c040000ccd04f04400411030000c00000330007c3c1044cc331040c4c00003755001c00050001003c17c0f3743170000c0031303d0c14571c000d00c0000340c704c0cc3003003d000000110c403d000f0003c00c1054000c04d110130000c4003000100054374300c00030100d0501000400001c0c3770c00000000d040c530434030fc0400c0c40f334010000c0f1c430c31300c0c100101041c4304000000034004000300c00540c00047cc170003000f4173c30101000c1c0453000030c40041fc70c0340447c03400000005d00003fd0040304014c351044030c1f0054d00000cc4c34d7500010000004f4c41c010c00110404;
rom_uints[443] = 8192'hf4000100310c0001d40004140c30010f301c001cc37c0100000433000c1c1003d0010001c0300340040411301104043741000335110f04314030cc3c5001440c0077c00c0010010c1400f415130c03f40d004c110140f001740d4010000c0c01c00c101300413700000c034c3f1170000c700003c00f0403001300441400000f050531f30c1004c000c0007104033d73400000c00000c4000f431c014c50c30c403000010000c0050000c00115dc33d4000c000000110f0301000007044c000077f010000d03051f4d4c40010c000003c4f44110000c17030f310100f075cc0010710040010711000c3000dc005cc0d303104c00053100c404c40100f0c0c0d40c040c30000d5cc00300f0cc040c3c011373d4c30773dcd43400004fd7f003c407f7c7007d01000f01004100cc0c100000300cd000c4000c14c700001f044d00030c3733d03d0003034033501500000f430c0dcc000d0c34fc0c1415700c0004400c100d04c10d47000cd000044340400007040c000f3f1003c110331dc005000cc4c301001000301f0f001345007300000040c00000d050f405141043000030500cc0014000c0d00c0c0cc037307304c31cc447d3f13c53400300000011c40004100101400c30f40040030cfc00d1303c41000c404cc74d00d400000d075dc300c0cccc004cc044f40043cc0cc107003110005003553100d504010cc50c370dc0c01fc447400340300f33043d0c0440340c33000107000c000f31017ccc004c0430010073cf00c70034150005000c0430051000c0014f10000340103400413c431300d4cc4000000013c7cc0c3ccc010007000c4d0f141004cd0000f330733c00034c04d3c004150004007f00040007cf4f3c4c0cd0330305d0d033034001d0004705c015c004070c733c003415d4c000c00f000710c30510000300051f15f403033c0d0c00030c304c0c03400070074370cc0c10cc0c10000300c50f4301341c0500000000c005030c00073dc0c3cd0c71001700011000fc0000d4000c40173f001c0c03004c4c00c40c11510010300c0000d50000400110c0701500c40f47010430c40d0d000c040c0c44000140014cf410301301003010cc0100041c010fcf14034fc0000d003030030c111000004c410c017c3004c5cf0004c0100c01c71cc005c00003d30c1cc13c03c50cc00c00401cc704070047000c00000cf17d010ccc0c130c1000010000014c0700000400c4d040400c0074df0c0004c005754c5c000d5c4000110cd0101c030f0100113c00003c034430001c00fc404304000c4f00cc071cc00c01030c0133c700000c003517074444331d3c0f3000330cd1c10003c10100f43f4010c434000144c00c00000150000c00dc500303010c0c000303010000041dc0c33307003431c4010047040303c00fdc0303000000000400c4;
rom_uints[444] = 8192'h4001000031c4d0000540701040000310c403000000c0300040f3c130400c4470014005c041d00040400d0400000034dc04dc04cc43d400501c0001c001000c44c1040100000000000000c71340c4414c443000d40cc0700c4443041c40cc104004f1000d45f3c040104035044c0040fc0010000c04fc4043000c71c30004001174f3000104c330031c4100003cc043c11011105000f00f4000000010c0104c0003000f030004001c00c50f443f00ccd00040001000003c00d0441404c344004000000c400000c7cc00cc0000c0c1407c403c750000000043003c000c3c3f0040c000107c0104755300c0007041c0c010c7000f4344400000000303400c0cc100c5105cc34403c00003fc10c4c0fd31c4f1c03405c404000017c4005d3c31004041c4f000fc5dc030c04d00c450004050c404047d010010c0c100050001f03004400cf0d04000500cc7cd10000001c030004d00ddc03500f00c0fcc4f040001000070d003330fcc0c0300c5700f40d1043100074040040500001450f00000100c07d40c1001d70100030010040300cc4100000101c000c50047413f00000030000c145043f4001cc010110ff044c0cd00704cc030000c4010c70343100c01300140000000001000001050f00cc0000703c05010cc4313ff040070ccc00cc000c0140040cf0701cdc11001340043d0c310c431cf101ff000c0133440c04004f0443300031440fcc011c11001004c4570c1334030c7d001104400c0c03000cc400cffc403c01f40c44300c030c04100004cd044000000340c000004034300004070c731004400401000f00043400000045000c1d0f0010104004034031d5c0c34c040cc00503000c074040d11040dc004034c003d00c00d054cc004c044dd004c4044dcf0300fc33300d40c470034d44c007c4000000c0c014000c30130034c30f4c0334104d410c0004033ccc13c14c47f45cc4100400440514c100c50313c0047c000340c00000000c1c00fd000cccf350c03c500f00030445cc10c0010300cc00c004d007030000440343c3003000310001307105cc4c00c4004c4057c0000001040404010c70c10f01000c041c000440011f000cc34c40000040500103401f40c010c340000310c04c000c03cd07070c0001c3304134041f0ccc0c510474141ccd3d043033005044300f50c1403001041471300c00c000c143cf000d04350040c00403143000000c0c007c0f0030003c444c0c5d510c403001300fcc0333c300c77c45c11004400f0c01301c00c03000040c10c0cd4013057c001043dc000cfc41c0cc7f07300c00001100f30000031c030c4414c0014c00c3001000c00d00c3c310cc4ccd51d444dc403f1004000cc30000c0001004c0d000c31410c004d4c013c44401301c0040d004400000cd070000400430000403000c1c01c0040010c;
rom_uints[445] = 8192'h7500000433001c00f4030c00c000fdc0fcf00fcc0100c40000c1400441010400d1130700d0c1c40000f0000000055c753004740f05003cd00c510003400333100401ccd00c03044000000fc0300c00003c70074f30404040c4c743700700dc7001d03401000c0f01f400c0cc3314f7f501000f05003d00700c004f40c0133004dd071000404000000040c4c0400ccffc00040c000400003300c303000013c1cc34ccc000301007c0d005c03c33300c4c000400000010010c03d00144000cf30004c0c0c70004d303f040c3c1000c30400307131015040d304543000303000007000000040f000ccc00000f7504dc314c34003030000000c0010503c100000f0c370000004c71d0f0c304540c504c00000d0cc000003100034d070000400dccf301000000c14cf0c0100000f1d000000000000dc00f0c300c001001fdc053000140704400070500000000dc003000c10d0144010100c3c031c40434710d00c0c0000f000c43d1c3400104c14403040ccc00cdc30700c100000330f004010540030d3cc0c444010003c040f000305c070c30014003100f0c0440dc400001140c3c0dc004000000010001c300100430303040011c03c0000000300400ccf43cc0001300cc004c000ff304c4000cd00d1744540c0004003104cc0c33c0000c31000007000cc00000413c0130c4030100000c1000001c00040c0103040000040107073000c750cc3000c703040f04000c00703cf07c45000330100101c1c10010d04c3704cc0011040d0000004004d0030c00c44454300d0300000041033f30030300110c3340071c74000c0000c3c0cdc14400005004010300037040100d040001050c0ccc40c1c1000400005c3c0400030d00000d333f000000070c00000014c3c040007000000c1c30c0c10c7077004003404d303c00000cc407003007cc03013c00c504d4c1010f000430dc1403001c40c503cc01c000cc0c0c0c070100070031070010c000010433fc000000010003040cd03c51340c044f001030fc0313c0000003c00f400000c0c330d3000004c104000001330010c003c00501c50c0040040430004d10c103c040300ff00c0004c03050000d40000400c1c0c0373c004c0cc300000300c4010040c04007140d0c00303004c007c0007cc3000d33011f011d0c40010d0c144000c000cf00010f00000cc0030f0300007cd0c3000c10073000000d0dcd03000004c000004c3004c00000c41550dcc0cd0c040004404004510c0c04d40700040c0c004000cc74000d1001470445c0007ccf1000000030004c000c10040c030d034000000c403440343000dc0c03400c0dc00341100c0000010c0dc4100d0001cc00030037c30c0300c000070c04014131c10333c43cd430f30f000cc004c73000c50c0c0440004100007c0c0c0c10cc013dc4cc01f00000c00;
rom_uints[446] = 8192'hf00fc0050cdc7034c041c00337c000c4d1030454dcc330c30c1f030c0c30d03400710cd04040007f1154cc1fc0040dd4f374cd030c30001304d004c0cc30f30070045045034500300100d110d030300c73c707c7400c043c0c03d1c303c040c00700303f4c0cd0c30330044030d030d00d003d4f0140400c000c3005d4403030cf3f3c0300040040010d0000f0301cc7c0050c4000300304040c03000315330030cc1c3003cf010d411f0030d107000110303cc00000f717c03d03dcc3f0c0f4344f3004000355000cc130310f041400100cc3140c300cc0c4f4dcfc4c174034c0070000101c4000040c1c03100d1c35c000fc3d4c130040c040053fc1100041347c4c4003c40403cc0f5c0c10401f0c0704030304003d0c77d000701033100c03dfc300c0000c570703cf500c0340cffc003d4f400c04101000f34300c0c4300004c04400cf00000d1040000cc00d1c004d0c300057c73f0c40cc00c1130cd4c00430000041c04c0070100530403fc500d01030fc1d040c053f7c30400c3404c1d071033505440000c10000c3000f300000c0d10300c50c137011c0147705c053f53440cd030051c10473000c001347030f013330c0400c34c50d03140c101c7f11ccf40f0d100000730000fd405c30c170040400430f31011003000c10df571170c010003c30c003040704ccc170400f0403001c5305547001030001f3307d730cf30c4031c0c01f30c00c40fd0034000c3f007cd4cc717cc0c5c4cf000c34d33440c34dc00705030c031d3003004003fc3000000c1404cc34430c5300f40304c7004c00cfcc0130001c00050504fc0003c10400034030cf7d0c04401fc00c73d00055c10d00f30c0c00101310c0035400410500ffc731c00504000000c0400003d000cd00430f017400c3f300dd71030f4100d0343c0001033c10004000c4150c00717c00000c04300cd3c03cc44d433f73ff4100000015c0c73310010170007153430c0050300303000c000c0c0c0005f3100070d03f00044d1c000cf34f040031050403000540014030050040dc040735cc0c05100000cf000044400c51315033c0c0350543dc000010cc300c003c0f00031401d00404cd330c3315001753d0c00307000c000cd0c00730414400d3c0cf11cfd01f30c3033301440c1f001f300144710401030500fdc00130300fccf010df341341f1413c010040037000100300004000001014cf000401c0c501000dc0f3444cc104ccc40371df00f005150d330141004d34010001c43030c000f3fc0334c014cc03d10cc103c7000cc3f3c04c001c301c370dc0050010cc1c0cc05403011c00c3040003c300007cc13c00300f0c143f4d73001c1c0034cf001c403c3010030004040050c43d351c70430cd340303d03000100cff00f4f0c0f00334144c00000100c170401f034003414;
rom_uints[447] = 8192'hc40f0000c01c04471f100371c3430034000000174400c7010373c000fc33d30703c003401c040c0014d30d015100c0d3003135f0c00340330c040010d7c0c0003010c300030d00000c0000140000c5c001c0100007510004510404fc303031d1445313d1c35c40c030313000c4df0c140000040c4cf0c0c03040c4030053010c0000c010310c00f0c0010000f40043c30400300100fc03000fc74c00c00c0334f0130d30040cc330ff1440071c0d00f0400403040041001f050000c1470003000333cdc31f000301430000d00030c7f00010c400d3f330d40004000cfd1000010c0030000d5c0c01431054cc00000d00c0f737c00004010013000003d304010dd030c00030010c0303c030f0143cc000d00f4c000004030c044017c013d4c04313404f00f300c0c3300001030300011033c010135c00500000c10c30c0c01030cd053034045300c013040331303345c00ccf014104c0df050f300dd11100104c011001341000310000f30001c033001330d343c0010cc7700c410030004714405415c37404400004d33cc70c3300c010c10030c00c003d0c03c0004103f00003701c303003040003c3f533f30031c30f000005d74c0030341400c0000cf000414300040cc10001c10d403c0c0f00410130000033504cfc0f00d4c30131c3f1033d00c01fc0140403c4cc03c7040000004cf0c0411c0007013511c000170c05000300c103c300cc4300c0c010ccf0d00d0400040400c01000f0051400330004c040c04f45c00371d403f01000500004c1d3030100001403cc0734c1cc001043d007d31170f041100304cf0c0407f7c0300000713dc7c51d4110f304d7fc004700100030cc5000401000d4fc300144000dc44500dcc0d3000000000000c00cc00001055cc0cc0010010c3c0410d4001300c011c4371035f01d00c00c00c1d0c1041cdd031700f170300333f30c03f00f5c047037f34c37f0000c0c4c10c3000cc0dd30c3f0000030043c030001c31c3103000010410c0000141404f010003f340c0c0033c00300ff330303c343030f00c5300101f0300030034c0d30000c0ccd0003c004c70c0cc331c103c113c0730c40103003f0f00c110010d070c00c00c700c3c70000d4000403101031c0343100001c0c30740341000315034d4fccc3041100041001c740103c0000440451d0113000c0f001105000d43100000010c3c00dc0000c1cc03d0013010140cddc00c00007c330c140d1544d00c00000c103471400000c000c0041000441c004300040c104043010c003c1004001300dfc3d001c074d03004413c0310c03c1d0410011c3300403070000c0c30f1d0100100430000000f73c00743c100011530005110101c400030030fc04cc10c403c30c0000c304011c013c0c01403404cf0001104000cc40000c303003d01f04703104000000;
rom_uints[448] = 8192'h100c07003c0014000c0000074300003430c0c04340f0111000400010000cf30c33000034000000c04037003401000c3030400300000cc04f04000030040c0400030ccff4034004000400c007c040000040fc000c3301f0001003001c0000000100003300040004cccc0c0f000f00030c401300170c10000030110c0377440c00c0001c0000000003000000000000044d0000100c00c00100f01cc0013000000cc004cc0000003c1000040000140c00043003cc040000f410030000000cc030007447333004003704040000074c01c0ccc113f300031d010030030c3315030c001304000140040400343000dc000c013c31133d0705040004400000000410000003031000f30047000c0c00400105c4003014f4c0c0000000030c0c4c00040d1100133c00300c000100000c54000030010034003030030000c10001043c0f0f0300343c07000400400400003c3001f00001011c00004000330000041f033043044404c04c0404c00c0100300c10001030000007000030001004500301c00010005c07074050040c0033000004c00053cc0040fc000000000c070000c00003c0000400001100041000040c3000045f00c1004400cc43301030400040c003c001000403040f003000000c77130041140300041040010c03001d0c03000c0300004100f1c0000303000050500300001000f057001cc41004003000100000013450c0030000440000f40404040000130130005c0c3000c000500c0000704744301030040000700004000c0000003000100330005400400041330c04f03000000031430013031030000d0000710001104cfdc0110404000001031410130000000100310004041004004000c00300000c0000504c40033c00001004004000c0c1000c030333004000400d000030c0004043070003040130740c053c00000000443100303030fc000c10000c544c3f0047070c04343c0c10040c0303300030c0c000000c0c040c3000000400100000034040000030000401f030f0000300010c040d0c007c0000001100570c040400304f105400f054c413c00040000040dc501c400000400c0c000c0c30040c0000000000100400410c00cc00070000000000cf34340000c0000000401004c000010440000000341c503f00010c0003030004043143000c0000344c00100004104000000043000c0f13000c140011403c000000440d54000000d0c0000030030004041c000c5000001404051034030d010000000f00000304df1d030000001c103c00003c00003014014000c000000040f000000c00000c03300004030c00000c03000700000c00340030540054000004010000000430440000003000c000000013450c00000000000000007c40340000c070c010c0000007030c0000440000000010440353004304043100010d30f00d00304d000130;
rom_uints[449] = 8192'h5300003004404c00c0004c0070000305c0000003f000000010c33c004443c000cc0c040000000000c3d30703c0003f1300c0c0c3000000c40040100300c0400101c001301040c4c000043013410400c00041000000c3c4c000c37300c0c0c00003410c03300003000c00c000c00cc0c000000c00c4000300017000330000c400c4c1000400000000000000004000100730c0400000040000c0000400003000100110000004c0040300c0030401d00040c3c00000000003000c440303400cc000010000000000c14000400cf010c100070d103100405c00000c000000501003001f40000fc004dc00300040c30cc00700c3434000f01000c000c000330000c500114c400c03f0000cc00300c40000000c000303cc0c00400003c0001400cc3c4000c030001001000000ccf0c0000d000050000f00c0c000c001001003431413000010404010401003c0000cc300041000c0004c00350c0041d4017100c101d00c0100000c400c00100c0400000c4c47c003f300000fd500003041d3400000010000401043043c00001000000300c00030c300cc00000c0000000c000011000000400c3c710c040140004000cc0000034cc000000441c030004004c40040444000014303010c00001000c00003c1100013403010c3000001400000010100c00c0c00000010130000c043c013001010000000030034010300c500c00cc30cc40000001000400cc00040000c00015004101111dcc040000000cc00003004000c7004043010000c0000c00004c704700000c3404c00010c0000000000000014004c03c0000404030300000000c031004400030010300c10013033411004c45000c00000f4010030310010000000dc3444d00300d0d30000c0c00cf1000000430501000410c1c0c10c00d30403010c00104c0f444c0040fc004300000000c4f00050f0ccc34cf000cc03c000000000000300d00c010c0010030cc000013000304000c10110c000000000004c00010000000300040033000000000003040103000300d00000000110c013000000cd0c000000430c05c0300000000c004cc00004c010030cc0001c0d030030110cccc0033c007c0040c00000010400000c05114000cf00041000301000034300010000004c000c001c4003c000000010c000004300300401050040c30140c0000000001740f0410000000010c000c00000000c4000000000c30c13c5d0040000000003000310c0004400000013f000c0c0c0005f004000c0c000000005c00400030c03400f0130c0044c104000400330430007c030000000000031f0400110000003010010030000c0c0400000300000c03004000103c10400400030c04c0c00004040c040000000c000000c400000c1c0c7ccd10000c40100d00c0001003044c0000000010300050000000013c0c0c04001430000000;
rom_uints[450] = 8192'h51c4000003d000f00003c0cc000003010c0000034c4410c00303430133033410401c3000d00000304003407c7c030010c0030070c4140f7300000000c13300c4c0400300c411300010000040c4004c00f003c41c00030700050cc1000404034c00043c004000d03400000cc00000010c0001000040371730000030000cc0400c0c30f0400043004300000133000000f000000000000440c030c444000033d000300c3040c0d00740000c0001414c0c704130000c000307c3000000c05400004030ccc000f0003c30400000d0004000400000405c00410034441100fc0031000003f0000c700304c0000101430011000fc4100000c0c0003010004c00400000c0040dc000314000c01000c1c3d1c000c0400c033040100003f045014010c70cc045f40f00440fc10c00003003c100cc41000330cc00000f004c00c13010000004000001040cc0c0001303c05041c13010c1000330c003c0d003c14c7010000f0044033000d1500300d00000403001cc000050d0000410100f00c07314000300004fd003000c0444c0003340c3000400f14300030000000c0001030010407170030100000fc030000c0001c007015d014004cc0f400030430001cc0c1c40000440034010c301400c470c0570037300000c7c00000304004030003000304d0140df1040003c0500c01031043300000300d000004c0f000074c30c030443013431c14d00c00100c040110cc40cc00411470cc010001003000030000033fc0c0000c004c30f1d4c04000000010030c00c30d0c4f1c10430f34400cf01430c05001000c0340dd000000000003107f30c500000c00301410030400c0011c0c0cc0044300f000000cc00030001000010c30f04c0430441400c4301cc001f0000030c030c010130000033c000d00004001050005003f300043007d07000533000400300001001c003000f0c00071443cccc0104c0440703400040000c40c0c00000011000400030045000003f0000000000cc0041010500000c317334c4004f0f0000300300000031430300000000c300533000004000400c000c030010c00000c00000000041301140000000410040d300c3c0cc04000303540c00000c113c0c30400f0000400040104cc4c0430c0101300f3004141c100130100000c030000d01f4c00c51c0cc0003030407501010cc1c0d40030034c040c041c0300c0410003003044c0000c40f4143000c03000001f010000703d031c10304404d0c000400000400440010710c03004d0030100030010404400000000f0010c4003c100534043f1001054000444c030c0300004c0004010113007000dc000001c30000010000404303000000003f00c000000000c043c1003c010000f0000400000000300c00100000004003c30000003c0031003003503304730000c0100003015000507c4000c003;
rom_uints[451] = 8192'h443400000000000d3000000310000000c40d000004010c030003cf00071c0d40000000040c030000001100043000000d301c033700c01c30000070000c010000010001100300c0041000000100001040c3110050043000300400d40d30c00c0004430001300403000c0c0334300c0003404c00c30000000c000000010030c00171001300000000000014000cc0000003000300000000010001000000000c4c0c1001000000400cc00040c0000000000cc00000000001030c0000004c00000004053000000000c00104c4010c0111c3000010301c00033cc0000000000500000c0000000000c000000004401f000c300001c004000103000004000c004000000000c000000dc000030003000050c00400430d03000c00c4100000003010c0030000041000050100030000030000000d010400300000001000cc040c000f4000000301c0c000c44c00000cc011c000000cf0c00000011f00000000100c00040d04000000c105040f310000c0070300000000730304007100cc0004c100000010100003000400000000011d00000c003c10300003000300100100c011013400000000c0030c00000c10043000030400030001001000410014c0140070000d13010001400001010500000000000041000100c40100000001c7040033000000300003000000c44d000c000c410c400401c0000000000c4301040ccc0004014000003703030030c0c0010c040030010007001004000000f1c00100003c000000000c0003100c333404c70100005f0000101100004400010000010c010010000100040d000fc40035300c0001cf0004000d400004000000000d0c0c1d700510344304340d00c30003000040344400001c0000000d04310000f10000030c40013c000004c11000040000030040c03540000454001f003f30000000000000000000050100307cc00c340c00000003c00000300030000103000c000c0c0300c04000040300c000c00000003000300000000000000400040003000000000400000000300401000004001f00043700000c0c0cc1000c03000013c4cc3400c00000000440300004300001301010c00000010000000007000700c000000100300cc00c10000001001300000000000100030000011040000000000c04030000003000000300400004000404000007000000050000400f0000c00300403000000c30c0000c30000c0000000c00cc0000c0000000000004030000000000004004300000f00034000000000041000000c00000000c0300000000400000c0100000c0340400000d00000401010d030000010000040000000300004000100000030000001c000000300c00000004000c001000000f000101000001000100003000430c000c0171ccccc0000c0003031040000047c001041030040000000100000cc031c0000101000000;
rom_uints[452] = 8192'hc000401140703c30000003000040c040400000041c0c0044c0400cc00010000000cdc0c0000004c000c3300c40130c0000000c00c0f00000c00033010c000034004c000000001c00001c000000000d04400cccc003007c00ccc001030001c3000000c0000c03101401c0040010100040c0403700000300f30c0401700000040c31c0003c0030000000400100040ccd30000000001c403000ccc00004c1000070503c0050f03040000010100c4004044000c000c40c0300000000c3007000c0410000000000c30030407dccc700401c0400030c10700030c0003000cf40c0c00000000030c1000000003cc05040340c0040100c01040000000040340000040cd00000c0047000400c4000010000003005004004f01c0010c000031701300000300000443010cf1440c00000400010f0334001333030000033000013000400010fc04003cc00c0f300000070ccf41005000cf000cc0c4c000030c44040000004000400d30c430004010003cc10400001c0c00100004400c00dc00100000d00030c10000500c400f0040000004c35c03000000c0000c000403d3000c0140000d0401c01000c000001c301c04000000000c000c10157c0101500070100000100c03f000000f0cc3100004100c400c0c134c10030404054c30000400001010030300040f30001400011045000000004700430c0040000000300040d04010005501c000f1c00c03100001000401010ccc001ccc0c440cc0000000000cc4030d0000c70cf10c4c0c0d000040040c50400c00050d00000000000c0d7310150001c45f3c0dc000000000500d34c0440400004000000000cc10000000c30c14c0001c40dc000003c00000c40003044c0001000400004d3d000440c0330c000c0040400d00040c000000c0c0000000c5000300404000000000450c40000c100c430c0c03300004070d0000400cc000400040030400c04000400430033f03c0000c070441000d1000000000000c40440000ff0400000f0000c403040c100c0000000c0010000c0000cc0004000cc000f30c03004000040c0304c43403011000cc01004c0cc0440c0c37000000c010030000c0000004100001000c41100c04000000070344cc40004001403c0c433005000001000d3001c4000300000007000cc10c0300030c0ccc4004000c0001074c0301310f000300000005000300504410000000cc07cc0000c104000303c40c0d0000040400441cc4473f0031400104040040100073340dc000030000000040000c43003144010c1000000700000d003c0413000c0c404cc4000d000cc400000c00000004c00f000cccc000100ccf004000050c40070504101303700d0c0340000c00000400c01c30340c07c4000000cc00445000d0104cd000000c4c040c000000044400000000000000c300110f0041c0000c000;
rom_uints[453] = 8192'h300000c0c0000000001014c040040000c00000300043100140400014c00400007310d040300030340000003c710000c00c04d0c00000000040c004c01c500005001000013030c030000f035000c00000300c0300c000c0033c00d0300040f000c000c30d10100340130c0045030010c41300f030003000004003c440c000c440101400c0f000c000403010100540c000000000000000c000300010004403100030000c3000030000c00000147404f003031cc00004c0030cd0030030000043c4c00040c0000030000000000000d0c001135c10141040400410030011d000c000c0003000c3c000014010300c0005003040c0130c4000000c30000000000040703000303000c000000303001c00330c01003130003c3014301010317030f30400000007031000301040003010c03010cc7000300000700000300f00030000c000c010c01c10c000000000110c00003040403407340004003300000c00c1dc003f0050013030000750750c0c00440c30000c04101030010000c0700000013310300400000404300000300403103c0114000c00100000d310075000c400400c01000000000000c0c00c000c44301050043303c11700003c040030d10000040dc3000000011300000004300044330030007400100000c1440003f01c04304400c0c00010c00010c004d11c00f000c07003003c000000c0c30000034000330410000004c70c00000010103400c3370001101f1c0103ccc0700440c01c100040701c0000d00074000000005dd0341000030000c0000100c1100000000331300003f0001c100c00001030003007000000c04003cc10000000c000cc00101315143040c0c00004d0c00000001000001c00000030c5005c1c04000000103000040050004100100400c043c00c000010003010003334073c040140c0030310c01310100134001377f0c330c004130030d40c0000774110f000100c100010f01000300041000171100000001000100c1043c03000040030000cc1f033c004000c3015000010000c30700000c033340c3050000000300000d00c0000d0540700f00001700c111cf00010c0c0400000537000c30000d700100c0000300000100d00430000341000000070310d0100d000100004100c0cc500700f400000c0000c000c310301f4c00300007000d000d00000c004c0001000110001000400003100c1c100000100d01c340340101c51c000001000c4f0c0c014d010c00c0c3f00000c000c000d03031001000cc030c070003034003003700301440000300c0c044010500000314000000c000403013030c1031c001310001030dcc007100000041000c00300400ddc540004c01c10404030d0004000c30c3f000000301010003301c0001100500000000007d300000500330000d333043003000f4cc004003c1040101010000;
rom_uints[454] = 8192'h4000000c4400003c01c0c1c10400147d000410001c03c04003100000040003010000000c110000c3040001000d1700111c0330344101070d040c0c3d00000c00070c0c0703c0c40c0004f03000c00000000c00330c170c000c00070000400c0c0c000c3c0f0d0310503f03040f030c0000030c0f440000004005c0030504404f3cc0070c07000c00c001c30000301000140c000040f00c4400000f4400c7505000070c000c0401000d0000000001c00050030c004000030000100003001000000c0c01000001000c00000c000c0030033c30030c0c00007540000f30c30000303d400f0c0f10041c040033100f3f000000730000000000304003147c0400c0300c04140000013c0000003c0030104d0000300040013000433c044c0c103f0c0400cc00404c0c330d4c00000c054401000d001104043c04073c300c0c1f031cc0003f110404000c1d0c0c04034000310401001c0005310c00400c430004410d0001040004410000cc000401110c000000004000440400000400701d000c040c0f3c3c1300d11030400000001c45001c3f00440c000c030c000000000d0c304034dcc000c0010000000c0c01c53c000704000010fc0333040c0f030430013f00cd1000303040013c0c010000003041017100010043000d0f0430300c30000d0c3c00000f0cd0c01d0000103c3c3000040000003d03400000100001000c313d000f00000001c15c0030cc0000330d000000100c00003000070c00404c0f000c4c0c0c4000001400030010c0370c0c00000400cc0c0300c0011c001c0c3f004034100430d3400c00010030410c0c0c134c05044d0004000cdc03000001c0c000300003010c0c0f00d003ff0d501000000d0371301d00003404041400000530034c1400c0000c0100dc400d4434cf0cc1033c0cd0000c54cd01004000c00100001c44cc001003d13c0747070c0f0c0c0011511003000433030000400047003c00104c0000000c000100000c0d00010340040034c1d4100000040400303c0000404043000c00103d3c53000014030c000300017403030000440330c0d00c040000003c0000000f44030d000034110014cd000330040c1c00310c00c03c000330010cc430001031fc400c000c000c70000000000c330c3c0c03070c0133000400c0c0471c0000103004000300100ccc03000c0040003000c400c4005003303c4047cc04000004030000300004000d00004f001c0400010404c130f404000434733c43303000003c0004100f0c10000c0041000100000c10000000c03c00010c00000040cd40501c00003c01400d73c000c000000d030130000000000c10000c3030701304c00cc100413c000c0401000300000c0c000700440010c444100c000304074000040440c00d401c070000003c044100c0c00700300f04003c10c003100400;
rom_uints[455] = 8192'h140000000040030000001000001c010030000000300c000001130c0c0040000c003c1c0fc000000c00103c13c304033434c4d5000330103001010f004000400f04041300010c00dc10014c33400c00000010043303043100040c1001000300000cc003f104000c300f00301d0400040000100f030000003004300334100000007d0d1111040000c0040000100c0d1c000c0c103000c00010c5730000070100100530000301300c040300100f03003033000c1400030001000c0c040137000c300cc300000c0007300304000000000100030c00000d037100000c0c0014000000000000770c0c000005100f3404f003003404dd00011000410034300cc140000c30703017f030c004c3040305501004030ff30000110d330004c004f04007040144d4100103c00c7000000000000c3c04003c000010000400000700003100130c0300033000000033070407c000101030c0300c0dc4130007000f1370340c00103fd01dc500300044010000000041040c17033c00010c5c00003f3000040d1000000d0005030f00000c00001000000313000000000000000c0113101041c00c004001000c03cc07d301330c300c015304000dcc00331000011c0000003f011f0c073303c00cc0c003040300003c00700c0100030c0c1130c00030030c3c00300030040301013010d0004c040430330f3400033c30433030f3300d0001f1110131000001400c0f01100d00300001030311100f3107300c00103300040d033c3010c307d1000004010c001c100000003003010400040c0007000114c300000c00000c11c00000030c001010010cc40003300000330c011034000c00dc0dc40c0c1005d0000c03000000300007c3c05c00000c00cc010c041c03103c00000cc040c1000fd00000000c00300004111d0433003044040300304c30030c00c404000037700000000030041111101013d135103d3d150c000003c3003303343001041304300100000000330033030c110003000300100403000004c40000000000300004d0000d0f300304000003040433d005d030100307300500000003303110400001fc000104ff04001300000400003300c3c100004400007c4030000d1c0700c301c30001000001000c00d00100003004040001530430c40030c40000010d3400040c0c00c00030000030000003c00000003f00040001d00f103f000c000000cc3c0005073403000c13100d01031c44100400001110010fc1050c1000d005001c040c35103c000370f300000f040000c00c0c005003040f00000d50010053300c0013033003010000300430001c00010c300000003010050400000510001c01330001004030300f0c140001f00004030c0100031030010000003033000033300c01000000003f00000010000d40000030034000040030003c003c0113400000000;
rom_uints[456] = 8192'h304100030300100000007000007000100000100300d00003100000010031033c0000000c00130000fd0000000c0340000000101000000000400003000030110000c1030d5000000013003fc10c0033303030400003c10c100000103040004310073010c000c01033c000100c010010000040c00030073003105010000433d0000030001500c03000030010300343040000000004003750000c101000c000c100000003010400150330000034003300300000001030143030030000003c031000001000400300001700004c000000315004c04373043c0004c300000010000040014c351000cc000031cc34500010001000000040000000443000000030000010000c5100d00000040c30003340d0300314007040000100cd00130c13001111003033c00c000010000304100000000000000000001000040000c00d000003010000403100010070d303000fc0000c3df0030500000000000f003cc00004030cc01300000000103c000004130101300c3c00000f00103f04000000310040400c00000c0000040004000000010030001304004014733001100403000000100c0011300c00010030004700010101c000c0000400300c0d00c0040033303404000010d0f000c0000300000c000000440000103c03c030000c00000111c0003700000f0003000000f0f004100330004130300000330014700000c33033000cc30013001433170000000c00001c3100d4100000030cd000000000000040d000cc001001040400100000140c04040303000c11040400003400001030c00000000000005030000000014dc00000c13040000000003030000c13040003301030f0140100007444400030000c1000000004004440d0104043000010003301010c000400144004001303040003030000400004334100300c003000300000c000100000031001000c00c0c0707c0c10f00000740c10000000005403034c70004c000c0000000c0000000040000007c400343000310f000000400003000031713c0010100000400030c3313041100010300000001013000010000003000c000d0113000c100070300d0c00000000100000000d0c000030100030010fc5300000003030d140000030c003500000000030000000000104100000003c3c03000d00001310005c000005300c4010400c0001000c0000100c4500000010013010100c000001100001103100101010001010c00000000c10513c4400000100010000003000003c03311000003100000010fc000004414033153700100c010000300030000040000033000300c0730040100000300003003300000000330300000000000130300003143000400c01300c103dd010000c343011000033300300004030000011d1010010000331331000000430c0004000f0000000103000f03c41010100000030;
rom_uints[457] = 8192'h303000000000c004000000004c00130410030000df000f03003000003013300400f00330c30300000001000000103030003000c4000f03000404f00000c0410400000000003100f0000034004df0f0003500011000301c040c0300001003000c03330000000000400000d700004d00403c0000000c31040100510010401300004dc3c0000503000c000003c000000004c40000000000c0001c000000043d1dc000000400014000cc000c10000000300c0004d00000c0035100000011cc00000003c00000000000000c04000000111100100f001003144ccc00c000d0c07d103000300000030c100000304050010330cc040030100004000100000010004000150c000010103000000030c00041000cd44034000010700000c0410030410d004000000c00c300004000003000c400310003000c31000000000c34001000130000c030003000cc0000000314f4cf000000410300c0000014c4c0000c00c311410300003134c43c000300c4004000100c00004c03000334001403300000400001c0cc0000d3c1000000031c0000000041100700000c0000001000c101300c00000041f004000000001c00000013c00001000001040131000004c4004000000c7d000c414000003000303003c0101000400d01c1000003c0003000001040c00010000330404404c00007c4433070030000301c3c00040100c0100010030015c00530000400c000000cc00031001000c700c030c41000030041003003370030000100001c00053014300400c000001010100400c510000000300c10030c0c0000c000000034000000000400053000000001000c000c000031001011000000c4400d00040000000003030404040000c000000070030030d0000003000010003000c00004300000000041030001003040000cc013114c14000c0441000400034000001c004700000000c307c00000030c01005000000000000030010000330001000000000c003000000000c310030304d310c030c01000100140c040050000c00c0400c3000400400c00000000040000000030000003300000100000000f40c440000000000000301030d10c000400000713c000000000010c001003300400c070000330100030ccc0000003000000c0000c000010c000131c340030100003c4041000340005c000000000000000300c0110001300000004300000300fc00000040310000030500c500c33cc00c4000010c00000f3d3000004133440070000000303c04010c0003c00000304100000100303000004c0303001f0001fc1130000371004000c030300003000c00000c40c0070f00003100100000400000001000000c3000000010000000004000170000054000cc40000400000001f00000000fc0000c40000340030000000003410110000c7000c00303400300000030c0000c0000000;
rom_uints[458] = 8192'h310010100c300003031040000000030304000000f10c00000000000c4100000300070cc0000030c0100c4003c0c413500000400070001c051c031c00c1003000010310034007130000305100030400741c00170d00300000011300cd0f4030100000030110111141031040003301000410003040000004000070040001030303071000c000000c01030005000000040c010300300400f00d033000000000000041341030000010c00000f100103300c00c0100010300000000040000034000c00c00000003f1133003100001530000031730003000300000003030010003301c104c0010030000110c7100f50003000150353c00000300c30300c30130303c310000310333000000000001040010030000c00000000000000107301c030c5010000004037004000000140f000310333000300003000010c014030030010040f00110301300001004300c30040304311c40000057305003005c311c30c0000000c03411c300300000101000010c030010000340301100031c10000000c00c03041f3370030030c070030000030c1010040400100034300000051c3030430001dc00001000003030400c00000001030000030400310300770040303c00703000001000013700340ccc03033fc0000450001003000c443040300030001f0d000c03000000030cc000c130400cf0c000130000304c10000000305030400001c00303031004000000000f003c0440000004000000f040f100311003100001000001501400f010043c0000400131300000d0c031000000000f000103300030104300005000c00c00000700005c00000000000000003000000005f03000c300100000000000001300100c4000301004340c00033c000103300100030030043000100034f0003000000373100310050011040100000003000140000c30301c13100cc00d0100000003030300130f0000073303c4000010304103000033003053c0d30000300000000103030c003c000f30000030000000001013750000000fd000c3340010003030f0000c0010000300030c000010c00010000010040c0003343300300100303000001001100000000100101f300c1371100040cc10003401400010700000700303101000f130430030100000001433101000000000c0c0030000010300c3001001000c0303000000c00c00300c11303000001c03330000000003330100353000040003330000500000000300030303000033000f0010330d0004100000103303001c0c3000000000330050d0041004100c13130d010000030c0030000c3000c314033070000330400110030010030001000c0300400000030013130000004c003cc1000300100000010000001300000010301300000000305d001307400013c034334cc401c0000400300730000040401000001010040000100030;
rom_uints[459] = 8192'h400fc0000f0700000004c000010c0000000044c0000c0d03704000305c001000c01c010c1c4c00003c0cc000300c0004c1341000003f4130004000000300c000000c0010004000cf3000000130c1000c43f4001c3c100044000c101040d40003c000f450001403000c40010030300c053340f3000301000c00470000003fc0300000000000000000000000040000c03c003007010f3f0100000010c400004350c13003c000300000c0000c140000000c000004000c0c000000100000c0000000c0000104c0030c0c00c00031f104c00004d43400010c000000c000000030c0c0000053003c0003000130c0110000000000000000410cc00007c0c03001c70031c0103c03c00c0c100430113040001ccc00c0400301400030100400f0000404400c000000104000010f40010000404100000000000004c00100000cc3c01ccc0c00400000004c40030043000000c4440007000c0fc400001c01c4d40054f4040c4373c01c00c407035040403c40f0500401004c0400000001304c0c0401c401011010303000c040030300000000000000040c05c044cc040c0400030c44030033000000000004c0000d0300134c00c0000f400043c0c070040c004c010040050c04c0300100100003c003f00c400000330001000d000400c740000c400c33530003004053303003000340cc70100000000030400004400314403c500f343040c0000c100000c0040000341103030400001003001300c00004c00cc100004001000000073030000000c300403000004c403010d40000000000004000040010000c00004f0000403100c1300000304cd000004000001000411413c4c00034033004000c0c0004010040000004104c000c03004c410004c0400000040c40000c00000000f0040c3400c0c17030f1040c04030000c030004003c0c040730440000000c004c0c1000114005c040455c000c0004c0d304000c00000000003010000000000300000c00000040000150000004300c0c0000c000c1041000000401c00000001000c0000300004d040044030000300003003030c004010004c0000000440c0c04c0005330300f4004c000000054004c01003101000310c00cc7f00003c04000000c3073000000000000c11404c3000c0100000c0105c003001c04c0040001000000000000030c4030000000c000040300740c1001c1c0000c0100000000100000c0cd0140d0000000000c30300030c0110030000c33000005000010000004d01000400c000c035044014f40030313000f000c0004c37000c10005c01000cc0004400000cc30000000c030c00000000500030c30000010401400c0040c00cfc000003c103040f00d0040014000f000000001070c10034000041000000004f0000c0400000140000004c00000c0000000f0d30101000000000;
rom_uints[460] = 8192'h430000000014d0c001c0300100c000c30000030c001c00040307000c000000c111100000010000013000404000400c00c0d3000301000040000040000c00101c0000000000000c030300430c0c0cc01010100d00c000c00000030000004000017004c033000c114070030c00307000000000030c00c0340cc0d1444000c00c0001000004014c00004000004000050000000004000f0000000000c4433c40040000c043000000000c0000400ccc03c0c00000004c010000003410001c0c5400000400c00f000003000010100300000100400f03410070000f00fc004400010030f4030000004000cf4010c4047003340001c0000030c10000000340cc0300c0001c00000003c3000730413c007f4433c0300000c007c00040cf04f33000130300034f00cfc10000500100c0730100000000003c0040000c4000000003000343100010000040440414170004c00404004340d000010400d0c000401000005003403004d000040301110743000070cfcc00040040000dc1130700003c0000c050c0000000c0004f0000f3001cc44010403c0c00c04c00140000040d0001c000c0c0cf0000f34304400030440304c30d0433430fc30c01c001040c0c07c000000003140340430000c000000c0033c0dc4f0400400c003003000100370000000000000100000030434030c40ccc00d00000c10000030000003c003c0001c40400f00f05100003054c0000c01100004010003100c00400c10000c100c00000330040013c01000000000c00dc0f1000c0000c3000000000005107c000000040300f11c400003000003c03010001300000300500003000c0cc40000304c00141000500c0c00100000300004000001000000000430c40400004400c000c1000101004000c43100cc30101c313030010050fc0000f100000000c330000100000400c0030100310044040470100140400107040104c00c04c4c3000040c000110c04103fc030400000300c000004c00000f431004010431f0070300000000c0010004001301c000000000c01014004000010300010300c1c0001003030c000003c000000c3c010104f10700400c000400c100c3000000003c0040134700dc004701c0cc0000030000434003000003000000000004100330000fc00400040100000cc003c000400000030305404c3003c0030000d0c040f0000c1c7300000444d400c00100000c040004000300010300041000000030014043c1000000c000000300000001000400d0437401030000040401410c005c00014300c0c30c000300000031000305000c047000d3070004300130000000c00300100000cc10004000000300400040003401010cc0c000103000000100000cc003000000c10c47303010c033300c0003c0001f040003030f04cc030fc00000000500c0040c000cc0000030;
rom_uints[461] = 8192'h13c00000000003000f10000070040004c000c0700100c001043003330170c000000304530f1c300030c10413000330000000001d10001030040100313300000103c1c0003cc0301000000dc1c000c1034031d01c400300c03400c03c00c4c0d030143370c01100d07c3400040300003000100000f31000301114103001100100f00000400000000003300404000100141c00000000dd01030d000304cc3003150130503000c0017300f4000330dc0004001030c000330c0c03000001d0003000c13003400000010010011d40000331001c0c0004000c74031c100431310011d404100000f031500c100030034fc00000003c0300340000300004c00000c00001000300400310504130cc0100000004c0000100f1310000010c00cdc10c434040040000000411d00000000003c0040040fc030030530030c00001c003000100003010310000100000310005f03fd00000004001130044003c000430300010043103000000c04370f1157c53541cc000300f010010010c353000103c0c00011004c0354001300001010034000100040033000001303004500d407c3030040104100441003d000400330300000c3300311d00000030043000000113c1000040304c300000001000c4c0010704000000000404f13300010307001f31401000013701d003ccd000d010000f00400000d330030c00340040c007c070c0000cc0007c0130003c35010030000100000d44d011d4c01d0000300d0030300310010300040003c000030fc00c003c0130041401010c40010000010300c111c1003000011010303c0073000d30010100100040071300010400011003c000300010100c0317104d00100100c0051c301331040c40000001cc01000000c34310140000000103000000c11017000c3400031f0001300030f07c000300300f10c0407405030404c003c3003001303ccc001017144100c4000500310000c0010030070c1003001070d03c711010030000313033310c003000014031c340403d00d43001cc70dc1400100030010000030d3101fc10c0513000143100003c00000f000cf40710043003c03c1110100c1000c000010130000435dd0000311300f01001330044c00c040340000c310000c0030f030000000011001030c0000400c01040010000300430c103300040c40c300000000001000000c4010101003f4001c0330c000300d10100101cd01011000f304100011300030003c01c3000000f300333000030c1c1c0014037100010003003000c0c0735d117c040500c1005003003700000c51000341710000003000001c00101001100301c4004f000100000000d00300003104f004003050400c00f4000030c0000c0000000c330300001c000000000000010f1003c00310000000031cf0133300404000410c00100c00104000030c1014c000c400;
rom_uints[462] = 8192'hd0400303000000300c000000c30400314c0000403300c000004404040030440c0100035d0000000030400c00000400c30c104000000cc404040000040000c700000c000c04c00000000040400300c00001c00010000c300001005d03004040000010040c0300000001044c400400003fc0c0007400000301c140113014c004c003015c000303000000030000000005000010000c00040000044000304410300d00000c00005001400033040000003cf000041300000000030000000c00040003003004000000004010400003c000033c3d00000304100030003000030030c0410040000000440000001100c30030000500000003000100000001004000000000070000003c400110c0c000001001000000c0000000304004c000003400c30c0400400000c0c400000000c40c0000040c4033000300400300c04003c0000000030cc1000000001c00500000f0430d00000004040d70000000c4044f440301410107c00400f0004f0000c30d100307031c100007c0010014040001400000000dc4000f004403d0040000030000040000cc00000000030000000c0004130000000404404010000001000001000000301f00000000cc0c000000c0000004030f13050c0300f0300000c0c000400cc1c04030010000000100400c00000c0100000040c0100c41003d00c31400dd0003010300403000014000010000004000c0000000034070c0340f04000d40400050004004040003000400f00004004c0004004000000415000000000000001000000cc00c000c300300030c30000004030400c00000c300004d000c000140000003cfc00040c1000034004003f40070000c00cc0530040000040000000000030404010000c41dc0c0c00004000cf001300000004000c01000000000001d00000003000c00cf0cfc000f30001000c1040053400303440c030c0000cc0000313c0c0c13014d1000400000cc03c0000100010000300c0d4040c40000010004430000000c400000004c000000440c044cc4000c7045100c0040440400c05000304410030f0000040400c3400000000c0000400c000700010c00000000c100070004c000f4035030500cc0c0014000040c0c1c00000000400000000c0000000313000000c00000000000000c00010ccd040000101c030034c0000400000000070c400000fc14000010000000000010303c300000c40100000110500004040403000100034051000000000004010c410c00000000050400000000c403000100c103000000340400340010c3c3041f0000000000dc040401043cf0c74000000c00000000000013cc004c000c11000000000000000d300c0004cc14404000000104400c4cc404000d000000040004000100c0001c013000400004000040000004100000000100010104000000000030000000007400000000;
rom_uints[463] = 8192'hc303c0c00700030330c00003d003d0430fc0cc0c0047c030000000c0040000003150000d0100000000c0030f33004100c01c010373c30c300001030300030cc101010c00010d0041000440f70000710c4303040c53c04003304303c001000000c0331000f04310000030000000c0f001400f1101d0130004030001cc03100000cc00c04001000011030000c4c000030301c000c00001030000000100400000c001400f000044c7010000cf00c0010041300300000000300000000041434003010030000c0000000c00c000000003017041030010c031c00044010140003000010340100300030000004000c00cc00100c000c370f0400000031003c0040000443103000040410340100340d3400003d301c00000140000430300cc10cfc00f4400cc0001c0c030d04043c0000300004000c0c0004c010001004503cc100100005040c4100c00030f13f0c1c0c0004000c000c1dcc04034c1000cc7400001030003c000c0000304004000041004c30004030340301000c001000010d300014000d001100100c004cc0000000470070303400001c0400001400010c300004003070d103010004140c00100c30000040100334c03f141410010500300010400c13cf411004300000033004000c13003c00150010000f0c000c0c000300104004010010c004174f0000c01000003000000c01000007000f1030f0d740140c4c043d10100400003011000400333c0c143034403130040f0044043c303400000cc000040d30371cf0040000100404c007503730307c00c003100000401c00000051000000f00400003ccc0300000d100c000c000357001400c4004440300cc00c3cd410c40403c00000300c000cd1c00c04301030c00cc0000c0c0c410c3c410400c0014c03401000000301fd303000003004c044403004003000000010000300100c10f03cc100c41c00003c140c000314004c00f03c000c3c000c003c0000050c0c0000031000000010000400000000004000003cf00030041f00001c300c040000c000300070100c00003c0d00400c0004000000300000040cfc130c003c1c0c000cc0f00010001034700000c000040000c3100c300010000c004014005d0400d0001100000cd0303004300434000010300030704c0c010400d40c0c40003ccc000030000430100c000010d00c4c0010000040001000040cf450000100c03c0c1000c00c00000c003003440c343d00c0c00c000c043030341450500cd0000300c00430010d1c0000030c04000c300001043c33000c5c01000034040440401f0c00c0040004c00c1403300010000000040c00030100140000000004040000103000000c440d040c3df03004d400c0300014000000000c0000030c000104d00100003003440c111410300c04044010c00c00140000300000000010311100103cc400;
rom_uints[464] = 8192'h400f00c04440001c011100003003040101000010030f000001040300300f30000c11003311050c04040100c00f0c0f3440043f0430430105350001000dcc000c000000100000040f000003340000f0ccc00000c000000f3400043330004c10000430100f0033000040000000c3000c403100043f000c03fc00310110010d00010c30c00000040000000f300c030004000075000400400c01003c000001100104c40c070000300c00003f0000c000d70300040f0000110004400c000403130000001433000000114c0fc140c30c000c300401074c000004000400030c000404010301000c030001000003033400030000004003300c050c0000014c0cc10000050400001003cf31000c000051f000c10100cc003c400f43303c070054000f334704000000000030cc00010c040c0c00434c40c33004040d00000040004400110c0c000304040100004c005c14c34c0044000c01000f0005030100c73300000104000d00040c0047000f10070c010f000000000130c50c0010c0300f030c4100c4030c1050400000c1400f000c7000000c3401f10c00005000010101030f013101c15f0000000c00000c3003400303f701000400f03d1f0c00c1000013110030433d0c1f00000104000c3013000100340041030c1305f0f31f00000000c304300d04000c3100cc04000031010c3c10001011040400000004350f00301000050433070030000dcc0003003430040430353105c1c1011c0100c00c073535004003c0f4400003c3050010000007133000c03000040c030014c43001400004030001003330350d1000000000c0040c001c3005010c000c00000010c00c3c00104400c40c04000000000c0f3301003000000cc01400013000c0010cc30d040c3300c10403030301000000003d013100000301003c000410303003c00001000030000000003c000000000710050300000433300170c70403554c0c0000000c010c004000cc0c0000000000003000000700000c0033100031f433000c07000000000f00010400030001011d00000c00034c1c03c0300140000010041300010000053433003003003101c0003033000001001000ccf404000c010c0d01000d10c31f030007f13001c0000034000cf00f0100000310000000130000000134010000054000341003010003033f00743030000f04c4000040340000100c0c00f353000f0713000001001010340005c0000000000004373004000040f0030c0100001440000300000c400300000000040400000f003d070000000c0011000043000cc0301300000103410400003031004000310400330000c40c0107000c0c40000000010740000c0c003100000c0003031d310517000300c40f040004040141143c070d310040050001000000000d33100c0304331000040100000341040c3030400344000c00;
rom_uints[465] = 8192'hf34300000003300003c00f30c3000000c0010cc10c000c0000041140030d0300030031d0030c003031f0000cc10400f10030400100c0030d040100c0c100700000001307003000000c00110040000000c0001001c10c110000000400c0410003305d0000300300000000d04000c00300300c00440040030300c03443c0034000cf0c0001040000100501c0000000000335c440c000000103400300013000c4000040000300c0011103c300014000000103030c4300000000000003315300c0304007303001000040030400001053fd3300c01c1400000433310101510033000344000003c003100030400030034c0300004000f0400700100007040300030000314c01004030040000003310c10004003dc000f3000040044fd030010300c0000000c000c30cc0000004c003c000c1000701003310c000000300030c0c10100011014c0001040300000303100d010001000c31030c1104c004c0405100d300000030000070015c31000dd01001404010030c01c30044030304004040010003013f0300c4031d0300015001340c03c300c100300000001400c70331000400c104040c01cd0c3c030000000c0000003100331000f004400001004000000101cc100001c0000330c003001400000f00d00d40000300c3000003010c000300c045c0000000c30403c403000400c004030001c100cc11010304c4103000003030000f030101100403033f030000c00304c50c000403040000000007c0c0d4404050000d4c100000d0130100c100010040013300c34303030100030700c0c01000003007301001030301030007000000030000003004000433c00d0043000000000f03001100000f0300c3010303000000130300c003040c7103c000040c30410001030c000000030005d304000040c30001000011cd30f00000c0000c0300c0003003c3cc000c00000030070c43c70300c4c700001300113c000310000310010000cc03001003000000c000030000000000c000150101103301c0303701033c01030440000004330443c730000300070c00310101000d0fc0c1000003300401c01c10c04003000400000c31001100030f00003300100400030043c0003f0f404c010005000030f1d1030c003101c40040000040000310003d00001c00134015000500000c14000f000c01c3000300c03f0100000000000100070f400c00000000f0d4000003070d4000cc4343000000000f1300c30d07c0003d00010103004710c30001000c010f00000c05040c004003040004070003010010004d404c0004cc400004100d00c4400003c30000000000000000c10c040100000000003000c001101c00c030c5c1034c0000000104c0030000000000c1030000000005000d03044100c01000c0c430030140304000070c03000000000c00000001dd0c000100000000;
rom_uints[466] = 8192'h1c400100c30010d1000000c1f04000d443c00010000f0000001010403f400100311040301000710100000000c03000003330000007c030103c0000040011430d30000500000c0c00000000054010c04c005cc301d00010004100704301004c0030f140103000403000c11000310001101c000500103040000004103010d000c170f340c310f003000400000f400000000000040000000000f030f00001131000000000100041000100300000c3330400000000000300004313400000001011000c000000003c04000104015403010000c351040033103d003000001001d00000000000c0400030050c4000c1437c0040000330c033000000000000c0000300c070030015c0c400004000000000701c310c430011000034cc0100c310400001c500d0000300c000305c40000050dcf014040000c034001003000010f00010000040c0c0c030f3c0040300c3017001000000000000110300435cc0c4004c00041000fc000341311001005000303440015000000c0c005000003f450000010c00c0005004c01000003010100000330d0304300c30000104d0c001000430c13c00000010505000001000003400003040000c0001f00000101c3010010000500c4030c0010010f03000404000000c1014000431d05033001400c0000c10c103400300070333410030d00003004000c3540c004c303104000004000cf1301001c0030c4c4003cc000300707000001cdc10300f0030043000300c103303c03d400341cc03c000703f4343000410c0030014c000001100000044300c103301c150040d100000330030030000c01300004014c0f033010031003000005c3000100000c03c5000c0010000070300010c40c0c00000130000100100f000f005c0010c0034c00c00000410c0005c33c000101101c0004d13131d03f0000003f13000c00000f3d30000100140c303003110c040000741f01000f0000004301003c33031000000314101030003f00c40000040400030000100043df1f0100f3003f00003004000500001cc30c000010030100014400434000d03100300100000000000000030030100d4000010000c4000011000000110001000410004000000000011c0c33d1000000003110350004400003000c001004003504000300001000c03003100501000c03000000c4000070000010330000040400100710000111c034000cc00c043cfc4000001f0005000030c431000000000030000c30000410700000330040d010000103100010004f40400100030011c40040000001c00033300030100c00104004c0015000f000000000030f0000033013100400040000000c00000000000000070570004033c400004000100000000300000c00300001000c41000034c5013130040c0400400300000400f04400000c4d000400301cc00c0035433c100000;
rom_uints[467] = 8192'h43000001010100d4cc0000010004001300d01003000700004f1300040cc100010c300000c300300001c0c03c00c01c0c0574400003031c41c001d3040030003103c040c14000303000100cc04005c000c101007c4300004000d3ccc040100000d147100400040c414f130003cf3040f00033450c30c10000530004d1c100000fc43040000000000cc10301cc044d000001001000000c1104007040ffc00d0f41c010000010c0d1010414000073014041000303000004001300000003400440000c303000004400c30104000000cf0043f0010000537010043fc400333c00c100c000403030cc043110000033341741000410cc1001000000000100f4000000035000010000710000c000c010c100010cf404c114143374d0130047043407130cd0000001f00c0050050103d301c30cd1c1400000300000050070001fc111c00c33033500004000d4030407000000000430003400340000c33447514400001013304007cf300440c003000430403c0030cc0c00001100705300000000004403c0cc0c03d3100301130040410c0130c07300c13d0004000031050100000140c00d40301341000c470000c0000103303001030103fc000341540cc0d40c00cf011c0ccd000400c0c0c4c004000100004054000143003c00000003100410300031003314050500c10034c110001d070000df303040003301c001c0c1000030100003034000040004cc01d0c00030d0cc14c0044100000c000000000101c1330f0140c41413300d47000003001007030c043000000303034104c0000704101000010011c05000400000040447004371c00034f144304c000040000101000c31300f0010010400f400c1300030003700c00c04300110003c00c10c100dc0000000400c00c300c704d01c340030c13c030044c00d31030045030c004040c434000333040031c301c10330f0f331f10000110c701c1040403000c071407714405001310c4000000400000030043310030044003401070000000100051443044003f104f00000107333c0010001c500c00c100c0000341c770d00000000f400cccc370303004010010404d1f01010c1010300003100001d01040000d110071c4000f000013100400000000113100341041440040003cc00007000101141c5400000c4004000100dc04000400700c000000c1040004101005040000000f04001f0c500000100c304034d003577c403110000c040c0147001010c43001001014c000007000300014000004d00c44004003cc3350001cc3031301001000f0300010144001017d0c334030c4000c00000f070cc0070014330000700c0d01050000004310cf000c0c4f000d131133cd0400c30d40301004044404003000c005001cc114041000300c40001300000000340ccc000000473501000000d0c0041001740000d0000;
rom_uints[468] = 8192'h10003c0df00c0000cc0c303100fc40f00cc0037001510000f00000c500404003c30343d0cc300000500004c0100110f1000f4010300440300001070001000034330030c00f0c5000010c010304430f444c000440000040400f33000003c30dc4c0000043004c0c00f0c07001cc4004000040031040430001f01f40f1c340010f400000035003004030400000400c3035000000000050c051c01000c3cc03173143cc1000040003c0c0003cd05000403c03c10003c040011000000450c0400440f300700004010040f05000c053033c000040c00d0003334f430303f1c000030cc030730300d00430000df0cc3007c04143000c0c000000c0440000c10000f0010d0c50104410c0101f40c030701fc1000000f01430c0c015403401cc00c10003d0000740000d000000c00300000007c430000350c0000000000000c000c01000400030404c40003110001040073070c4c30000f040c3301c5c0170c005c00440c400030170c300030040400c0c305041030c04c001000400000c00000f10030cc0001cf0cc10c00100400c400cfcc1430030404000430000700301000043cdc340cc0034c01310004040c00c500110030000c1c400c133c00000c000007000c50430d30010000300c0000000000c4443300000330c03c30100000c300c4100c00c110000c000cc1473c10cfd10400010040000c1c0000cc01c04130330030c00c0f0430fc000c07030c3c00c00005c0303100c4000074c00000000303fc001c0c0000540004003000c400000030000cc0c304000344033c0450001f0030000f3104c03400043c0d0c000f4c00f4000d054c34010304000034000c341110070035000c0c000041000100011c0001c015000c70c037c03f0c4c0030000000000000000500000003c00c0c30d00100000c3300c510c0d0074005c00c1f0700300307030104f43034340534700d047c0c17f00f34000700cc0d0f0dc100100300c0001004000000fc0303000400c00c3100310f0c000c0dcc010c40c00030400434000030d00c000000310c40004c0f000c3c370c0403040003c00cc03500043c0d07000c300f05304500440c00c1000cf000053003c0000c00f0003f33003000040c040001040c0c0000470000110000040430c0000f44c004000d00400c0c1c01c5013500110c3010f14340710ccc030c730f000410034303300400040c3001c5040c110400000440301030700003003cc30503007443304404003410030f004f04300003000700101070c34400400f1400c111070c340003c4310c701001000034007030c0000c300c0004300000170003040330000c0c03004300f00000cd0c34c00c000f0f0004001c00301000000300001c0c040431cc4300040100033c001c05cc300110030050f0341300c100010c0c30c004300000000c0700000403;
rom_uints[469] = 8192'h400c0004000100fc0040cc300330003c103340c0105c400340c400c0000100004014cd0017004000104000c0c0000353c010040033500014001100000c004103000010d300000470400071c0c10004000401044013c0000000c0010c00d11303000cc01013f001101c07440050400300037000c41051003c000d001cd400c0101040000040000000c0d00010d000c3cc5000010000000030ccc10cc05034f00000000000004f0c0cc010040400c10030000000010000400d000340004dd0000000f000d00000c0c1c0004050000014404c04300c1041c414004010d03404300000c0c030f3c00000000000c10043001c00013f0000304000c00c00c0000104c000013030443000c013c10c14410004ccc01300c4044111003004010c4000030000d0030000d0000d0000404013030010c0c000c00c34030000000410414f14004c00014c00c303c010000140c000c300141400100c14c0000000c0041000340040d4d01041d400cc00013c7c00dd014000301c00000c414000ff50c10c0044001ccc4310045400001410c01050300030030010030000001030000300c1404c00055304d04000d040d03c10c0303001003000cc4000c043c00400c00c44100030040c0000f00300000c030000030000f000440000fc0000000c30400000100003c000403304000400d403cc0303040000d7c000033004c00c0400000c1000047c4c04130d00c0000cf000c00030cc030010ccc00040c000300000f0c04000140400000300143c4010004010c0d11004c0c0c1c000400300c0040050c4f000d1004c00cc3c00004c00000410d004400c00c000000c05000000c0030c00000474c000301400000000400000c14c1001c00c44334001d00040d0134110000d00c000143050001000cc4300d5330040400100c01070000000c077100f0000d0130c100cc000130117c00c000c10cf004344c45000c00000404004400003300c00004c00c003000000c0000c0010c000c0400000c0d404f0c000333c00000c40c0c0c00c00034450003030040c0330400000050444d04010300f00000013043c03050000004f403004300501000c10001c0000030c3c0040030001c00004c001004014f001004000c001001c00000000001000000001110010c00040310440c100c30030ccc0c303134000430c10004c41c7101c0300f04000cc3017c50c00000003133430300040c400f300c000440010d0000000000100c010f05054005034400100000c430000003000cc0130040000d0000c0011430000c00010011c04004000d04010000034740040000000ccc000444c0013004c0000100c0030000030007000403cc001000c0000100c040003100030000000c4000c0043433000004c0000300400c000c00f00c005c0d011044400030400000010c013c00300454040000000;
rom_uints[470] = 8192'h110000400f400010300001101001c0431000100003f0300c011f0d4c114043053030c0001040043030701f0304c3300000c0010371d0000030c0300001003000011000004030400000003540cd31c0000010100300133000353030c003f3c000001f03000c004001c0c0040300f004053500c3d4000030000000f00000c00003f03010004000700040330070010000300100100003f000c0c000003140001010404c3004f003f10130100c43130c500c001040000c30501300053310c0f0004300c300000000030013300004104100000000700000040000004303400000c000101c1f03000f0044d00000003000f030701540001000000c000030c03003010140000103033000030011c531030010304041c107430300154100030010100500d100000030300500c01030c0003100700000c0cf00d001030100f00cc1101c03717030c31c1400c00003cc004403004000301035000330f34043c000000030c30033007050c10540c00140004170c00303000000c040001300c0004014c00300000f40300103000030000500003030100000f0400000c01001010045300005301330000000000c70c00050033173300004344300300000c117005040103000037440010000000001f3c3003001031140c04000304d3400cc0000d0c0700cc013030fc5034301300dc001000c000003103c303350030000073000c0000500104300d03001000140003000040fc010030314043f40c00000400010104330f0004404403c70c31000013c000003330c4000c0703113010000014300000000030000400c004000000010000500010011c00340c0003400000131303003f030001f00010040030000100000010cc070c00030100140000d107100704003000000d50043f00133030c3001130000c37000013730c00314c5017003100031f1003000c13000f300434300f000c3f3c30001740001d00000003100100c700005101400010005004000c00ff0dc00700c0010000043005005000330040003000000000c3000400300003010000000cf4130c001c10f003000030000c300c0100071000c01c01100cc30043f53000000000000130000030140000030c00000300000010c40000000500000104030000040c000033003003043c00030c00000303300f0c10c334404c000c0033003f00c4030031000100000031010000c004000304300f0c0110014c0400c0330433040400030031300307500004503500000c100d104c0500110000000c0030000000030107403c00043c0400c0000500000003c00cc01000000003030ff110040001040010000005000504004330000010000300300c0300000c0400c033370c0100c0040030430d00030c00003c0101c004000c10000000040003000001040001070c1501300000000403010c07131150030c0400d0;
rom_uints[471] = 8192'hcc000040f00100004000c000000001001d000c0000c40440000100101d304007000403000040000c07000000700000c0000c00c0001c000100000000110000001004c0030000000000000c010000c0000000403004c0c400400340c000d0c000004300000cc0000c413001004000044000c300c004300004004dc00400000400c10cc00000c000c4031000000100000c0100000000000000c04ccc000000000000c00000300000000004000c0000c00400030000000d000101104004c001c0003040000004000000040000040004100000100c1010c0000000c0000000cc00c30030004007c1000c000c00040000f4000000cc4000470000000001c0c00c0003c7000000000000c0004030c0000000c4c01300000c000100000400c0017000cc0000c0003c030004000000400300cf004000000000004c004000c4404000000403c0000c000cc000013000c0c0001300c1000000000000000010f4010000c00000000000c443300000c4c04000d0c700000001c4000030004010000040400000c00010010100000000340000000c0300000040000000000000c4040c0440c040400f0004400000c0000c444c0000c400000400c0c1c0047cc0004040000031100110d40c110403000030040004000100000400c000001cc300000000040000c0000000c00040430cf4c040030001004041c30000400c40010040c0c40300003cc300000100c000000000d000000040c0000400034c0000041c0c00004114140f040c00000044030300000400c4050000ccc000cc40040004000c4004000000c400000303004c000c0030400000004c004000400000000010043400010000400000c000403000410000c3000000000013fd40033c00c00c43c010400001000000000000040104404000403cc43404000004c7040000000c0000404000f00f040000c00c04c0040c0030030c0000c0000d0c3014044100010000000000000000300000000000000000004300c0000000c4000000004100c0f000010c700c000100000000404700c0000000000c0000003000004f0c0000c000000000010400c00000007000030000040400005c00000007003000300c0001300c1000c004000330000000030c000c0140c0000400000000c03000010070000000300cc00040c000c0000000300030000100c00000000500100000c1000c0000300c00000000000473404044030400300c0000000400014003ccc0c000000000000c00030040300013000300000000410000400000000000440000c44100c0c047000000f0cc0001d000c00001c4000110400300001400000053c0000c00c0000000c00000000d001000c00c0000400000000cc034c300c0000000c000c0c000404c000000c4c4c00100000401c000130000000300004100f40040000000000414000000c0000000;
rom_uints[472] = 8192'hc030300c000000c330003004003370300000001030c00000d1110000c030010001c01000d000c000d04000500003103c0000c01030004000400000005070000001077070300000c0000147c0001041003000000410331000003040000030100004c0100030000000010104c03400000030000000c340000000c00030000cc000304000400000f000403000c000001100000000001000c040000000700401033004d0400000000003030c00300c00c0003740000004c0070000000000314000300070000000c000003000000000700000040c300001003000000030000000cc001c00c01000c0004000000c047030d00c01004300500000c00000300010000c00304040011c0004040300340010000c000400000030300c103100c004c000c0c15000000000000040000004007000000034000000101400dc100000c0000000300000300014d000300030010300000030c004070000003030000c000000000010000c0470000030c0300050000130000000301030c004000010f0c000000044c0341000313c0030303000017030347c000040000000000100011030000030c0304c00f0f0000001c0cc1404c01030000100304c1430f1410c10f000000c0c00004040c0001000005070000010040300c041000000030cc0301000100000cc100000001cc0c000741100f4c070100030c410000030000030300000000000c47c0300300d00300030c00033c0011c000014040040030034000000d1c0000070c00000030010130000000000001030c000004d000003000010000f0001040000c5330c30401000000000001000000100000000011030404000000704c040d00010f40000001001000700000004000c010010c0300000c0300070701c003c010000011030000000007030c0003000043000003073000000f00400cc00300000000cc04030400404f01c04300000f3000030d03000f03400000100c00010c0cc00001c000103000010007300000030f00001400400000033cc00043010100c1cc1d330003030c030100c0030000074c4000030344c700000010070040000c0104c0cd00000001c74f00013000030400c700000c0c100001000004000003031f07010000c00d0000000c00043000004000000004000003103000070cc0040000070031c0000c03000000c00030500014030030070041cc00000103404301003f400000c0000d400000000000c000001003c0310000c01c000304000400000104013103030011030400030d0103030000000dc00300d043030c00040000000c00c00000000001010003000000000c0cc4010c0000ccc3000001030030c000000c030000040000c00013c4443000300100000000000000000030030300030c40000000000040000000100110c11110044c0c000d0300300000000300010010050000010;
rom_uints[473] = 8192'h5030c000c300134c0c40003ccf0030c3f30401000c0c00300000030040000c0000030030000c0000001110005000140030043700043d047cc000c0337000c004404d00303014075c100040cd00c000c500300c410300c4000cc1300c07000c0000003340000030f030f000c030c0037040c030c0130000000c00301dcf100cfdd470400400000d00c0300003703033300000c0000c40113c3c0c3034047c04c433101300100000000000043114143c10000030000c0040101040011d4500000c133040c0300ccc10c4c0004100043dc0405070100c3414401004000034007c007cc00c30101cd0000044401004730300074001000010003c0000c000c0000c70034040111151c010304000000030d304c440000ccc000040010000cc0c44043d3000000030c0c000c14c000453040030c0c0cf100110300040000fc13030c051700400347001000f0003f003400c0000f00cdf077d003ff0c4441040c4c30000fc0040fc4014000cc4000c0c3141400c0000c00031c744000c107c304004c0045030300dc0c0c0000c0007004000fc10000430053004c0000030103c0000cc0004f000000000c3dc003cccfc040500104000000010fc70001cc000414000001cd0d0400404c0dd3000300fcc0040c34c01010400fc00003000d04c0003f000ccc00000100c130c0010d4000c00401400c01403d000040c34004000001001333ccd04003cc030000000000013001c100c0c0c00030003000030000030c000ccc3d47004034cc400c000c10140001c0c00f033000000c1430000c0c00170003003000c04d303304000040400c41f00000fc00cc01010100011104c33300cc00c314100c04010300d444c0c07c5300000011c010c03c4000034000000007cf0003000000013400c1c0f4001050dc110400c0d3400c004300d300c030000f034000000000017300c1040047034c00001c3004004c0f0d070300040334c433d0003000010401c0000f03430400010301c301400c3304300f110701034f010500c310000040400000c040010c03440004031000030c50010000300004030000000300400c03c0404c030000030c33004000000400000c1300c1c110cc44004704001010040000f1c047c0c34100c0000404000c01f0000c3f10005c30014dcfcc0d400c070cc00000150000014001c0440000070c030107000003133000000003030d0100c135404c000004000c004c000c00cc00400000c170001c430040d00fc1c00000004300031100c10c00c50c03cc14000340000040400c000001d00c40c1001d0103cc4c001750033000c4c100010f00410007040010300300500004450c0c013070cd0340000103400c30c0040101c7010c40040c000c003303dc00000f03000010000131c00c30440000000030cc110000130340413d01c0000140c04700;
rom_uints[474] = 8192'h70004000d000300051c3400540400f00d103004033000143010400c30004000100c0035100000003004d0011c1030d3100d3000000cd03401003c0010c0001030140005000050000000010140000000f004000c031c13c00cc10107140d303c30070030400c00f400c001000007133010000000100000144000104014c40c300104f4c00000300c0c0000000c000031300500000000000400000040001013cc0040f130010c0400300110400000c00440000000000100c40000000c000000c0005000c400000430005040033000045400c000c30000040c000000443007000c00103030300c00040000100311ffc0003f7c0c1014000000c0004c00030000004041304400000c003000000d04c0300000c0f034c1013c33000c001c44100303050314000c0c04701d00073d03001c10014cc04000013c0000301d000cd000000c0013004c045040001000344010000000003c300cc1300cf00f0c440c1011000000000001cc0000d0c000000030003c10c01d100030000034004550041c1cc00c0454c00101700030104010001000174c0000030130000030310400005470004000d0004400500010303011103cc0c000f13f0014403000107410d00000003301305310300000001004701000c00100304100000300403c700404004400fcf05c5040004000333505001403004d00000c00030c00010010000c000000cc0034100d0031f330000430340010c03030c404cc01f0f01000000cfc00400d0c44030c0c00c03000c1000000370307000440c000010100010400053cf10000000050cc040c03000cc0c001010005001ccc101c000000004470000041000000340c04000c34500010d014c000004c304c30100001c00c1440000000cc100c41000400000414034c0004100d01303000c05711075c3fd10010303000400400c0000c3004d0040010413c3c0000000fcc334c0c31dc04000030000430000c300005030ccc30443000000040dc04003c300d10101000303cf0000000343c1000c00c000100000410431cc04c000000dc0c50400c7c41010000033110000440c503c00100003000000c30000500c0301c1400f0000c1400500000d10034000c000c700000043000040101301100000f00000440000c01c03c7ddf1010001c34c00c005004c007044300c00000c01340401c0403c400c1001100033000c000cc000c30001c444c00c34c00040cc00d000030c000d000000030000000c03000c0000000d40040d013073c0001000030001000cc0c0030f0000d3000030100c030003000000c0000001c3010003100000040000c00100001d00417100d00d000100000100dc00040144c00043001c00004404c1330040000c0f00010000000000000c030303000c504c00c404011cc00ccc000000010134104001c00000033100d040c00300c0;
rom_uints[475] = 8192'h400400c400000040000007000010100000000000030000000400004c00000000001d1000300cc0001000040000103430000c300c04044c0100400cc00000000c00031004000000000000001000040001c0010000000000000400000000000004101000000c00c0340000040100304000000000010000d10001000000000000400f0000000007000000000000000c00300001000c0c4c010c00000c001044000000000000000400000500030c00040000433000000cc0c04000001fc00000000004030000000c01000100cc0004000c0000040000043c000003000c3400100c000000000000000000000c11003c000000050404110000100004000110000c000f0004300c0000c40000000000001c0001000000000c00000000040d0004c4000000d00034040000000000c030040c04000000000150000c0c0001000000000c04000404001000000c00000004c0c004031000003010c1344004400034040c030c00040cc0104000000c00000c0c04040404000100000000003d000010000005040340000430000100c5000c0000cccc000500500004000c304000040000010cf000300330000400000c0000040c000030000c00000000040000c0000c0c04404504000004000000c3000401000000405f000001000c040000c00043000c31c0c0040c0c003001004f0100110d000430000c00f00004000000000000003000000c0000000040010c0c00000000f00cc1010000004c000000000404010007000000c10000130000000000c0101001d000000000040000000000300345c00000000c00030c40000c00000003d00040111011003304000403000c140000001c0c000f000011100140100004d40000040c0c10000110005037c0040001040000000000c0c1000000130c011100170400c000c04000300c0001c40c000000000000000030c400000c04000d4cc00400003100100000c0000c00100001101000400005040c00000000000c1400070000003004040c000007cc0c04404c040000000010c0000000000c0100000000043100010000030cc000000000c000c0010cc030040000000004000000000004000c03040c00000000000100000300010300000040100000000030000c0000c0000000000000cc05c004c0000c0c000c000c0300004414000003003c00000430050d00000c00010000000010f001000000010000001000000000300c0000040100000103000003c0300000000000c000000c0000f4144400400000000103001c0000040c0011000c00300fc00000400100cc04000043c00fc40400001000040c1400000000000300d0000c0103000c00000440001400104c401c000100000400100000003c001001000000440c0000c1051004c03000000011040000040c000004000d4000000410000c00003c000003000003000;
rom_uints[476] = 8192'h7030000440037c00f500000004040f403031030404033f3c00110f0010701003001300f1031cc03100041030c00c0340cd300cc1703013d4001403000c030c000030100c00103030030030100300070700000174100173c430c0150033d00704000705f03f00f0341c4cc00000f00301c00410001044c341013130c0034000001f314c000000001300d0003010004031000000000030300073000c00711037101533f0110007c5d1000304000110005c0145cc00000c000000300010f70c000000353011f0305000d00003000003f0077f000f00334301044f74c0c0c14d3010000f0000133001c00100004700030c0f701030170034000001f010001000000050004c004c00c40513010dc4c007c03000000050003c400cc707011333010f3400040c000013000301000003010050000c101dcc71c3004057c1400c3f03d03c30100ccd01f54c034f0c0013110104f0035d0013374c01f304c41dc000000000c30c4000434401fd10000d010000001410c100000c04004301340c0c0c0114c11333471143004330410c1c401c01430f0d0041003400013004d0c00000000c000000c113301314d0001033c001c1c34c3133c470d7f0031100000400035cc3d1d0110300005300070c000cc0440000005c0010c0f0000d330c3340f3101000c31c4c0000043434c11741c50f00c40c0d5400000d000c11c310310c333011304c00c3700000000d07f3350c31f00c0d37c0c0054001010c010303c03c01300341f50400001c73000300d0000007c300c00d0f5003040cc40300404004410000340c053130f30d00000d000d30111f00500130001c500d03000051104c05040c34033010d001330030314010300f0dc3c0133010c103474101c00000000d0d1c0103c40000040c000100307001401031040300070c0000430f003000004001011700c01c14c110007074335dc0c0000c101c113700000000571101cd430f1011014310400400000301000c0cc00004301001c03f1f0143c030070101cc0007010300005c0103f0c30040c10000117004c01f00114f005d03000000100033130f301000014300dd7570f00100cd0c04c11040c0010cc333000003c30fc10100d00cf55300003000703300d10c010400130c030c47110cfc001031040453c101030043331434130301000330f5c01300300c03010411034d0071030070000073005340f00003730d00350d0000703400d000c3000f001030c013c55c01c1000110400f304f0000004c0004f000400c000c0301010f0301cfc00333340c3000c000c03013500000403300430014010d000001003000047100c30040c0f0000040004000304cf703105c3c1c0000f3040000c00330cf5000301030410d40100400110103300000d1d001300c35130104001403530000300c001001003fc040000c0000;
rom_uints[477] = 8192'h1c4000401140001000000000000c340000000c100040000030d0000df3004000403d0c00c00000000000000001cc000000040000c0705000000c00c010300c400f0f0000300c1000040c3c00000c000c34304040307000c03c0030000343000400c0100404c0000c43004c00cfc0000cc0c00003003cc004300cf03d10c000003000100000014000400cd04000c3c00c040c000000003000f0400c0010000040c400000000c000c000001040100030440440400c0c30c0c04031004000004000f000400040003030400030100c4c004034c540400c030300043c0033100100c0100010c7000000000001104440043000cd004000c03400c00040001000003040c04400004470100040c0f430d000100c00f3c10c00030403000040400011400010000c0c004040000007c00000401000007cd004400004003c43c0c000000cc07cf00000c01000cf30c000c00000000d0040c0100000c004034000c04470000300c04d00001000033004040ccc0300000000c0cc000c000474f00030000071100c410d3030000f0c000000304c310000000010000c400c00f00000040c000d301040030c0000000c000000040c3100000130c00f0003000c00c000010c300c004040d0c00c00c00000000c100005f0d0c0000cc0c0ccd000c04040c0f00000004004f4d0c01000c0c0000c00000c0c1c700000d040c00400000000c001c0c034400cc00030300000100010c30000fcf03004c000c030d00007344400400c440034000f0c00004000c4000040cc0000c00c0000000000100c0c400cc0004000c0c0340400000c000000c0d04010000010440c0400c00400000000000000041c44f00c03c000001000000030000000c040c1001c00c000000070000310040040c40f0400c0400300100000dc4040010cfc10f0300c0c0c004000c044330000c0400000c0000c14000000000400001000004403000040000000000010000000d000000000000000000c0004000c00000c00c0000400400003000100ccc0c0300c300000004400f0c0000001704000c040000000000000f00f000c000c000c4000d0000c054050040004cc4c00000f00000cf0c0cc0c00000003000003004000100000400000000000c0000000d030003000c0c05c1044000004000170030004c1400000c030003000400040c400c03000300030c0400c03cc0c0000000400f000403000400400000030000000c00400001004c04cf0c0c4404040000000f000014c0000000c0000000000001dc0400013100030100d00c00c530c000c014000054003000040000010000000004c4443000745003000001000c00000000000011440c0c140ccdc0000440010340c44000cc70000404c0c030001c00400000c00f0000c000310440404043010000000c000000000100000103c400000000000004;
rom_uints[478] = 8192'h104004c7040453000000047003cc50103d40003003c003010c1c0004040030003c001015100000f0010441c0010c300000d040001c7d3330000004104000030003140000000d7400001100500101300000074cdcd00cf30103dc3000c00303c4370300400300000040d000000c00000cc0f040041000301c530c40033c040c0c300c0030c00330303000000004003033000010000000104003c00d44c000030130c1400f0001043c00350000c43431040000000010c43010404033c1004044004344000004001140001007040cc0fc00540370410000045000340041004303000700040f10034004400c011c110ff00000c03400400000000030000c00041000000441010300010001100330000710040cc4000000cf430100401c3740000011043000054c007000003000410f0000f4000050010300000c00c44c000000034f30040c03001401100000000330c000040000043c00100cc13dc3001c00130f0030c1430040c3000d45c303000f11100c00c003400410c3074014000c310301c3f30dcc3040000c0130403000004000040040000c0070407000000000400030c040c00303000d30030440040c000010070007704c00053000330c0000005d000f4c10d000400c333054000000040034001c00f0044430c00fc1134010d010000000000430000014000000741c500351c00030040040000011c00c034000c710300c011c30444000030017001070030c4013000050000303400504000050c00007003000470cd000000c0c105c040c00010300135133010433c0430c000370010c33033440440011000004000503044401004000040c1030301044000000041c0001000dc0d01300c000cf40100100310443c01000305041c004f4000f04445000000c0000030c070414544001030c0330ccc1040c00c4000443401100433101030451100000dc000cc001c3500001c014000c041000500300400047000000031041d330000000005700000013105000510010c0103cc70300dc0c00f0f1100000003c0f300000c000300cc100d03fc10040313c0000001c400010000000000c0040100c0107c403170300000c30550034000403000350001140cc005cc0300071001000000017000c000070c04c000000073000c0400000300400f004001c010f00343d0000c44c1c00100dc300000044030c103cc010110400000000d1c03004400100001000000c00070000000c0000cc000303000300f0400d030050040cc00dc10344510000fc000dd004040010000004430331d100030007000c40003f00741f70100000140001473c10700400cc03300c00000004000c00001101100c0030474c000700733c1007005cf04d00140cc0c01010304040030400074000d10000000d00001c30000030004300101100000044100d01c00441007c0c00000;
rom_uints[479] = 8192'h103c0000c000000340c000010000004000cf030014001f0000000510010001100035003130c0000011000000f0000000340000000fc000033410000003300000000003cc0c000000000010001100040300013ff3700cc3040c0d0133000431301033000305000fc05d0c3c00c10301000141c133c433010010cd00c00c43000371000f03040300f00001000310000300000000010000000c33c100000000540d0c140000030030300000004030040007000c03050001040005300011dd017300004d0c00000000000000010f03000c10c00cfc1030010001000030774000013403300c000103c30c000100d700dc000000010104400000010000050007500000000101030003700f0c1430011043040303534000010000c00cc00004d000000c40033000103513130000030c03033c10340140300f003000c10cc000c143040000040300010000000f0030f0344301c0110500070040003043003330c300100fc100440010043000c1030111f0110f30000300040301100f000730c000000000044000044400c34303040000c04c000300000000010014300571040f0001030310cf4300033300f00400000050074007100103135435400107f00101004340514004007010300000007134031300000475400103000f040000400f0100500073031003f4100f004c07010c0073040000c0000003004000c13d004dc0035005411000330140000300010003004040040001c0c000034c000000030f00c0c000330000301403030100000003cfc43043014003d0000100040037130004cd000c030c00150000cc000003030f3014c00101000004c007300003034c30004050c3000c3544010000000300030501000c1100f0000000040003004304c0000030c1f0010040143003100c0100000013104001c10001073010100100c00000733c10c30300010440004000001030330f0000107530010c00c3cdcc30000c00000501c1d00310000300000c000300000030000400003400c1000430000f003000070c3000003d00d7000c3000003c30000000000000010031000000014040000011000c03c0cc0300f10d300700000c00033100334401300c0c0513100d0100c101300043c300000f30000c01010000040000cd000303000030000441330310010c0700f003000300c000000100000300100c00c3000c010010014c4cc000000000400400100133d0000000007000030301000003007300017c01050c0000030103030300d00c000000300004010003040000010040044030004004141101300c030000143043c100400003010004f507cd04000035430c0c3040030c00330005d50007030030050043c103c0014340c150000000c003000000044f43070000431c000305010131404400cc304401000000030007000300010c3040c3c3000400000000;
rom_uints[480] = 8192'h100000000010000030000c00000c000300000c1030040000000c040c0c0c00100100000000c00000001003f000c000c100003c004000104000cc000370000000000333000000000000010cc00000c00000000c003000400000004000000000000cfc0410000300040cc03000041033400000000004000c0000401000400000003034000000c000c0303030001000004000001000000000000c1000000001000c000040000c30c0300000100000c0000000411400000000000400001440f00010000000000000c05400300004c400300000c030111054000000c004300010000010f0000c30000c0c1000300010f0000000103c40301000000000003000100000f0101000c03000040400000044c40000040000000014d00040c01334104000000030000000f00400000000100000000000000040000030004004000cc00c000000400010c004001040001003000000c400000000c0300130c01040000000c000000001d4c3cc00304040001000140000040c040000500000303000000001100004c00000000000000030000400000003300000000000c000000000000c00000010040040000000500000c0000014400c00000000d4f000003000004004300040c04000c000f03cfc0000c000000c000400004040300f313000d1140013c000c0040c00000000000030010c34c0c00000003004c100100010003000003300000000000040c00c0000cc10000004000030d00003000007000000000c04000400040c01400300300000004010001000000c000010000000c0300401d0000004c00000000010d004000003000030004400c0001070c0003000040300000004410c100c3000004500001000d0000000000c01f00c307300c00000000000001c0000000050f01000c4004400f4040010000000000000000000100000000000004004000000000400000040c00000300000004000000000000000c000000000000000440000040410040c0030000340300005000c04000c0001000000103000f00074400000000040cc000000c0000000004000400400000000000000000c1034000004c00c30d000000004400030000000c000c000007000300c000040c0001000c0400000000000000000000000004c44300000001400000040000c0000c00100001c041040c03000400000000000c0100000100003441300044c340c00040c1000c000000010004000700040000000000000c0c0303000033f3c00000000100301c00000000000003000300040001000cc3000c000c400004000c01000007000300000000f0c0000000000000c00000000c0000000004000000000003000030c30300c0410c0c070c0c00000c0c1003000100000000000040000303000c0003000000000000030100c3003000010c000c0000000003000c00000040c70c03000c00;
rom_uints[481] = 8192'h41100000030000004100c003000000c340000140c10c30030000c0000400040000c3c010c0010c000001030000030c40000747c001040c01004300404001000000c0cc0040000000000c000000000000010d00cc4cc0000000401cc00cc0000c4441000003c00cc000030300c14c0c0c00030000000ccc000040000440000003c30704c0003000c00f0103c041000000400000000c004001c0000000c1000301040000000c0003000cc000041c004501c301cc00000100000010c37100c00404c001c040000440c401000073c50040c3040c44c500404c000000c0c5114000c10740030c0cc0030300004d30cc3c070d0051c300c0400000000300c340400310001c01010cc0000001034047000c0003400000c1050310000f000f00410300700040000403c303330100c000000001000000070000010000000003400040000000000c0c00404100c140c1c000100d070f0301030040004fc0454043000000000404070c004c0cc0c10001d440000fc0434003030cf50cc000d0000000030300c300d0c0000000cd5303000000c0c4cf000040000000000c04400c000000000040c00400030007c00300000403410045000144030c00cc04000f01010044c0000000000cc00001c10cc04000c00cc003000c000300c301c00340c004030104400000000141c100040000c00003000c40000d033300000f0001000000410300d00041030400c10403c0030400400300c44c014000dc00000103044340c04041003100030000000f00000300040403c00003dc000100000000c00700004003c111000030c0ccc00000000003c00000c00c000d4000c40303c04103c0030073030d0047040c00000c010000003001400cc1340d000300c000c000c0000003c043000500004001004d000c000c0c00010c0d0c0c00c04c031300000000010004000fc00000000c0c00c40003430040030350d100500000f0cc0c400000d0011000cc000000c0000c0000c00000000cc000c00404000c4c0000c500040100010000030000d1010000ccc00cc00c0300330070010d00c000000003c4000053c001c1c00000c040c30000c14000004000c0004fc501c001c4c3000c0dfc0000c04c0347400001000400004000700300c000c30300400103c340030c3f41c3010044000c0c00c4000000c0c00000c0004000000401000000004003c0074400000100030c0040c00c01000100400341030043010500030400000c40d103000400000500000003c0000003c00c400101030000c0c000044c000d000303401001000100000300c000c300044000c00000c0000400000343000d10000000010440000c0000000000430000ffc40003004703c1400000010000400000000001000000c00f03050000000040c100000303c1440400000000c0000f000cc1cf000000c103c0000;
rom_uints[482] = 8192'h307000000030cc00007c0001300074000040010303c00004004000001340c00000c000c0c000c047000000007503d1000030430370004040c0c00003c00000044004c00400000040c00300300000d0c0000cf001010040c000c300400000103041400c04c00000340c700c0330100c40401040c04c34030040c00300004000000000dc0000c000c040c00004000000030c0000c0000c004cc40000004000000073000001000c41400010400030310000134300000003003000c00f000000004300d041c00000000cc0400c00001007d00004c004c7150f0000100300004000001000c04000043000c300000000d01000f000400300d00010000003000000c000000000c05031c040000050d01004004013400000030040030000007001001d3410000001c700f14000c040004000003100400100303040004000f10000d00003300310c00100c000050000100000114000003000050c00c00000d0c0c0c0004044030000d00c0000000000c030400f31c100c0000300000c03c400014040000f3cc0f000d00003000000001000001c1100004000004040cf0110004003004000c30cc00040000000013000000100c04000c003c003031000c00040000000c04c000100000400000000100003300000c003d400400330dc404100000110c0c1000003000300030103c0c0000003c0100c400010c0000000000000000033d0c040c0cc40d300d0c3000300033100c0001110433000000000000301c033c010f0c1c373ccc50c0000400cc11001001300c00003000c030000070300c00150000c000000c0000040c01000c400000700000040c0d0c3c0100000030013000000300000c000003000004000000000c13003000050f3c0040f00400004030000000000100c00c0c0c100000c00004000004000c3c000011003053004301000100000004014c0c0000000401040c040f003c01500010030004000430040433440000000c00000103000000f00000000000000c00400044c000000ccc00005cc03c1f400d0010f300000cc40c034004c01000000000300000031104000041cc004c00300f300000300c003000000005007c00000c0d0000000c0000000000004004030113010000cc0c0c340300000000c0400000103000000404000c0001030c0033c0000c030c0000000300000010004000100000003c00143c3005c000000307004cc0000c440400000050000030000040003000100c000100000403003100000c0004fc0114000000000c0000300c040c3000305c00100c0f000300000c0c000000330004000c030c330000103000001c00000c107110000000000001000c000700c000110c0000043c1000111c000c00d041000000000000040404000c000c040010004c000c0000001c000000000430504f4000000007c4000c103c0300000410;
rom_uints[483] = 8192'hc040f0000c0010004c004014040c0400f0000c1c304000000000000044131c004101cc10c00030003010001c000310cc1d13000000013304c04030f040030c30c443500c1d000c000003c4c35004003c0340003111503cc000100000040014300c101030000c0004c0031c001f40303c07c114f0031010100d3c401f14301001103c004c3000410010c00001305001330c0c001000103034d0001013040003040f30000003c4003010004000000c1000c003700004d003371000070330300130f0d0cc3c000070c0343157f330573730014c3d30000143c054003031100c0000c00c04340001300004001c14031c0030c7144410404000003000045c331c000403c0d0c30c3c03c000000c034000703030cc007400010000f313400c500030001c4c700050100004f0c43cc4000d03c000050c07000cc0003030340cdc443300fc0101d010405003000040013010c0000000040313040000c411101c0000fc103c4300103110071000c0503c04001030030c0c54300000000c70d000500f74f03c31040000301400001000070000c07410301430004004003c040400f4040033fcfd3014104cd500000c0c003403d0004014dc00f74000014000100400305004cd4010044c000004704000303030c00c10d03010003074300c0c00003c030c003c000c30cc3070300140c0304714c01770000cfc00c01c1010003001d404c000fc300017740c0404470040011431443c404430351004c00407101c040000140c30d00c000c000000100070d3403004007c5c701010301f0034dc0000300140f303f0f0300404103c0c74100c003100504c50f0040033f0300c140c00d44000700010000c500050100144140c40100030100144304004044400c0c00030000d43dd401450000000c033105c40010cc013170410100410f00000410017000430f40d10115d00fc01000000c00000440031d10040c04000101430fcdf5071000404013004010000001c004030040050cc44047f40c0040c000c4c440000007113000001040004301010040000d01000043004f03fc0000010400c0040f7000000045304005c1dc314007004033c0030030c000050340100c00c1000d0c000d0030373704430d0cc10040c30400033ccc430003170100c30000c03000c003cc0303030113c000001000c100d00310000000000000140c4f01004d00430101c00003c0000013035c00010001004004001100c430000300300f4f4ff1004cc00104000c00010100000003c10015013700037c430311070030000000c40c403c4000034000014310000c004004004010cc07c000500303c1000300000000000c1003011001c003c00010030003ccc3440300c3400cc30100c5010d0000c00000040c000000000003d00140c0c10f300000410401000000c00c0c0c03000c4c01000000;
rom_uints[484] = 8192'h10030000c100030037c0c330300000043d03000041000000110301c001c003010300c0fc0000030001c001f14010005500c00c013000034470000441fc40100000c013000001000cc0000015c00001130d050033010000000000c000400cd0c3410cc0001000f04000704330d03000003013000140c0c003003013000030100005000f0000c00000300001400100000d01c000300000000043000330304330100305035001c310100301000001000c00000070000030f0c311001041c433000001c403000001c0317cc30100010000c0300400401041001000000100340100c0000170c00c0000000000000cc513f3000310cc01000000040cc0030011000030001440c010400c0003000000300010300117040001c1004d000100100000404000130000001004c0000003100f1000400011c0c030d14300004c11104000000c0c054cc04000000031cd0300430000000400000043104000144001c0401014c0001c0054033040c00104f3c0d01000430030711040c0030410c30000000010307031000c011cc0d0000011000100d003c000c04000001010011350c004c40c00c04301000000400d00000041030c3000444000301010c00c010000c0000d030500040007c310c11400430003070004110d00410040003c43000000cf11000d4c300000c000c00307011113c04f10000300000071004000000003400001010303c141404004040300c0030003004c00c314101400c00000033c003d70d0000003400003300c030000000000003c00140030000010000003000000001000000cc404c00370c0041000000c000030400300030001c34000313100171000130000300401000c303000d40c100f17400001c0110004014c04400000034c100d004100070000d0140000c003c00000d11530000000c311010040040000c010c0405000f000444c07c000c303fc0033c0c300c00404031040300030d1010003c3c103c00000700300000000c0030031100300104041000cc030c0040700010d403000010c0000000000100f0104c003135300001043c01003f33c030c04000000300003100000100340c300010004000000404c70000000c00c0100400000c410001040033d03c0d0014000303030414000310400c00300014c000000c0140000007100c400c0300100014001034001004003400c03030cc0010300d0010300000403510fc0c00300010000c00000100000000040c04d0003030130d04000c10c01000304104340c0400300003103434c00000300d45d1404400cc13c004100000000000f00000000300001004011c035400000007100030000000030004000c00001000000d04c000003400000303000f001c4d00000000053410c00c000c010433000010000404c00003c100043040000001100c00001000041051000010010004003;
rom_uints[485] = 8192'h103000103c3c33000550130050000000f0000071f00010000010300100c340013033c300300100000000000030c0001000c003030000144100000000700300c000033030000f000f0000c0117103c30403000030cc11430000c0310730030c100040500004004000ccc0071003401310051004030043004000110c130004570001033f003003000000f100c000100430034c00000000d0f74300100cc33000000000110000010000000110c0dd000000c043010c00404440403010113fc00303030c0c0000c03030cc0000003000301310073301c30c01033303c30310100000c0d00000340000001030001001510000033f0313401000400030c040030100100303000003f00000c01330c0d13330c4005000043000000c0001c033511030010044030003c000310000051003000f00030100034001030000030040135d003000c1035d00503c4000000c74130010d01104c040000010003010303c0001110000000f1033300000c5c0004c10033070000151330000cc07030c330140100f5103000073000c30000003000f1000d4433000c4c00000dc1000c3103300000050513ff40430c0c0330033400130000100100000301d0003f00313c1010300010001c1013315c01300c0d003000000305c33c33000c00000f30030f03000c400c0ccc3413030c3000100000000000100c0054cd00c10313000dc000030d0dc10cc00003303c0c00c00004000003030c017141041333003003030010050d000f00011400000f44070cc0010133000d0340043f431005000400300410c404100c3c00000500330c0c003c03010c300f1000001c10030c330c000005000110001400303400000400000300000c000100c303030000030f0d3d000000330000003c000000010100310010100303100dd0010330301d10000003100003000101000d30005c1010300c07000041303301073000033d340c111c00033300000500030000031030110000030030f0000300030003c000430304000410c5d000000333000000300300000000030c0c1330cf0c00000011300cf00004310c01d00c03301303000003000f0004057d000000000700040c30040330030011100c03300c3413004c40000400033010000010010000030040000040034c0010000100030400000c1303030000030010000c0f10000c01000c0c0103030000040003000c03051c3c003010144c10c00001300001440000070330330001340303c303c0014401c034040c000d00000f40030014030705c0001c0103300003173c0330f0010007000013030004031c000003010100003100110300037c0530000000000000003100000000303c00030c0c0000040fcc01100c0004030110040f000c000030000100017001d0000c30001000111030000003030030000010000c1c010c330d000c073c0;
rom_uints[486] = 8192'h50010000037410031010101430010000141100000c0011100447140004313500005c03444000000003f00004031030347cd000010c040000010004031d0c001c31001100310000001000c03015000c300330000047030330000700050001c40043f0100d3401dc000f34cd000404c03300fd003c10d174000000f00304d0000047040c0004cc0014004413000007001f0017010400301c00c0310004c4000c04301c0107030c015000000003330401003000310400300001040c04011c0310000fc40c0c0000dc005c03441c1c040331000d0300f00100c1101cc30d3033000c1c0400000700000004310135304314cc0c34310040c40001104030000000003307001c0f00cc0f00003c00130101040103cdc33014c03101cc0504003500030300c1100000340c010000000c317c431c7c040300100000000d045c07c0310001000300030015140000000100100311007017400000140014403c14300000001300340c3001130400504000001300013030070001c43c40000c31c40c0500c01000301013041014304030700c310c77cd1400340000040401040430100c071000010c0f1100004000000000341c04010003000cc13007010f00010401301d74700370001030000731001440003c00330504c0003c3c0c333d00000c75035300701011004c043c00d30c03cc00000000040400010f0077300337f400040303c000301cd0c01030100104300301301d1701054510c033000f00010f7003f50500300c35010007100000030f0c0005011c00000c33000510c001000c14004010000c0000050c030340000c0014d100440504000c31000f01031c3c030c00033c010100d00004d40000003c14431100130000070404100014300c030c0730c0100004c03f0f001104010000140500405411000510354f54041d0400c1c004733001330000354000031c3d100501700071c10f071c3005340f44d40000100001041004010000001c004434f10500130411007c04c31014c300df0030300004040d3010030000003d4034000314003343f4003037c00330004f0030043c4000000074044400d0000313cd1510014414010c000c03f13d01340c340f001001000407100530310001001f0dc1001700051c0001310c000d4c0c47c004140f0c030030100030dd030004300100440c030010010010310004000ccf04ccc0330000000c00300c30400d014300c1100c3001f00007000c11cc0c040013310f0f000300000400040c0003c50404000c00040000341cc01000070430001300c0000300500f3050003033300333010400010031170000010010cc0504000d0000000000400000030030015010003503000c33004411000330001000000000303000001300c5403000043400000c071017030110033003403c0004151000040f1311000035100000;
rom_uints[487] = 8192'h3010004000c0000000cc040030111040df04000300000000007140d00d0301400070000173770000034700c130000000c0330c0c043f00040f054c030c0010000011c0001004033040001057cc0400003000034c00000010004305d00003c000000010300cc10c00000c031110400f100010000037000001000c300300043300cc350030003300300000000cd004100f000010000030040c0c1c000010400034101000300003c0c4f0005530000330000333000000000350430104003000000411003000cc003003fd1c03005c100c14407d03330c1100100040c0133d7400000c30000000cc040c0c011000040c00f003007514004000000c0004040000000c0011300003c0335c03003000510044cc400000000310003010000037c0c00c0c10043000003400040301300030040c0400431d0030000000000c0030f33104000001103f0301cc000c0010f3d0010003110c3430000403037300141c004040000c0000040cc00000c000c10d34c00003000000f50300113004c1d30000004400344000000010300000c0c000100010043000003000030400040000d010500400503f03000f300004000f300331030d04300c0010000000f00400c00040c0c10040d0c0400030040040c0340050101c4400100303c0c100010070770130000030303000004004300f30405c013000000f11303003c010340300000c0070f010011000f0c070cf0050001000010030343010c4300070003000000030001400001000037000c1f0000c0000140c0410000001f0000000730000740037043c003c0400040c3000c3000c0030000cd00000000000300004003030115d0400000100c17f030000f4f3c00000303033300300c030c00000033010c00003400400f0c0c00300014000001033cc003f4343040437d400373700c331cf000c3000010d3010303c0000d1003000111037333011031100331c0010000c004fc000354c00000003040100000000c0d01000004003cc04c0c500000300043345000030c414fc44c0000d40130301000034000333000c53000030003030030003c10010c0000c00300000000f07400c1c0c300c00000030c00d0400053000140300c34010c03003c00c30010000c30000000000000000300340740000f000000000000300003000310114f000c00030300cc10c000014f000130d4000310ccc03400000c00434730001004300d30030330010400410c00010340500000c1000100000000dc00100000001300c00c3001000000df007ff000000134c007000100c010440003000000010303c0010030c0500000003007000003c3040010010030000100001c01003000040c00013df300c0030c10c0030f000730303000000f00000000340000000440000000005003c000f331c0101033004000000c0c0001040c0430000003000;
rom_uints[488] = 8192'h3040000f004ccc114000c110000140000f4c300c0331dd000f000004401130000c000341cc000300000434770c033cf0301cc0000c3cc00000300130c0c01100103330d040c00cc0000770540000030c000000000cc3cf00015743340001c000000013300000d4c004c500070330cc330500003c0c400c03034c3c0fccd04004430707c033000cc000001030400d1c0cc000004004c0440cd430c04330f013443000000000000440000c0cc00d541c000114c40000030c4310130130fccc0000010c0000400004004430000cc40cc370c0001cc01400034c03d103cc4000000c00000004001044000340001c00f00cccf43f00c100100004010101114400000104000004c0030c0000000c003c00000d010005c0031030c141300cc03c0cc105500c000cc0000c0cc0000c430300d30000000033000000001000d00c00c030374040330c0041d0030c000c000c40c00031000000c35c0c0cdc0010c300010c10cd5000370440034c1003407114540f7c300000000c010ccc004554040003001000f0c0030400000d31c00c07000004041c003100000cc400104040fc444003044fc0001041c00f00444c0c00074000d00000730500c000c30c03400004d140751000310000040000351400c00141504c4404cc000040000334000004f414c0000000000300400c01d50c0000c100c00000000100010c7dc51040030000000c414100c700010044004044307040d350c00040400001010c300007030404040030010c0304c3030f300010c00310000040071040000cc00010000c0114400331cf34004cc34000000f3c10000000000c400c7000c14c40ccd0004041704000034c3000cc0000c000340c0100040100040cf0c01440c04100003003444f000000000c00c04143003c00005000c0c00100155114c0d1d00401000340000010004c0301040fc0400c4c0c000f00300410f0041fcc040043000000c40c00001f10100000103040400c0303c40101100040070000404400c0f4004040000c000d0c300f00040040100c5370cc000cccfc0040f0fdd300d10c0030000100004c3100000c44000f00cc0040d40040c00000c0c00c04cc300000c040000040004400c04000d000040c30d000043100f3000403003ff00330000100f04c401103c30000c0000c00430300340c00cf001044000c00c4c001400cf3c300ccc040c00c01003404f0400000cc00015004000004f0007c0c0000dc0c0c41044033f00f00ccc3c000430300000000100f44c00000cc4dc400501011d00000400cd003340040c1010f00f10cff000051c00c000400553440c0041cc03f400000000000c00100d040d00000d4110f044c4000c3f0400cf004330c0000f003300f000c011010300c000000004000000003000034000005005c0400001500c00c0d000000770c0000000;
rom_uints[489] = 8192'h4c0000c03001030303c0017d00005001000c000403300000c7400d0040c300000401400f010000c040004c0000c00030003010030c00303104000000000100c000011c00c000c0000001374003c00731000d03030300c00c0713000401c303007100f310003d000500c100c470c00110c000c00300033303711103040300001340c1010000000c00110001010000000000011000033000030013300040c0010103010000031c010110000003cf000300430100000043041000000453070307c400c0310000001d030c00000000f004c071113150000004530d0d3000011010010000030c00d000001700f313f10330030d00f400000000030030400001c004030001300030001131010dd3c40f000000fc30f340030100c30300017003303013730300104033000003f03014c00400000000030c1000c0000340404104070011001071cc000030004c3033300033003070f00c34100f43c301100001c0c40c0000f100530d330000000d0d310f5134000001034d03c030000301404c003030c3033040030c4c0f003040c051000300c0000100c0011053000140000014c00330310301c0300000004000000001101000005103040303310700c100000d534d0331301000001c0301c0000003030000170441034301f00330331000015141134c0030000000c30c3004c303000c3c11441000040400400500030003101c0400d000c04135cd00000304f0dc00010030000503140c000000c00030301100c300000003040d0000c101c03003070013133030335030f300430345007f100040c0000131310301cc0003f00000c05040407c040000000000300003130000000c04101000000040011300003c01000103010c40000c30030100000000530d000010103103030300000100031031c003000000400003710731000010c0003000c0c030c0413400004c0003000003000003001f1034000c10000c0c410303004001c00d00000300003c4071000c0114407c00100433c030c00c0003000f1040c03343400030c0c330100000010000300000c0350700d00001114031000c304010330030c0c333000c0c017100130000003104100040410000000001030007410c1000110100000c01313104d1000000000d0000030030004d011307c0cf0100003000003000000304c0000110143040000000400c0001c00d400003030c00000330100003c4c30000001c100c0100c00040003300000050000404cf00001000000700c0d0003100003c704071003070400c100014113041004000004000000000000000010333f0c0c3000041100001000101000030000f00170301ccc0000001010300c0011f403c4d0101314003400000015300000100400010100331000f0000001000100001030030010001710700405003003003711000103030c10400010000;
rom_uints[490] = 8192'h3c000004003000000300010c0300c40130003000031300107f030001300c0000000010000000000000000300000cc00c00300000300350000c0000d10000c0030003000000000c000035040310404001040000101000000000301400040300300343c0c0100000000051100003c000700000000000000000c1130000400100cc00000000000040000000c0c0000000003000000003000303000311003005000000000000000c0c00130331d10000330010cc030000000301f00000070310000000000c000043001010010000001f10030001010c011100030c010437070000c4330010f3013001c00c00000c043f0000004c040033000000000001003000000300000000001133303100400010c700013c0000100030011450003013300cd000003c000303000000000000f00010004000000c001100000000040330000030301003003050040000000073400000010c310c30334103000000310103070030001300040031000100f000000cc0c000003c0000cc40c30000d00100c0000000000000010300300000c70000c00303000000c0000000050430010c0000c0004333c00000001104010001300000103c000c0000c010141000c50700000cc4100000000c700003030303c001004c0001140c00000000c005010000f0d1340d0100030000000310143c140003033001000043000c110000000001000017c11400c0c000000430013013100300d000c0001003000000c11103000001000030d0c5c3c0030000007015000000000000c400000040100300304f300344001003000300010040010000c000f004000003c030c00c00003300c00001000300300400031333410030034001000010000300c04403000003c000000003c0300000000000f100040000000000043343c0c0c0c43400000430c00004100000003000300000000c3c0040c1000000030030010007001131c000030000030ff1c0304301000000100000030000000000000001000001140340000030000133030000304c000000300000000000034000000000303c40000000043c0000410300010c0130030300cc000000c10100000000030000000c000000400003001000000030030430001cc1d100000001000003fc000000c001000300041000000100000000c001c0c0c000313000300000000000d000000301c000d00000000c03000c100000000000000c000cc0130000017004000070000c0004105110000010000c010044003000300000000c000301030105000000000004c0c001c3000c7001000004100000000000000c00500014c000000003c1000000001001341000c0100000c0000000d10000040010000c0000c0c130111543010000000100000c00c0003304001300000004000030010001003000300403f1010004013000000000010003000301000000;
rom_uints[491] = 8192'h40c0c140000004030000000f000000441000000110014000030140100cc0003015700300333004010300434000400003c13310c0c347ccf41c0000101000000000c03003011c00114001400c1400c00000dc030d000100f070c3400003000001035f100d70130c000400000c01001000000000004c4c030033300c034000300031304030130000700d030330d0400000034010300000c3030003f00003010340000c0000010f40000000000000c00c1000c00000004000c00000011050c000c1c030c00000031004370041d001100011000000004000413100d30c3000f104001000000113c0010001f30cf4f0110500034001400030000000404c40c00000fcccc00000d0104073000003301000000041c0300040000000c1130c0000000041000c10000000030000c3f070000510070000000040000001300003700304004c000cc00c03404c000300070100010101c301c300300701003c0000430310004000fccc0010030000c0004000c1c0d00000030304c05c003c03004400000000040030c04030404330100000011300c0470000300000005003dc30f000c1000c00c0d0c1000300404400004300051010c000103030c0000300100000340f01041c34100030c030400010c000000c00c1031c040104c001000000030000d04400400c730000000c0040c400000000304003040000d000f7010001303041c0011331c500d30000f340000cc010300000030c0305c01031c0300107000f1c0010140c100440111d55103030004000000300c343300001000000c300100031000301c00000d0000401003000050000001000000c01f000c10000000f30c30c450000c01010303030000103000c410300000001431014100300000000300000100300000000414000000c70100040003000004d113dc0c0100111001330c303f11100c40010004c30c03c013d00041001c0053170c000300010000000c000f005d0403110000100100003000000c0500014400040c0000300130133c000007030c44070500000010cf3374100130000047005004500cc3000005c010033700011c0030040c00310d3400030100004400000c00300000000003000000000307ccf00010cc310000c01d3d3c00c501cd0cc00c03000c304400030000c1000c3c3000000040c4000300000f300314100044cc01300c003000003300035000140000dc370d00000000103d00000f00100dc1000100000001000430114144340000304c703c3113c31300007f0013000430050c0c1c050704000000000005050070000f0014010c03503410000010000101000000f0001000d000000c00001c530001d0303044000000c004000c010000c0031f30001013000f00c40404400401110333003c0000000000f3c000003000030c410000f303c010cc001c10cc3050001000f000;
rom_uints[492] = 8192'h400300050704c000100f00030440f1fdd400000c0d0c03000c451000c003cd0000000533007404000c30057540cc70000050000c0c0c0c00c000c0c313c010c4000371000dc00400c00000fc504c0d040000000d4c0d43040000c000010c0140c70400c00c00104c070f0000075f00030c400f00014c030001d40d0c00013300000fcc0500100f040d0000c00003c4041400c400000000c000cd3000c00c003403c034f1dff334c40c10040cf0070000010ccc400400711000100c400100cc00d4c0c004c00c0c00000d0cc0c0d1cf4d00030300000004c1dc0fcdc000f00300c4c000400000c0040100003ccc705c0013015c700000001401000044000000cd00310c0304044400c0d40f7311500010107d0fc0d0d1c40c400400c05404040c440000000fc010c040103c3c71c1cc0000100c0140300140300c00100c400000000cd10004410c0cd0d3430d04001000c300004c003310dc403400c0d04003c01330000cc434044000350540000f1030031cc40410400040c5003000141043000d0cc003000000001fc400cc00c01cc410053c0000044004c0f00c5010004000c1fc300f030000c00500010704cc0c0700c70710f0001700d0c0004c00000000000040404c0000440cc030cc400404c7d3f030440cc030304403140000d00107c0304c000000400c0cc43000d4300000c00307d0000401003003c004d0500010fc0f00c0cf04ccc450c0d703c300c00100c017d50100c000100000c1c00cc05505500104c0014000000f0003cccc000003030c0011d4404ccc0100f47000c00405c003f00701c00000c050100c000404d4041000d41c4c0c300000cf30301414c04000000040c0407103f0dcc00c00004713c013010400000c03c045d003000f000c0c0010000c00545400c30dc0004c001c3c0110000d000400cf0c01130c040c500c31033001700c400000003007054cccf04cc0700401441000401414100000c0fc4000014001c0c0004c0000c404043fdc00400000c0040040074c1c3000000004cd0000040004003c410004d0cc00ddc70003c4000000ff000c5c3010c7c0000f0430c140d0070010d00c7000f0f30440104d04c0000c3340c0fd0004d4f00c0000001000104103540c0130000c0ccc01cc14140404001c0001c0d0cc000c00c30c33003c0dc040d400c30c000c00c0c00c04700c00140000000c0000ccc40c0c0c400003f00d0005d040041000c003f0044003cc0010040340000014c741c0000000000004530100000110c004d000c3c010c040004ccc001d5341c40410130000403d14d30010c4000cc003000400034d400c0100000010000037c40c017033c4370404d00ccc74c00c4c00400410000c01040d700514c01343000034c00d031000c00400c04c0cc01004010ccc300143540040f01f100c0700c0400;
rom_uints[493] = 8192'h400000000000300000c0000c300340000010000030000000c0000050000000000000040000000100070c0001c14405100000000000100001c0400000c0404000300000c0034c000031c00000000000000000cc0000c000000000000c0c400ccc0000000000043400000001100000c00000403300000000400070004c400000c400c000c00000001000003000131000000000000c00004000c000405000000100c000000100c043000041000c00004300c0000040d04030000000000000413d00040000004000c0110000c004c0c0cc0000003004003c33000003c1000c00000000c0cc0c000000000300030003000700d40001d000100000070000c00c0330000040300000c000c040000000c000014000400100f0c0100000001000000003003000004000400f004030004cc0000100040300c0000040c400001c000300000000000000000040400003040004041000004004c0400d1000c000000c000040340103300000034100000000000d0000004c00000030c00c310400000c000000010304030040040400004000004500000040400007400d400000000000000c04cd00c030c003000000000c03c41000000000ccc000030000000000000003c004c40000100000000c00000140000007000cc110004313004001000c400330c0000000004300000000410000000000001004004c000400000000000133000040c0c0040003000000000004000000c04000000000400540004000cc103c003000d00000000f40c140040040030000c000000300000010040003413300000401040003300c00004004000000000140000000c000000000c0000c444000c0000c3000000000000c0000cc00c00000010000000c00040c004440340100000000000040d700000034003c0c00000000040000cc01c04003400c000000000c0044000003440000f000c00cc0003000cc000c10c4000000000000010000300c4000000300cc0c0300000000300003040030400000c000000000c000000000000000104000000000c00c0000003040c4010000c0000004000300100001031000400700000000300000cc000700004440c00030000d0000000040300040c0c000300000000c0000001000100000033001c00000000001030004000000c0014100c404030007000000c001c0040000c000c3000300000000c040400300010000000c0031000c400c000300000000000004000000000000c000404030c0044000000000004000000400000c00000000400040004c4c40040104c000000300000100100000cf000000400000100000000c00c000c04000000000c00c00c000000000000c0000004040c00000c00000000000000000000000c000030100000040310000000000c000c0040cc00304c0c004000010000030000010001c30414000c0c00000400;
rom_uints[494] = 8192'hc1c3c0004040c00300c30000ccc0031033cc3000dc03cc000030030c350f000100410040350700304c0000431000030f03c0073c7c0304000033010030017c0410304030000d000d0100735000c0c0003100030c3d03033000047c0c400004cc013000c403003000400403c0d3c00040410000c050d000c000f04dc0c4100c0003f03700010f00003c0c0000030000310000010000cc1004d303000003000144300c0140040c431000000330005030c10010c0000000400f1044000f4f30440000f100000000470001c300c3c1c40c0cdf004510003110c0c31300113003000300c30071c04050000003000c00f0c010c034030c74c000000003034000000040cc03c00003c00331404c00000dc01000440c0000d30300000003000fc000c0c040077100000100c040c0003f13000700040000550c1000000c30404003000000c001c0140041000003030044cc000301c3004d13c34434c041c07004041c0000cf4000000000c0404f010100030000000100470104007000004d0410c000000cd0c00540004003000411000c0405000400400701000003c100040c3f010000c303450ccc40c000510003010000000450000000714103000041000000c000c000400000403340303c300001400131000345c00130004d00f0c000450001401330c000000000030c33010071cc1103c007c000311000000300400f0410c043c340cd100333c00c10000000030c000c400030544c0313000300ccd0f0300c0004c001c0000303cc00004103100010010100303000c0c0013c0040030000300001f140433001170001010001c00500cd00000f010000d0400c00003000d000010300f000040c3c00000000010014000010000100303000c0c00003cf110014c04145000114c00c000101c004007130c0400000401010d04000000040c400c4000c030005100031014040f303000400c300003000010c10fc0c004c30000003030f03cf0130300000100000140300304000410000c040d7cc50331000c01113cf3141000001005c0330040051404cc3c30003033440f000000000c0714030001003000030700334010cc30000c043000cc4f000000300cc3000000043300000c00c13401140144d400c000301300040001000c0000c0040fc01300005000003004100c00005d000c35011c000300c0400c100d0000140c10c03000040030003c00cc1df0c00ccc0010141334000304300770100301000000c00710c4740000000cc033041d53000000100700000000003c301403c74fc4d307000400053004300000c3010450c010170300000c443400c00c0004010003c0000000310f00000ccd00000cc300100044fc00050004d310c000030c014000013015150c3c03000cd004041c3400000410004c40030100300003000400040000000401000001131000000;
rom_uints[495] = 8192'h1000100003010dc000030005000c30000000001cd00040000000030030010040044033c00d00000340c00c00100c0d0001100030000010000000300030300004003000000103040040003d104000c033c3004030150301010000cc300014300001100370003c0c0000c304003f0c001404000300000001000cf03c0003000134300030030030000100111033530400c0304040000004030c3130000c3007f000304300c00001300030c010001f000d013004300000f4c30c000033cf000000411003000000000c0000330003300f0ccc0f00300000305430333cc00000000333303000c0003000000010cc000c050000010cc110c000003000000101000001303000100030c110003f000030c003c0000441100d0041400404100030010c0c10403f00000000000001400301010f01300000000014c10000000000000000003c3010d10004103000000000c0010700004000143f301f041140135f0300f000033450410030000100100000000443301013c0c0010030100c0330700401033000311070cc303030310001000c01007000000000c100000031040310c1004000301c70000000c10000000000000301130c00001103f1303100100000000cf4000053c0000305100003001000004100300540303011c13000000000300300c003dc000d03003c3000140401340000f00400c00c0d40310000030000000103000400400fc001c000003001300c00000034f00cc0100d0000013010341010330c00001303001001000130000c0000100d0000003000001c40f0040000334040003151000004c00100100000f03433031000010000000004000000054d1101331005307400300100303000003003c300100cc100f000c0010c3010040101001c03c00130d000003001000500c0330300050000703301000004530000000c01404c0d0000c700040030401303007033043c00f54003104303100431c103000041001004014000f00000010000000110003c003003004330040330301000000003c00030c00000031c0400000c0000101400001c3003003300400000140c000c34000030c040010300000070d00003300c0000013430000000300000000000333010301711f30501000000000300c0300c300000c0c30f00000000301004000100001c340c00000040000003c03010300c3c0003c33f00004010000371c00000004143400000030050000000100000000300100000301000010010d3110000000c01000010030c00000030000c00003100000040000013400cc3c00000000000cd0100f000010000c0000f003000003000c3c000c0000001100430c400340000000c0033101000c0013033c0000c0400005c00047003000000fd000000000000003000f0c00000000300000010000c000000f000300005000000100000c000000000000;
rom_uints[496] = 8192'h14000c00104400140c4300000c00000005cc171d003310f000003000301040000030000d004000c00000001000103c04340003340c0100001403000014c0010000c33f010000c017010000150100f7000c000000001440000000c0f01100c000000d0130c101030c070c030030403c000c03f0010c4c0003000410000000fc004530330000c30000104000cf03000c10041500000004300000310c04c40c0033d034cc100000c400004540000100000d000c1000001100c01001000300c3040000f000000000000405040401c400013400c0c044110300c010000430c0d431003cc0000101c4110034300000504000000004f30010c040000400004000000004c13000104cc00500030000f0433070c000c4c0c0140001c0dfc00030450c3000c5c34f00300000400005cc04000004041404cc0000c00000000104003040f000300000300c410300711c001700570404000f5300313000300010c0010440000000004330c031f0443030c014c3140000014c0100c357cc030c3d01004004000000310c5000030000440031040010400f0013000c00c040c0c0000c04c100103c10400cc030000000040000000300405400c4300c01440000030c0003c4004041c05403130c0c003c0ff00000c400d140c4300c04000000fc001c1300f0d0044c0500041c0000c005cf4c110c005000044d0000053c00404000c00100d1d70400c00000c0001c0d0331040300000041c4300c1001dc0004000c04003cc40040c400001003070c00030000001030000000003004000030c003000000c03c0004cd040dc00301040000004000c4013d3c101400013c0000000000c17000000000310c00c500f034c007000000000c03000c140100c0033c14301c5401400000d000000300100000003301004103030014c040f03054400c040004dccc007000000004400000cc00c34fc0c0300300cc0004cd0c0c00013c0c000007100014010003410000f010000c000f00000000301100003c03100c00040010000f0c07000c003c0000110000100d01400400075010c00000043f0c0000003c0037003c00101000000140300030c003000d05000c304000c00300000011040f0000c4333100007c044000000030300f000000c00c000100000044047000004050c00c001c40c30d030c0000004000040071000cc0cc404000c0c10014c0c00041000000c040001001011430c400c3000000c30c00300000c40000000c0000104300005d0004000500000301000104dc101500030000c00003000330010c00c40044d00300000c004400c045000000004040100700003300f504001100030000040c00300100c044fcc3013001f0031040403104000031c4c040100000cc000110440c00c0000c30c0040004404000000404c0001010400c000000300334043010000d30040c00;
rom_uints[497] = 8192'hc053f30000001010000c0000100000003000c0730000f0c303110440003000030300000000000003034430300330f307303001d04000001130000303404000c00100004f0000c001000000f00000000500c150c10d0340c1000c3011401c03c0f3030010c303000040030003000300001313c0c0c3c00001000314c3f300131f07c000500c01401000d100100101c4000cc004030000000300430cc000034100001041340000030040010d03000300311051103300c40000040300c00300401001d3000000005303000c001013010100004443f400d00000340011051c04000001c040c00001700003030100070410c0300300c10000010000000c00170000000101010000003103401401000300040000000117000040f404411013c50003300011c00031c000f000000000d00051c00d330005c04010000400500300c00c3000c10101c000c00000330311d4c000040300000307113000cd01313000000c3c303301007f0703034301700000175000000431140000001030c030033f0030000010d0c1cc10c00dc0c50000c1001001030000100100f100f0c001010100f3000353000300000000c00303301304c00040300f1004c00c0030f0100030100301043400000c3030000001300010000030cd1000c01050000cf0004040d047030310010070cf000033000733c3000300c001030030730001c001000030031c0f0303000304c00110000c00401010c07301c0000000f00cc01d000031311003400d30130030040171c00001c100c0c10500505011000000000cf00c04000400c01000000dc1030303000000431cd11033304141c400c100700101cc00c003104304000000031400000041000d013003001f10300300c000101000c0400000c003000f4405c0000030010300030003c0f100c101743103705104003410000003d00443030301000001010400300300000c3730010000770003d0000070c333001013c010004004003000471000c100c1004100400030400040430040c3d0101140033000000031c3000000411100f0000000000013c01000c100001103000c000000101050f100313001000030000040c3001300000000000400c00000000130030113044000430040403300c104400010000133000101c00000005000c3310004000100c1000001453000c1000000d00100f0000340000100000007430000033c040100000043400000000030000000000d00d0010cc300304013304001000304000c0010c000004040000433700100010034d03007003040000300c10000c3010030000001310103c000000000401000cf004301f0c100100000c100000000c03000c1110030100300000140030401000000030300400000c5f0c01c0303001000440500000401c0c000c5031404400003c000000000c0c340000050003300c000;
rom_uints[498] = 8192'hf04000c000004400c0400000f00000000100005400000c00c014d0100c400000001000c01054cc400c5000c0c00100c3005134405000040040c00000001030c000c003400050000000001ccc3000c3030004701103c00c00f0cc0c000040c001c0005c00c00001334000c0003000d04000000000001010c0c0300040444c00c00c3005c0140c0040000cc0300400500000100400000cc340410004cc0000400041100300c03c030040004400c04040400000300000000040100400001d0050004000404440000000000c0040c00030cc00c5040000d0000070c000c070c00000c0350000c000c04000000050004000400000330000c4000000010040c000000000c00000f00310100040f0433c000401c0400300c1c4c0f100403010d00ccc1000c0000033c0000100400010c1000433040000004000500040000c00c0c40300f3c00040030031c0f141001040c03000c0c04000c10000c00050000300400000000030043c0c0030c0c05000040c401004000c0000ccc04300ccc0003000014c00d0001100400000c001000d0370c0410400c0c00c0030000007100cc30c00003c54100040000000000000307000304040f0c03000c0f030141003700005c300c00c0c0010c0000340f104300000c0100030000030c00300c01000c0f4ccc011001000040010c01010d0d00cc010004040000cc03000c040c010f000004c00c04cc3010041c05cc00c00cc0d00c0c3003400403400000c304c00c40043000340c04004303cc050100000005034c011c04cc4030000c13040c4004410c400c04000004000f4001000c000000000100100fc0010400c34c0500cfc0000f01004f010100000000000d0001000103004004c13300010300070700000c030c400f0300040c010000000c301c0f00000c000dcc0cc0000000000c00c040000043330000c0c00004000f040303040f00030000d04c004300000000010c1400000004000c130c3004000000330c0c01000fcc0c00303c010000010c4403000000040430040000000503000100000000000c30400003043cc00401000c0c00000000000c0c0c0c0c050104000c000c00c001c0004400040000010004030c30f30044300c000410030c00000f0f0cc003000c00c000040c010f03000c0f00000c00000c10c004040c4d40c0030c0c1000054000cc400004c00014cc00000c05c004040300010f00c01000040400040004050003000140010004030f00cc0303040f00030000c0004000cc030c0c00c0040000045cc010c14c03050400073c00010700000c30100f051c01000d10c300003000c003300c0500cc000c000cc00300000000000500cc4d00000400400c000c000700000c004c400000010c00040ccc00000c000140000f03004c003000030c0f00051000410400000c0fc330cc0003000000000;
rom_uints[499] = 8192'h400c0040f04c7000c0100c0000000c4cc00c403000103010003c1c004010003404c40f45cc3c030040440000c00040f0001030301000f4c00030fdc510c0040100cc00c1003300300000400040000400c3100030d4c0330300c000c00000300c007ccc4000010040300cdc000c40cc00170000310444c0c001404030c05cd400cc003011000300170000c400740000c00c00440000c004000c400c400040100f40005407300c00000cc03c0c00c70030c0c0000000d0c040307000044730c130707001c0100c0c7035010040c400c10c3c4000400044c070c5000000047000004731c00003c00004400d00f07030c00100400d04000100c100000340c0440003cd44440434003310044430005044000dc10c14cd003c4c30d0cc0000400000d000c1000030000c0400cfcc033030c00441000030010034cc00c005004310c0007000004000001300cc330cc00144004403df40000cf00c00c000f300cc0cd3000000000074500014100000730f45010c3070f03504504000003c030010004c003000010040004000c000c0000400cc01c0000c040000030d00000404000005f0417d0000000003300001c0c300070401030000340000c0c040c00f10001044000000000010c40c0430c0c0000000cc10f40004c0c000c13100c3040000070101300030c00c4300cd0c000cc0010c3000ccf070fc00000cc3c07f00047c0000c140000c4401c00c30010dcd4f10f1c0c5001fcc3c03001344310cf040005c1041133fc403c5000500c00034000c0000c01c0300000c0c50c00c00033400c05417043301000d000400000000010cc40000c404cc00010004100000440c00c0304d00c00000f003003000000000f040d00034000c440c04c040d003404c503030017400c04010000704001000007004000344007070c43c001000070000ccd1403c0010001300041004307004fd1f0001cc0c1540f40000c0310400f140107c003f4000004007001c0000c00000001000300401dd0c10010000007c0040c030140000000544f0c000010004c00000c0004c00c0010f007c30004000c030333010001100304000040034c40000cc00030031ff010cc040030c0040110310400000c01035000c03000000034300c0004404c000407c4003c4040c00fc00310c055000c000d00003007c040000c3034400d00001c13000040340003000030040c000303400504c30c00004c30000c10c0040040c3c30003004c33000c0000003003c0010003410410004004c04100000040740c04c7004040004c00045003c00000000000000000004100440043100c004000400c1d01040000c000c00110001043cd0000074d000c01000044407000710000000030030004003003c0c0c1c00c310c0f004f100f40000cd5703404430000001000000000300c010d400400100c01000;
rom_uints[500] = 8192'hc000f03003003000034000000300f0400040000004c000c00000035340040004c045001c0000c30c0001010003003410300c10004311000733c03c00000000c003cc0000000003000100400030034c4000030100c0030c01c40100131710033043410000000007000001dcd030c1300000000000000fc030330004030043010cc3030043000000c00000000000400000000c00000300433000c00000400301030100000c3c0c03cc130040033000f0400000000000010cc40400130000004c00000000007f01314000011000114c000400f3003004104407410340400403000c4000c0030c0000050053000301c34000c411030c00410000c000000300700000044001c03000040440c4c0001000000f33030c0c070c430100004040c04d000c4300c4c34000000503d01104c04010c00030001c0400300004000d0000c3c0433070000c4c4000070c03c10010304d40c43f00100304f34111310000fc0000d00fcc003000d30c0401f0001400f040c14c0300000404004c017040010300d0c43300d3333f00c14330400044c00ff000ccc0c00014003004030cc000c43004044405300303c0000043c0000d3003440010003c0000401400cc04010041000c330003300300c0004c000003407c0033d11000c03303c000000310340001703044cf4000c004334c1340003000000d0c0004cc0001003131d30c001cd1110011010c0f44300440c00033d0003c000000004050350001140030004c043c300001011004c000c11000000000c0cf10004000100001c3000010044c0045004350004000001c3100035040c0cc00cc00004040c003004031000004c0033300031c041100cc3000004000030004300d0000040053c0c013330400f0cf0040003d00004005103001000000c30c0030c001000013f00340c31001c00c3000c1350ccc30f030133534100050d014c01500100cd144c0c0400000330c00f00f0401c10c00010000000000c030000001c00000000c10c30c31010040044003c00c000304040004cc03000000004034c5c3104000000104c031070003313cf04cc3d0000c13c00c53000000500400000f0000f001cc00c04034000000000003c4c0000401303300004001c0400004003f000c030000004001c03100100500007f0047c10040c00043c000f000311071000c0030c00031301000040c300000000000c0000c540001c1c034000011003c000c01c0c000403c73000fcc00c400000040404340f0000f00000031c000000c00000040c104100cd4c0000000f1005000050c0004140003003c1003000003000071c000c000dc03005000010040000000301c0000000040c1000c3010f030003c30140041000c40000003004031cc4303030404330c000400300300c000100000c0cc003013030c01000001400340000400004004;
rom_uints[501] = 8192'h33cc0000c7130400f0000030700000030400000000d0cccc000100034540500c041c0070c0000000107c00000c0f000c1001014c10c10000000c0000100c0330000003d00c10050c00000f000000440005c4000fc110c00000133000c30c000000000ccc01300700c11140000c0c043000333c33073c3c400070001100047c0cc00101130010003003000000dc00070c0030fc000030d431000040403030000f00d41000000c404003007000000d0c0004ccd400000400000c000014d0c0030c0310100c0000400107100000040f03000440030cc000004000c000c10403000c00300000000c0000040000500c100003c300133cc0700401300003000330037c00c0c030000004c0c33000f57000000040130140001f000034d0001001f004d0010c300c13111300010c34c40c0c00c31f0c0100300c0040044410c0310130fc3000031c004130003101001031340010100301c0013033c0c10c003004004c100c3101100c030c010d04040033c3c700000000000401305c007f000c00000c0050030001d0000000400000033c01710130033000000000003d3d0310000000035f10c10fd000010003014c000041cc00d10300304000100d0100300f0c01d00c001000104d3c0430301c30040040403c00100110130070100000001d44013c000070043003c03d1001000034000000130000001c4c000300c00c000c000430f000000c1030000c044c00401c110035414d03000c04010103000110703c17d0100004043001340f10010130144100d100041000000000000104004404000340dc0c0000030000c04100404c0070034000001000330c3030041004004c05c0004c1410004cf00c00c003300000000704c001001c34000003030710000010300c00050100007cc000c30373f0030000040c040301100c000010004d00007c101000010c00000000d010001001c00041004cf0c0000c10000300300c3173400000f44c00340000000000010d3c30040030cc043c70030c0010cd301101300010004000000c0c0430000000cc07c00c4000004c043303c0101403c010c04d007000010003000310040d0030040000040c00440c00010300000000d0f0d0030c00010030400c0334c000000030000010cc1000004010001000100400000fc03c10003053300cf0000c003000011000040d00304c00340c3400000000005030c330001000000004000001c074000001d0000000441d1010c03f000c0c303c000c0100171301400c00007300000000d1c400044000cc0c3c0f01c003c0000c05ccd030004003003740d10f004000045cc001330003404000000c3030000d00043040100314004f43000f100c0000000404dc400040010010000040fc3030003000301030000044300000cc0c041043014d40000c7000001000041510003c13100100000;
rom_uints[502] = 8192'hd0000040400d07004000004400cc000c000000000d4004003c300c00000c000c10030c17000404c451c10400030000400000000310040cc30c0c103000c00004000c000040014000000cc1010103000d10011341440c010000044004c01cc00000004010000003000c004700400400000430c000040c0010044ccf0040500000034400000000040010000c0000000000c0000001000000d4000004000000040c1c00000004c003c35000c000c000300000104000cc0030c010100500000045300c1c00400300030d00004c0c04500430c5040003700001c1050f0004300000c1310f000c03100c44001c0c130c4001000404410000000004030003000001000000000005010f000140304000431d00000c00c004d04004303040f041c3cd0000430001041c000c0c00071040000c0003c10003d40000040c0001c40c000000000040400070c0001000000040003000010340004040cc1cc00df0300410030100043000053ccc0c0f000400000c0440003c004100c04014c010cc0d000700034f4f5c000040c4140c00000000c04c100500c30c00000c003c4c044400c000003f0ccc40300c40010c0013010c0c00030d0c05000c00003041037301040c0001c40044004400030000000000d0040005004c100100000c0401c01ccd040c0300000000cc00001c0c001001000c104004410f31400000040004010d0d300c00000011000ccc0c0c4f000003000d340c4c410d0400000017001c01000c30004c00003f0c0105300030000340cf4c101010714c00000300013c00000000030d4040003d1003d1004001c0410004031001c1c3550000000000000000004c0304400ccd0000c040000007004000100c04044c01c010104040040004030100303c00001000430c10000c4d0031004c434070000c130d00430101000c000000010000430c0c17400c0001cd04cc00400140c0000d00007cc00010740103d4010001030c10000301000d0030300000030010c00000441470c100c1c010400c104400c00000010703000000c00040010700100000000c0730000100004040c0050000c00c4000000dcf000d40000004001300004430000100000c004c300003130c040c03450300000d43000003410c0c00000c00000043400000c00c0100dc0401030300c00c0100000400c000004d0000000c0000c4003c01cc04040004000000000c010f00000001000c0000040c003000000000404c00c4000cc505300100003d41000c0040c00000f00dc100c00404000c0dc04c0c1f03000000000004000c0000000000d1c403000c000c0031000000000c07c0004000000300000000000300c00000400c0c00007c0d100700404f300d31c1c1c30000000d0004f00c0c0000004000040000000c05700031000000300000d000054c000c0c00014c73cc00c4010;
rom_uints[503] = 8192'h304c00000c0c0000000c000030000004100c0c3440003c000014300000040004004c04d00c00000040c004000c003400043000f0000300040440000cc000100000404c0c0000000000000414d00003500010000ccc1c4c000c10030000c0000c0404cc301000300040100c001c00001c000000c00070c00c00d00440100c4c00533000047434000c0c0c1000100030c40000000000003001303004c0101c04000404340004300000001c0c003040cc00000430000000003004000004041c00000000000000000c0404000000000c1000040000300070000000440010040000000c000000f010000000000034104040000c00000000040000000000000c000000030400c4100cc0314c00040c0000000000003000c45000000000000730c000f404400c0000104c70000000140000dc0010000000001030040010000007100c4c00000000001000001f000c30000ccc0400c000430050010c0c0410000000000000000c1434c000000000000cc03000100400140000000c3000000004004004005c10cc00140000000f0004004400500c0000100000000c000c40000000000000107c04300000000000000000007c34000004007000100c10100c4cc00cc00405100000000000001300340000400010015340000004001f4f0c00000c4000040000040c0400000400000300300000000c40403c00f0001003d03c4400040440000500c0340000c40000040c0504300400101000000000000ccc00141010000000040c4c000c400040000040000c0c000000754c000010000c00400440040030440000000004000000041000000c404c000000000c004000340013400004047c10000400000c4c00300413100c00000c00c0000c100003000000000c00100cc00c041000300000c0000c3004004c04040000000400003030040cc00500000000400c0000100010003004037c0c0004000c3400000004030c0f0c000c0130040c0000c0300000000010000000001000000400140c0c0100c000004030400040110c0c000c0030000000001c0c041000000410040c0c000000000c0400c0740c000c300000003c00004c000000000030000c00040000000cc00c001000100c00004c01000000040c040040004000000000c4100c04000cf4f00000f000040414000400001c0054000004103c1400400000000000c000000100304cc0040040040000340004304034040c010000000004000000003c003000000c001c0000040000000000700000000c0040040000000030030400040c043001103010040010c00004c00f00001c001c0c0c0000000400040400d0040c000004000000000010041001001c0cc40000fc000000c00004300004700400040000041400c00c000c300010140cc00000c000cf04000000000004000000c000000040400c3044c000100030;
rom_uints[504] = 8192'h11c000cc30000c000000c0000000500030000330400000003d0030004000040c4400075040000c0000070300530313040100c01043010030001000304030000c0054000c310000550014c54300c314c0000044c0005cf0040000c000014001c00001304400100001c01400500400300010c0c0104c044c3104100300f0000150004001c0d0000030000400000010000f003030000010c000004030034017500c501003001000dc0000710004c00301000f0001000103405000000030f00c31c1c00c0030000c30030310004000001045cc00cd0001007014400f00f000040c0400c03013001000fc1040074140100103010034400400000400107013000000d000000014001c0013003c0034001030001d000000410000c00000113010003004dc1000d01000f00300000000f03000c030c000030000000000100c00400003443c00c030f3030000433003cc00f0c050030c5000130170500c0c331050010334d00d31030300000004cf0c0c401f5010300000c04001111403444c400c100071000500444040040100300070005000cc0000040000f0000000c010f05010043041c010cf30400d00103400000c331000340c031034543c1100c00000100031c0014c100004103000f00000510000c0cd001400c000d4000ccc000400100003c30400003300004c1000130c0050300c100c0c3000c000040303400400c0f0000c00000003c040000000004cc1000300304700c00300c0c0004004303000403003700c004003004000103000030000040000400030c40030401d00c0000000c5400030c0000000001c4010c00d3050c0100cc000c01c000c00050001000010cc540fcc005000000400000c0000cc004043000500cc0540000c0c00000c00c000040000004400c000403040030035f400c00750100000010c0004005410c3f00c400000040013003cc0004c00c104c03003003000000040000cf000040001c0004001030000000000cc000000000000003001014c0004000307000040503070100000300030cc0c0310035000c04c0c0400300003cc0c0000f0005f300000c0000c30000150f000f3100000000040c0000300001000001100fc501c50000313c0d30c000300000000c0300000000050000013004d00f40700003c40100000c0f00130c0100000004c004000041003050f300c031045003000d440310000010414c0c01050000c30c30011c05000000c3040340f3c3000f0c10050000000c0001c0c004100f030100000c0005300c0c0040301010400005300f030500013400004d0000c0030c710030000c1fccc000000001000330c00003010c00000000000100c4000c700000c00000000c0f4c0001004000f0c0050004010fd000051c0000000f05700000c00c14c00c700f10c50040d03c1400000001054f0100030000000;
rom_uints[505] = 8192'hc0400004000300000d00000003cc00007100070003030c0000000040001400300003000f040000000c0040cc00c0f0ccc3c040034003401c0000000c5040c10040dd0304007400005400c001100c0000304000004030000000000301000000d040070007700000300000c1000303010000000300000001000315f4c35004c0000100010c70c0004400040000440000000c14440000c00074cc010000c0000d00140034cc000c1c0c14000000400100550f30430000c1cf10100400004400000011c100403c3000c0cc13c00000101c0400054044343070001c0001000500033031c0000100310040000300c040041c04d034cf0000c0000000000cc300300000003100000c0c0030400000c0440000000043000c005143003010300000cc0c30010c7000330c0003400c0001c030400c0003000007000c0000c10300370000401c30040030fcc00040000c3cd0005c3000000000c311c0c30030000d40074000000c03004d050f054003030000354000000000071004f00010c00d03040000001f0040c0f30434001003000040000000003000c0000004000100000000040c00100000000000004400000000003c0000300003010400c00007c0004010104140055010000100030c00cd000c0301010c1f0144000005000c003001000001000000000001c007c00cc0001110000400131c0003000101000030003cc0c0401cc0304c1cc400010044c0c10f00010c000100000000f40cc00070030030004040c3000f4700000f0070000041100340044100c0c000010c000f0104003cc100c00c000100010300000003c10010070000000000d040004c7010000100130100000f000d0000040010c00004f000003000000300c3400004c003004403000000404c4040c1000000000000000300010000c0411003c01cf0005d40c00000004030000c3403073c41000001000c0c003dc0513c00050c00430000001040c3011000c00300c100440000c00c4000740c4001003f441c400010d0c0cf0c00f01c03044100000300330c01c0c03000010010000007010000000400000300000140040c00c000c000434003d000cc0000000003000c00cc0d140401004001300c3404001370100000014000000007031c00c0400c00cd0400000c0000cfc10010000c30000c0004c00000010000007c0044034d00000000070004000001000000070ccc00cf0c40000c0c4000c0000c0300004400c0c03c03d0414c1d4ccc010004c0001c50c1c0400c034d10000403d0030c0010ccc004033f10400c040400c1000000f04000010304000000040000004000000000000040d100fc0c00101000013400004404f0cc3000004000000030004700000c0c400000c730c000c0100100c01c010000000010440004000404000c44c4000001000000010c0c00041c1000140000;
rom_uints[506] = 8192'hc000040c00c00000301c000000030030f0c4004cc00000430001000dc00d0001000c0440000044000007dcc0000c00010c0c43f00c0000000001c1000105000cc01010004c0f04000f0000f00c00f000c00010743c3300300d0000000001000000c004f01c00c0c4400000c0010d40010000000040c0c4c00c0030000000c00000c0000400003cc0003000040030001000301300000001040c000cc30000000070000004000000000400001040c0000cc000400c00040c000100440c00c000001040003c00300000c0c0c07c00130c00003c00cc03003f03c0303cc0000054440000003000c0010c000c400c00c00030000c00000410c0000070000000140d1310c000040001f0cc000004cc0000010c0c001c0100400000040705030000101c000400040c3c03000000400010000000000010000040000400000c040f0c30c00400040130105300f00000000000cc1100c00c000c00000030c000c00c30fc100400003c00400d400c40000400100000300c04344d0c0440cc0301c0015ccd00010c0400c0040100f44c0300f0000000041c040cd40004110000f00103000040501000000000f0040400f04300000030c0001150f000000cc0100c04300c300000ccc04400000000000000fc0c004040010000043010000400c40400c4070010000141440000100100cc07000013004050040000000000300c003000004cc04cc000044000030c40000cfc000030100f0000c0000c0c00c00c0004f0003c04c000c10000030010000c01000c000000c000000c000404300000c4440400100100004c0047040003c000cc400050c0000004500cc1000000c0010c304000000c0040100000000000304030c540f040c03c00c000400110f0004301013000500c000400000ccc0030100300003c05500400400400000100f1c4c0000404000400000c0030f0c43000400031004000000000c1004000d11001000300000004000000000000000010000c000c044c0c5500c7070cccc0000000000000000004000c00010100040140000000f0040004f0000000000300014003000000000040004c000040003000c000ccc000000000000100000000000c300c04c4003c43000040000c0000373c004c40100000c0300c0004040c30004c004040034000dc0414c1000010040c04f00000000000003000f00400400140000000c00000440700410040000c0000000000100c400c3c5cc0000f00000001000000030c403000010c00000000401300000c40000007304cc000304000c4c0c040c300003000044000000400000040003000043000000510f004000005000c00000000000000003c000d0033000400c3041cc00000000040c000000000000004031c000130000301001c0100d00c040000000351010000000000400c000040000040000000;
rom_uints[507] = 8192'h34433000c0c0c04103034000030000cc0f4c00c0c000100000f000d0001ccc000070f34030cc003000141c00c000f40400400430410c400d50000c10500100300003733c10070000130000c5130074f0013f000c0c41000034404000c0410c0000d00000f400170133007400300007c000030000000c00c300170357004c30035030c0000c070040000c0040300000000000c000000044000c000c00cc00d4f000337c00c050000000c01c015500000000000004001003d00034004304400030030000c00c000c030d400100010441300004f013040010000340010c70c530300031000030c00c00003c100000c4000300040c00053d0000c000013d300300c0040000100000d0010c0701405030005110c30033030030c043000343041c0040030403000c0d0000000c00003c0c437c703c10100304cc0014003d00f31300030c0c00130001300000101c0010007000100c113000310c50c00101040000c040530cd03003440c43000d10d34004500001c011c00303004003cc041c110030100d000001105c1000000300100010001001000ccc0000000030340050000000c0500f00414301000000300cc0c0050f00001140c3f40030c0400c304000003400001001707033007400403000cc00d101c340cc001110374100c0c10004300cc11030c004c0000010050c10003c3134403100c003040400300517300305003010000003000300100030104304313c0440350c000300700003030001110040715000c30030c0cc000000000400700003700101400004000330300703010430004013d050143f40000003000033003d73c00130f430413301104000000c00c0003c03043033c0f0040110037013d0000003c10f400c3c30040c001300303330c000003300003c0010403c433f0001000334007cc001040340400003030031730c30cc0c000d400300000000c0c0c0c03004f05f000f0000001000030cc40000d0000010003403003005043cc010304fc331003000000004000300410300010c000c0f001041c10000cc00000041013c0001403000c37310110000f40404000003000110c0c03301037c001000d000c30300c404d040000000000050404004cf3000f0c000030000c04000cc000c0103000c00047011303400010cc0040f1040010400401c000030d10c000d000000000000f003c001000000473300000133c00d0013cc000300100010c4000010000000c4003401400050c0c40cc0c00000003500100dfd4d003004c0d0101c430333000050c00031134740303f33cc101f041030300c41c3d00100c100014400004000c000400033400034000000400000c3d00d1430fd01001433300c00d0300040004000007010005dc1cc0303c04003044000c51000000000c00300d0300030c31130073001003cfc004c1c00c31f3d130c00;
rom_uints[508] = 8192'hc00000dd00003300330030d000045cc00000705c1c13010301500000c304c0115000740070030400d0104010cc0dcc014cc0030100c000000010d030010030101004010c0000000000441430404c1003000c0703f3500d000c0c0440d000000033f0003c3c303c0f030040000730c00100400c70303330c4010000300000c7004cc010104001c00400000cc0004030000104400040c0ff0400c00000001100000141f0004001110010c40050d00f100340000000007cc00441001053300700003c30000000000040d0c0005c1300100c4451c43c13000c0fc0100010c431000100c000000010300c4017c00c0040d0c1d1c07041000000410c0400400000030010f000cc0140400001400d51401030d0f00301000010007000c10030001474030f0000010030d00400c1307030305d05c0c0d030000000000010c00c100000000cdd000470400030c003300030400000d00d004051c00c3003100010000d3000c00101c0011100001c010034d0c0001010004010701030d03400dcc00140c00000100150dc010000c5c0c0103000cc300030104000340035d00c00d03000c0dc431443000c00c10040c00041001cd4404000501040000c400000000c1040c400d0400401000071f30000040040000c00111c0000c0c0000040110011101d41c000005c500c00c3404c73003003f013c40c001010f070330005000510cf500010404100030000044043d030014010c035004040f00040003c0040f0c004000051004c50f43000000043c0400cc000300040d000304040c0400540c4300c0000c0003001400cc0c040d00003150101c0fd501000d050030c0500010c0400c040030004037c0cc0000000c1c0c0000001300011103000c03011c0c000c071c10450c30070001c0c013c007c07100400030000d1000330043000000000044500004000137d500c3c307000ccc0304c40c440040000001000c0c0c0f470c0440000100310010000400c3003c4404c00c010101300c0cc00c00c00001010c050400100003c1013003130141400f0f0000000cc0330f000300030c050d0c40710c031100311000c00003fc00070c00000003300100001c00003100440000000c0400040100053c01cc0c100030010400010000f0c7030010010004c03f0d03000303c00f01040000413c4004c510451030000100003000400000040c3000c34300010c04400c010d00000000131c30c014030404000500c40104010400040001c0300000105000000c00c40000f0000d1f4700000c000c1cc0000f13310010000014c0010f0c3c04000040cc1140000cc00c00003030470414c0000001000000c000003714000315dd140000300147040c04400000000c000004c1030c04010ccc01000c000013c00c000071000c077cc013003300005cc0500111cc140514000000;
rom_uints[509] = 8192'h47000000004000003c0000300c000cd0030c00f0000400300370170340000040c000c0030c000000010000c0000001c0005000cf3141003fc0170000000104000000500101000000c30044c007001c40000700c0f00000c001414730007001c3300c00000100c044033103000004f030011003c0005400c0030000c000c000000fc041000040000000000000400000000000003000000040cc0100000031300000400000c003c00cc100000100f00100c000700300000030103003044000c000c400c00100c00334030000300040c00100003000000041c0004000303030000300c00001fc000000c000010410000000005410100000000000000000100400c00045000005c001000074310047011000c0c00100000044000cc3441c0410c10004000c0010000030000000030c00c0404100000cc000000003c040d010000010000034000030011000c000c30003c0040013001140503010010003701010004003c030000400010000000303003440c0000000000103400010030001410040c04300004050505000003000fd3401d000300000000100000003003003000003c004013043010001000c10000040034440700001030c00010010300000c030c000c00300c0000000c030000c00d000c0035c00000000005d0003c0000000c0000d004000cc0100310000030140301004001f00030100001003010071000070007c03003c0100330010000100004130c0000000c303c0030101700001000300000100cc000310d00000000003005003000030710000d0000000031300003400041d01c004000000000000f00000004110004100c00341c10c0300010000000003d0010000c3001010014103000030404400c0000300001000403100c4000010000c0440000001000100c03000300100f4000471d010c00701000001001000c0000001001150001101000057c1cdc040c0c0100000d0000011000000c000400000030000310000000003c33001000000000001003cf01111000100410301c0300c10000000007000000000000000000100004000030000000000000100000100000040000d140103000c000000f00000000300010000c50300030000000040c000d03030000000000010000000000100500000c0703003f30000c0f0301000400000c0400010d00003000000000003003000003000f0303d003000000300000c03d0000004c1000c30010000030003401000000000411003c0c3c000000000010000f0000c00c000030001040100034040c0000047511dc30400034010000000040010c00003c003004000400000000000030000c0013000000cc000000000000010c0c0410313c000f00030c4000005000004c00000005000400000f0c310403033c00000004140000f50000044c0c01000300000c01010c0000000000000003000;
rom_uints[510] = 8192'h4001004000000c100400c00540000c00003001300c0040000c030000c33304000010310010c0000001300034000ccc430000043c3003010030c300c3c0000000000010c000104300000c503cc000400c0c04000003d0c0000030030000045040350033400000f100c0100014c1030440d43000c3110013000c000041d0c000001000c000003000d00010000f00000c4cc010031000003030040c0040400000100100f00000004000c00c40004001004003c000000c001040040000330310000040c0c01000000030104010c0004c40000400301000301030403c0cc0f17400030030000040c010c010010034401403c003044410130000f030004000c0c00000c04000c000301000100700c50070c407c3403303043c43c0f1c0c0010400050400c0000000500040003000d3f00010400000cc000c0030000000300400000c00300c40104430000300000330c051c00c101c4c00c4d00004000010c000000c100400330040100310000003400030300c410fc30f4000d044f0c0cc00000000134144300300d0000f3c001000000403003000d00400000c0000cc001040c100050c007cc030d0c01000470000004000000001040ccc0000035000c00070c00004015c103000c3001004c0c0073000004040c4700fc33030404130000301000110d0c0450003c00000000001400d00030000400001c00f0310004030004030f0d070c000c00c00d00030700040fcc003300040743013400c10010c0000f0d0004000340100000000400000d000000c003003c0c0000cc000c3100000f4c00fc330400c411403c003004c0c0004c00043000c00c0004030d000c700000005f011300cf00003d0100340300010000000c0c1000403000470411c041040410000c403030cc0030c01431040c3dc4400400007c0314010000000000003404104c3400000c003d134007007d470c7cc010041c310c40c000040147dc04cf000340114c040110400c00003000100c0000c0ccc0000000cc30401f0f1004003d0403c00c000000001f00000000c04005c5140014300fc0c00001000400c00c103f1c0001c54c01c030c100300c14000c00003c003c03c0000401c000c0400030f0dc001003000c04370c00030c00000703c000000000c301c400000000030fc414c3cc0c000000000000000301301d30c003000c0c0c00300043000c4c000000041330000000c00c040c000c00300007c0cc31000001c0300034030447000c00000000401500000040000000440c0dc4cf030c40010530074000ff1c004033c3000c0100003035300004c0c3310004033500000400104700450003d0000000000c0c070c0100cf01007030335000d00070d0000000000c1000c00034000440007000000400300000cc0c00f0310c3000407c0400000c0000407044300033000337000000;
rom_uints[511] = 8192'hfc010004c00740000c0000c0105000ccfc4050304cc44000500430403fc0000030d0d40111004030110cc104f03cd0c001300f0c40f170c0040013c000d000000030cc03004004030050050000c0400104c3c054004303001000033000000040034004c0c1300ff000c00cc0000c10f00030c07c0000f300cfdc435c000000c00040c0c4300030000000c300004c00c70100000010c3c043c0c0d4c70c10c00c4c010500c0300030c00341d0454010304fc01400440000400c0000300cd000005c0c10dc004000d000001c0110d0004fd00300d000c3000030c013cc140c0100d1c1400140c10c013000f000130c004f74300041140000030140400070000c000130003531c0c030d00000c00001c0d04005c040300330004400c45307c010000000003014c070003030703c0000c0014100c34c00700030000040c0c3103030c40000c010c0c03c0030700330c000dc31453050f00307711004f000000d003000c3107100c0f0c0c004310000105c00d040c4003cc07030d0ddc0000c4340000000415300704013040030cc00c0d0c100c7f00000c0000410004fc0d00000000cfc0073c0000700f400003000c01330c007f0100040c41403000041c0100001c41441c041041100cc003071000004304c0570c7c0330c3040c41100c0c0c0c00003c10003001f00c40300c045000c70c0c000000100100140fc40000000f300c00040c0cc003000dcc00410ccc1c0130005f041c0010000001cdcc0101013d14c0000007300300110c050000300ccc0130000104044f0007000111500300000c010300d30f100d0c00030033030c4c0c00000f4f0cc401071000010c070c4cc4000307040703003040cf10cc104cc400000c0c01000c0d0c00000c00c0010010710100c4000033c00c7c510ccd04030043c401000300000c00c100fc0c000d0000c400cf10000404c00c0d30f00103010003000300f4030c04c14030000000c003000c000301013000040100cc0c4c0440000cccc410410303030773c0041000000300000010000f40c040040000004d0c003100070430010400000c0340004c000c0c1c33004c400010000300313cc4000f00070110410c074d0105cc010d0c4004cc010c0c004d04007301440700000314430c00000101041330103c404017401003c4070000030d0000100130003ccc0c00044c0300c1040003c0c000d0000000c7c304000001040001010d340d000040040f0003100c0004f3013130010440c00000c3000f400100404100051c310100000c0000030000000d0400001044004715040d3d5c0f301c1c0c0007300d040cc700000503000000010004440100000d10130f000300040d0505c500001443054003300c0014003007000004f04100c30c400000cd004300010c074d00041004c00f010c003f440c000303000;
rom_uints[512] = 8192'h30100031414040001000500410004c001030040000cc301033c0100003f0c0004140d0304c3000c000400cc0c0c00003040031c07000141040000040f3c04000c0c0004070030d701000314c3030c40040c00333001030c3101371f040c5003035101030003cc4c0c0000004d0711040d170d01410cc00111f31701001500030100c003103c0300000000000d000c0c0c0000f000f00f403314c0000505401c0c0c0c40003d5d0000c7000f04ff000c3007300700010013000000030f4400033704007401003403174c00473cc30c330c000c35400001c4000000000d0400040cc30100000310000003043f03010c04ff0333300d5400000c0400044c03015530c414000701000014051400030fc0040c4300040c4c000540cdc40c0f330f0001003000000c0c4303c400140303301030040054303c0400100007503033000c0701c70000c70300010c0305c00000030c0100003d0c074150403c44050354c0300fc001100d303f10450cc0000000c4000404000c0055010041414c0c0c100000014c04cc400004043c0004010153000c00100700010f01073c400f07c4ff05073f03440100003104c00c000c0c030c0004010f0703010300000c0003000d0004010c000140ff050d0001007704010cc1030000000030300001000c00cf0100010007000340c40004345c00c0000001cd030301010000c444030c0340c0040043000003c100005c0313010c10c1c3c5c10004c3443007443401f401055101300cc00003001f000f000007001500cc003340c40301040c01030f300f0104130444100035030c01003003303c050ccc03030137c1343fc33104133040540c50000df4000c011f010f31000400010001013f103c13cc0cc000030000000000034c0031c0000303005c0d30000013000703034500070400005d0000150700300cc033fc00010010000c0403003f34000307410d3043503c000017f033c040070400cf0040000100000400400cf040110cc3004c015113313f40030000000003004710000000430453cf04d00410071f130f04005d400d0330104544400101010c0cc00104cff001c4040f04500340fc50300101f10c00000100044d00504000c4031f450000034000040c07cf0400c30c0003c00c0104c00000070310f0043404430f0f050400700c0100000d0c050f4400413d0700cc040c1f0c44300cc040330004001001034000ffc1010000fd0000400000c003075000040fcc01010ccc353011001f00304c4000c001000c1007c0104017c00c50010f000044c70003fc000300000001c0003401000f040fcf030c10003041043000010350000c00000c0030000f540cc73f0d30005100000cc0001d00410000000f00300000030047000c000000401003c010300403040051030000f005000000034c01c000014c03cc0c30;
rom_uints[513] = 8192'h103300000d001500000cf1c1000405004030cc500034f0010c00004f540010000c0c00c14000c004d00d01f00003c01400000c000043000000c1000000700010f00c000000c04000000004400100000c003004c033030400c300000400c040030c011d0c00301010003c00c400000000314d300c00044c0d40500d157000400433300003c0500030300030c1000033c1030100000041cc000000001010c000300c0000c000d04c000010c01400013000000000000000101303300300000000ccc0110c0001000043300d5f040c003000f0c370000110cd003040cc0030010004700030000000000013030f0c3304430000500100003010100000041000051000004004040f000400000c303d40004cc400410030004403000004401300f0000733300043400c400f400d005010000000000000000000001000010000000000c300044c0c100d0010c0000000457000c00c0000000040000f5cc4300430cd00000c4317411c0004003003004003040000044000c1000f100c0c00000000004000011447c10440100f0044000c00f700c00c10c01000c001c03070040c04044f0c431034000003f0005000c0040010000000330400c4c0000000d050004c00c1000c403400000c003c407000d000f00c5000d0040001301003f0130010f00c33030cc0000304004000c4400050003000f0037335c0c0503f0c30000c00003c1c00000000000c001c0000130004704040041c00003000041100054000014c301000300000107007c00c00d0000000001000341c00000000f00c00000000040000004004040303c000140000f0c0c0041000d0c0000000000c0c10104010100010301000000004001400c500300004000f1001103000f1004030701c0000300c500c1c00c00100000405c0000c4003340c00040000000040300004030430f3000010110c0c00c4001d000c03c5103005000f000000c00c300000c03030010000033007c0000000000c41d0003c040001000031c7fc1c10040c00130c0300410410000000f0310c0c0000030c0300004c31000c370103000c0d04300c300500000053070f1c03300c000000c3f0040011f300f003007000000010040c5010007c10070000c050005000000000000c400010c043c3400031000f10403000000040040f1400000000000000403001000400103c00050cd0000000f0500000000000001041001c0000003000003004c00000cf0070000104000043c00000cc001c1c03001000400d0dc00010000307104044001004030040c0100f001000045030000c003c14003000000030001004d0c0000004fc000c5000f00000403000010030c00c004c300f00000000033000034440400030001000001100fd00001dd001c30100000301100140300400c00cc47400000000040000c31000004c004050c0000;
rom_uints[514] = 8192'h10000000100c0c000700000cc0003d35700003cc3040d500000040c400000000c300003000c0010000100030304030007c3030400000c0d05f000450701140000c7030000c00c0d0000000030000c300d4c00004c04c303000113300010000000f001010100314100000000040041c303030c10c010414000400010043340043d001d0c010300000000000001000001100400c000043340400104000303300403100000401c0010030c000c0003030300c045000003004704010003c407000004110000000000030140000c001c430303c044010141000401c31000000000000700000c1c4001400007003cf3c00033403030c304010040034130f000000003050100000000c4011300000015f7000010000103000000000c0c00010503000c010310000130c41100c000040004400c00c00000000000000c0000100100c40003000004000443000000030010030ccc450300c3100510c0300c000c030f0105000300004d031c00000140070005000740040004400c050000300c000c001000dc100c30300000010440030000000c4010000f000100f010003000007003000000cc400010c000010000c0010001400004410c04c0c44400d404cc00c000400c04c00004400d0001000000000c0013c01300003f4045403c000004044c40c301000300c30c0400400cc010000f011433f300c300040000000000400001c003040c000000000d001cc05100300c0d00400c000017300050310000040100010c1000c00d004140000c00004c030000040004447000000100070c033400030040cc0004053100040000050540400000cc0c0c010c0000001c0110370000004c47440140004030004001c00c0000004000100000df001030470c0c0000000340030000001000400000000043073030000340400133040430003001c04110410c100f010c000c0100310c0c304410c10d040301000030340fc0040003030001000c030000010c0000040000100300010d000000c000d3000040401340334f043f000045000000300c0100000400c0300c000300030d3300310000101c101001000000310314033c0400014100041001000700100d000000004010040cc41d000031414c730100000104000440f0010c004f000000c0040030400005000c3c1134004100010c410000170000c04100003001c10c300000310c00450cc30400030433100d00f00c3c0c00000000000033000000dc0c010003001cc0dc330000040304040000010f00000d030403007004300040010c00050004000003030f10000300001310003d4f0000010c0000030040010c004c0003c4000c0007040000001c0000000300f100034ccc0010030000c3000d000c000c0030000100040000100300700000400010c400040c00004003033c000000033300c0cc000040035c3c040000;
rom_uints[515] = 8192'h1d1000040040c4d01003000100c1003c030000003100f00000c0030010c000000003000000011004301030c101f03ddc50001000000050c000c00c000001000011c000000c31003030040340000500000100000d0010c0000c140000000003440c510c10300014000010000300cc030f00400004433c03c00c0c0100130300414100f000000003500001000c0000000000c00100000040501c000403c01043f04501000000040040000c0001000f01f1030300000001c0c00c0000000300c000001c0c000c0540100040010011000430cf000040000c0001c0013f0c130000000000000004010010000001400401000fc4c0c4070c0101000041471300000c11010f030017004c30000000000403003011430410014c10001c300c40c1c00000000040000300103300c700400303040c133c00000000000001000040401000f30000005000c00000c30004500001500c10000400f00d0043400df00000405c0100033f0cc0c300171300000000000000010c003400c030000ff0d450000000043d0c4000040000400c10000403001c014000000040030003c0040010000000000c030000401400c00c040000c0310001001005007000030c3000000001c100074c003400030430100000300400000c01000c0000130100000010000101040043000300000c03c0000130000c4f000300371000000000030030f000004030040d000d031c01040501030000f01c30040c0343400001110310000040400000c00d000500030fc0000030300000c0000000034400000000004403300000300004000100400010000040140013000030000000000c3000c100040403100f4001cc000000000310001010000c0003410000001110c0000307d0000044004000110c000000000000040300001033104cc1c30c0353330003100c00000c1000000000000c00440c304c0300000f070c0000001c00d3003000000000300700001030000031c03400000000030011003000000403000400101004104000c010000040100c000000010000000000001000403000300000c0f0c000c0040070000c000000000400100d407000300c00000000c0000100000030400000c3001300430000401430000100103000000011043000000c50000cfcf3001010070d4000400307003000c033000000c000010000004100100000004401130003100050000c01000c300c000350c030003df000000c10000000340004040304000003000000c1100000070c300000000001c000003c00000c4cc000c0003040f00000040044c0000000f00310c00033000000010110151000000507340010000400001300010104000044000040040c00300000004300000000000000000010030000c0000040000000000007010c3000d01000040001031001000070000004141000030f401000000;
rom_uints[516] = 8192'hc330000c10001014f000003d041ccf1f3004cc40cc0000300400c00c0d304010c0030300004000d400100307400400f3010004003c3c0c4007001000300c40300f0004c30104010c000c0c0f400730400c0000003f3f071c10434c70000f00c404300c00c40040000004000400000c000c0c33f10c000c140c70cc0c004d7c07c1c3440c01300c70003004c0000000700c000400000030004c000004441c01400544040070f04004000c0000070003dc340c00000100c04d0cc00c4c01031004c00000c00c401c070c30030d001f041c0400400cc40000040040010000370000034000300000000c33400530050c0d3004d40c03144c0000004000010c000c000300004cd400300c7004413044000003007400f0000000c4000000f017030d000c1cc0040034c74440100040000035030c04034f003000004c04400c0c04cc141cc4dc0c000c0000440c0300000340cccd00003c05cff300440731c00c300c400003400000c0f304410c4fd000140400001cc4000c0010005000cf0004005004c1cccc340d3c70000d03030404000d4c30004c011000000c10000f00000000001417000000c511cc0f001000c000400430400010f00000430c00c450c30000c01000000000c0000004c0c00040000c03c4010000004c00c000000030f3031300c0f01000000c0c3c0dc00cc1c034c03cc000300000000030cc040000c4471001c07f00000f003c00040300010433c03130c044000c334000040300070000001000c05014cc300d000000040000001c0301044c000c44c11c071c040c00000c3c0000000000f010c0030003000011c003040410040c0f1c0145c010040c0f54040000043470000cdcc30c0c0c4041040404010040c137000001f540003300000c04003c0010070000cf40c1000007f00041cc1c0000c4c0000c003ccc03000d040300f0003d14000030070c000cc40cc0c5410cc000c0ccf010034f11030f004410c50040000000c00c1c0000010d040f0100340c40131c0430303440041c4d404000cc000c0103300500040c070c400c0c040c07c41c040700cc000540001000040c0ccc00c1134040010f40c030000010000030001030140c040c404010045440730c04040443005f00c01300c4003c10443f1000c04c04c410001c10cc40004f0cc30000c00d540cc00c01013ccd0c0c0000301404400330c0000f0d3c010004007743c0d0030c007007000c0010040004370c0450040c00040000053700103070300043000031000000035d33c40403000dc73000330f0c0000004c304c070cc400dc00c401000300cc000c04000004c10000d004000c0c043000c000000cc130003c07c0f030000404300cc00730cc03f0000f051c5000400c031f0734000dc000030031cf4c000c00440000000d303003001404000003404c010003000;
rom_uints[517] = 8192'hc100000110c000c401110000003d1000500c0000004010000014000030000440010770001d1000000000000400000310300034f00000c5c0033004507000000010300f00000c00000004ccc000000030134ccc030000c030c0c4c0000130000000300003700000330000c030c310331000c10031440040400d10333000010c0010040005000001000c044000400c000070040000004000037c100000400c0100044030cc0004040cc00ccc03400030001c00000000000000f34c004c003010033cc00000c00534000c0004100c0c000c500cc00347701000c1c07440c40000c000000000140d00000c000c4f01000c4c47c00c40300000500c0000c000000dc10003030c044c00100c01c0004000040300d4004c0404000f0c0001030c4000033000100c0044030c3040cc000300d300300050000040c000c0c03cc0004c3d0c30c0c410030c0000400cc0301005100c000c010001070401f3045f0030040010101170c03000000030000cccd003c004101007000cc7000001131440100000000000503c700100040030730300cc0cd4000000000000000c1cd4000c0c1004000340c4c3cc0003c00004000c04100c0c31c000c330400c000c40c40c004404f3f00744010300045400330000c00c130c010000c4003c000c030d3000c014110400003c303f30f1140c04104c0003001c000010c400000d400c00000f04001d0004f000fc04100c000c0010ccf040cc000c04c003300c700c4414040333410010000003c001101000000c144ccc3000040540c0100cf0340c13000000000d3307034000c000030000003000000c0c04400433c000000c100410f400000c000000040c000070000300003c0c5cc40c430c33004000000003040010000070040000043340010c00c00045000004400304303c0cc0000444c00000300005d003400f01004c000c104050000000c0d700fc07300400000c1307001050dd005000d001001c0000000c44740000000cc0000000000000c50c040c3f004000030c013001d000000c5000000c30c0100000000000000300030000000000000000fd130000c00000c00cf0c071000c0403000001c04700000c000300103033c510cc4000055c400c100000003041d0c00c3001003004100400310300000004c1040000c0c0034c003c300074c0000c04010014c1001000000303400400f0c004000100010c0000c14cd00c04c010000003300500000010c030000040cc00400000404c30000031c0f5000c0c000004000404000d04030003034004000700f3770107003010c030300c0044c00000100041c703000417d000d300000000000c000010d300400c1400300000440c1000000c0314000f04c00c4004c0040c0040040030cc0014c3004c0400300440dc0c3030c700300c700000400cf0c41007407c700000000;
rom_uints[518] = 8192'h5d0c003c001c01c00000c00000c05c1dcc00300000000000004c000c00fc000000110100dc0043c7000010010137c44c400000401c030401000301000011000007101c0000000c00001c00c0003f1000000003f00cd00400c000000000000103030ddd100050000c1f0c031c10100100003000000000c0000d011404cc30000d1f01000c4434fc0304000111003001007000430040000c04000703000004140f043000000004000c1c05030c3400c400011000000c0030000000070400000000000c000c000d0c00010cc300c04403130011c01c30f00c01ccc0113341130f0110c1000c00c0100000003304c0110c30000010400c0000400100104400000f0000000d001c0d3010000d1c4000400d14040cf004300c0304100c1103000000005530000050010000010c0301c1301100000071cc0307003f0c0c010c000400d71d000c150104001c0001700000000000f3000c03d40c0d0030c31c1c0340000100140105003043030003030f01101c00051104300400034110cc70fc400cc0c004004000cd0004005400000c0000c403010f0700000f0cc130000c00333000f0cf040cdc0c003001400c000001000370013d0704001033300004031c0300001400cc4c30010300000f0104000c0c340c3000007f04cdc7000000100030c0000000000fc04400fcc000307001014013170003c104c0001cc307000c040d013c0c010301050c003300000c10000c04c0040041400000000030010d010d03dc3c30c0001d410100040000330001000000000c3d00100103030c00000730000000d1040dc04040f01400014000000f00003d0100103003000100004100010340400300000c0c0f0d00f300cc00000004dc04010700001710010ccc0341cc00331000c00f0c0c0c00dc0154c3300c430400030d33010000000000000000010c03101c0c00003cc00500c003000501300107c0000c003000134000403c04004000c340c003300000000003030001410d000400001c000ccc000d010030000130030031000304001c00000c1000000c3500003c00ccd4030c0500030703000c100c00100031000000301d4700005400000c0003000c3100000c00000030010c010d4003c00003401d40000000000d0404031500100400107101000100d003013dc50d0001c100070007010c0000000c33040c1d000fc03c01100500450100c17007000000000fc30c001000000000030030401cc0c44cc000104440c0001100c00d030010030c0c030c00430c0c00044c0103400c30500c00000000011030040033000c000000cd30000030001c00303c310000fc0000c000c10ccc400d00013000400f00c14000414f000c0075000c00000c0140400000000400c410004300c00307040c03300d03c0000000000000c3010144000c00110001011045040c40014000;
rom_uints[519] = 8192'hc00000103000040004000010000c30410000c00000f00000f00c000433000c035003c004c000c00000000c000000c04c00000dc00c0dd50000000340040003400000300000000000000340c0040010c010000000070004040000000c00010304c0c00c0000000c000c030000430040030000c000d0004004c0040d0044000001110014000004000010000c1000041c030000c00004000c00400000000044100100000000000400c00040c101000000033100000034007c301000003000c00000000000000000ccf000001ccc0c00000000d01c0044440003c0dc0c440000301c004004004000000c00133304f4c34400003010051000000f00000000004000c0c00c045400310400101400340400000c3c10003100400dc000030000000300401c00000000000c010000000000005000f01f00c00000000000ccc0007c03010c0c00100000c0000000300c30000c0030c00400c00141031000dc4000030000000013100000000040500c13d0c0000000000c00000c000c0033000040000c0c00005434300401300000000000300040100000c100001000000000c003000000040c00404c00003004301500000500003d40c0d00010000c400cc1400c0000000703000100c000000c5000000000000070c000c00f0300c000000000c0010001000003000030044007d01040733040000000034c40000c000004100cc0000700040c0000000000c00003000000401000400004f0041c3000c000014cc00301000400c00400000c1000040000001040001c0c100300c004c1030304044000001000000000300c00000010c00f40040000000dc0330c00c40010000c34001d0c000c000007c300703103d70c1004c3033cfc00000004000c10c31000004f000000000040c4001003700004c00040005c30504c0003dcc100400c00000000000000001c1400c0713000c004c0d001000001100040c000cc040c0300c0c00033401030011c00000c000c007000f0004000c00c0300401000c40135003c04cd001c04d000500000c0c000000004c000c10000001000100000c4c300000000c00cc403c04140030c00cdd0d40030003000301c0100001000c0300c044010000400c00100000003000000013000cc0c00000c00c100001404ccc0000cc00001304c1000300c00000001040c01000000c001040004000c0000040c43000000c40300c00000003300c1000414c300000c000104c1c400003c00000c003000c0000000000040041300000000c1110044d00f00000d1000c0cc000110000f0c310403000000c000003031140c0034000000c0000c400c000f4f00000000103000000c1030c0000010f400cf04c00004000003c010000000c01044000000c00010d0f0400001d00040170000300000c0c4000c003000f00000000f0c0053410003000003100;
rom_uints[520] = 8192'h1330c07303c0000004c000000c03c003f1c0000440307030c13fc043010100400ccc337f40101500415114000040c1100c00040d40c030d0330400000040000c0533c301000110100000300cc000c0001140000430f03004000f30c0043d000000c331c04304c050000cc4030100c500c00c0c00dd010cc003c0c143cc0100303103d00410c00035c440000d73001400470000000000c30040300003035f40c0000100100d30d0df040000034010c01c000c03c0003004311040c0014040000070000c3300004430c0f005010140d0c00c000c00401c0f0c0001311c047c40c0c0c004700001d000070100530430cffc1c00000040000001000000000303031303c00c4dd00330d001400c013cc304000530c1cd0503300f0dc000c47034041c0004c00d000100f00041030100030000000107003010c00040300000004034d000c0310540004c000000c0c000740100010000c44dc140300001103003c00c00c000030000304c0fdc5cc704c00440c00100c10c00004570c0003300303000000004070c130400000001000443010fd4c00c04004040f003030003c330000300730f00c00003c03100c00040154000330000000100000030000d0d000031000000c0000c0004001404f3000d4040000c700010000c00c01014434004000440f0d0cc40c0003040011d1333c041003000c00100331130130431400cc15030033f50000c00543c00400300000c00c000c000c0000170c0030c4003c3f070330034110000014fc00310000041003100100000d7500c0040c00000fccc001003c0cd700030101000400004000cc7005011443000d01c0403d00041030333c011c3c051740300f30007c0000041f00c000001410140c030c00c3000f34000c00000c30000300000000000cd0c4313731400041c400003300001c001000041f300001140000013c003014f0000cc037100c0cd0cc0300c04010100c030330100303030040040c00000f1000400043003d073010c003040c3000c07000c3000404cc100c0000003000c100000000000c40000500000c50340400100300000000c4000f7003034000fc00000000000003c40004370000000cc01330000c03cd00c43c100dc014103000000030700303001041000c1000000070c001000c0030033001307c3c33700000000400013c0000c3d0000300344001c73c000c003300c33cd101000001004030004000300000c000cc04000cc073003c400010100000003403003c0000043300013c01003cc300000cc01000c014003010000c4004030c400000ff03d0007c35d01400d000c0044300c3003010300000000403100c00034104400000d30c0c0c43143003050cc040100000000010001c010000000301c3dc0100010cc030003c103cc0000000000c04c035c4000c31000000000c0000d4010c04;
rom_uints[521] = 8192'h4cc001010d00333010000101000c00000c000001101c00c030300000014010400000010300000010104001c4d030004373000d0000000000400030010010000000c003300040003010043040c0040100340000400700000047c0f0c001f30100100000000001f00c00ccf001000010c000030f00d300305300000cc014cd0003df0cd000007000114000004100004000431000000007110001000000cf014c0101040331c70000030000000101400400f00c40c000074cc04c400c3f000000040040000100030000f000010300c000d0400c10003010030c00c0c00005c44010c1f000c0c7401000c1c0004cc170c001407031100010000300300000303001400000000044500007000051d304030100c0301400300c770333d0c30c0d04cf01430000004300100d0310c00c5c430000033cc000d001000000c00c33500000d0440c3300433d3007044005000040c40000f403d100c00fc0400cc100c7c01000c3013f4c0133c0030c000000fc4dc0c00c3d000340c100013131d0cc0041c47103c5400001000004000001cc10300d00330f10001003000c03c504300410017d3c3d413cc0c04010300403000100c04c30100400344c000c01c01040010300d00000040033300007d0c0c000000c0003000003700104c0c001d1400300d0303000413330001010c043c414cc0075c0001410003110003501010010004cc000d00000c04c30c0001130540003000004371000300130d0004400003c01000d0041100030750f500340000c03c0c01054001000f0000033c01c11f00007100f3000f3c040c04300000030004001c44f4030044030c0c000040017000c0c401dc1c00031c004c0cc0003500330c0300330000003c0f14000c300c4005300cc30100003c3000433300010730303c0f04c00c10c5c0440f0010c10003f0000f0030100f300c051010f10030c0f003c0141013d4c0010311000070100030000c30110000005140010000040c00000003c0c03f040003d1130130c01f00030110c700000400303100033300000c000c0303101c0030100000041400001031000030030c07110004750004c10040305c01000c00dd00074004c400040000400100000c13430030d033ff0000000c0304c3000310303004003000003000c300f004304c0100303c0410013004000100007c041f010d00004104000010703cc000000000340003001700100070cd4d000d0010341400033000410510030c1000c004f00cf0001004030c000c033400000d000cc30511c000000010453031003c00000c0100034030403004300300300340004c033f003070003000c4331000000030043033004d01001300c30c001c1013005c004c03000000000030c10c0f0c0300000100000000014300007030c003000030c7040300003330341d4c330c003300005000;
rom_uints[522] = 8192'hcd000000010d1000504000004004001c3c00000c1000d0000c000030300400000c0c3cf00f130040004c000c40ccc000cc3400000c000c030c001000000000007030c03c000000111c000c0030c000c0000400000044c010c0340304c0000cc100d000000cc00c1c0000300000040001001010d404f00c040030c03047c0000c704c400010c000700040000434000004007000000040100c31cc0000043000000001040010100310000000c000000c0000cf040000041000c0000000d0003f0003000000300000040c4f0003d0043040300c0c04100033100cdc040004110000003030000000040c0000007501c01000c5000014000000000030000cc00000000401100c0004d000c004000410040c040440000330100004f0340004400473003c00c000cc0c00040c440c0000c0430d00000c00000003003c0c10031300c0000c300040040cc0000000001000c0401c4050300404300100ccf40404d00c0000003dd4400c3003030c0c4050000040040040001c300000050cc00000000cd100144400f30c0004400c041c00000c70741000000000000000fc004c100041dc0000d03c00001c004000000304c10c040cc0000011000400001004034000041047001000000010000c000000000000000c041040000fc3000c0000000004403403c000cc1000cc003400400100040034004001c403004010c0000c0400c0030f340140303004010000104043c000c4000430d00010cf50c00c00103c7f030004000010100c330d00c00030c0047000000071c1300c030000440000300d0700c03000310000f00000c0c400000c003d00c010c0030000504000000d3c00000c0000c0cc100000ccf0c000403000003000000410000c0000c0400c440000f4300030c074040c0c00400030f70011d11040cc400c00cc33001d70000004003c4fc000cccc00540000c01000031c0300000c3c4f0040c0404000040c00c300001c003c1c00454000000010c04000000c0300d000300c000044000d301004004000303c00003c0030c0000000cc100400400c50000000d000400c0010300400033000000cc030114000c0001000044300304403340c00310000000c400004010404c00c0034004c00000000003000c0000010c00044c07010030c000000000c0004f4000f3000000c440000000004c000003000003000300c0100c000073000000030100030000c0c00000c01043010043300000001000000700ccc44cd003f01c4001040001c300c000c101000303134c0c04000003400300c31000010f30030000c0c000000003c0040c00004c000300000f00030003400000c0000040c001c00c010000400f30003c0cc003444c000100000c0000400000000c330c045070004000000340c1c001000ff040000000074cc0c000000cc000c4cc00cd104000000003c;
rom_uints[523] = 8192'h3000000003000000000000f0300000000000003101004c000044440000003300000040d040c00030100c1000000000c000143004d000004d3000000030000400000043011000003304000fc10000304000040001c04700000d04000400c004d000314413000000000c000000703000000000000000c400c004d3000011300000003c0c00003d0c0004040000140010040100c00000c0100000000000043000170351000001000c000000000cd000c00310000000000000000000c0cc00000000000007000c000404100000140000404c0c0000304000c40040c010010300000000d0003000430300c44c000d000c410034cc41003000000134000000013000c00040070000300000000004000040003c10000c1030070300cc000000000c400000c0cc0000010440030040040000000000c0000c00013c0003003400300401c000100c030004c0000000007c0043ff0010000000000c04003001133c00000c000c13001001030004004003d4000030400014100004000c7333c03c104040000000000400c0030000050004000000030c0000340100040400c00c000014c00000307c0000001000400000c00c001310000140c400d00400440004000000001d30d0000300031100c0401400003c00c0c0740c0100040130001430100030044030c000104c000c0000000140000000303011400004001304000c0c040c00003340140000000000000010f03c0c000000000000000010000c004400c10000c4033000dc1c0000f3000000000c003000304000003000001c00c000000c0c050000100cc03c0c00000c300003000010010000003c030000001000cc0000d0fc4011005d0000304000000f0000c4000000c101400000c03c000003000030004000070000000400001300000c003c004c31f10000303030010c0010000430100400004040c01000001c0000c000001cc0000000c0000010100d40000d044c300037c0010003300300000310d00010000000000000000030103000c01100c00c3000000c4300f0005cc004000003300000000000000000000400000040000000441000000000000000300c100004004000c00000313000000340000c00004c000c0000004000000001004040403100300010000300d001d401300000400000300003c4304c00c0300001003000000c00013c1400000043004000000000100000000001000000007f0c0f00040300000030000c00000000000000c1c00c000000000003000100540300000c00000000030000003c0c034000003c0c0030010004100300000c10143030000050000000000070004400f04f0037000300100000000000410100005400c0cc001004000000010c000000040c00330000040034100001000040010c00000400000400007c0034ff0000050300000000000c0c00004000103000;
rom_uints[524] = 8192'h40c4030000440000040010000100cf030c0300cc00d130034001030003c331cc00c40300033cc0004011000003010000040403001000004c000040000400c3107cc703004000004c0000040c00000d030100010c4c070000c000074004011001300100500c0034010000c1000340004c00c0074005000000114343c0001300034004c01041040003400000c10000051101030000003300c10f3000400fc501433c07c00400034d00004100103c00071103004d00000040c300101100404300000c1c1001c3000040004101000100c3000030f0014c0f400000034003c401c00300000000c1c40000000300ff000d000300303301c00000000300000c40014000000143c0007c00c14c7000004403011fc7c43035c00004405401000000f31300c00000004300110d00c000c0d0000c0100010c030f00030074040104410c0340430000100d4033014000000305000000c503c0014cc0d340c000cc00400000c40100400413c30307c400ff11c7c00cc300000000c0330040334030c730c0030040010000414f03400f0000000000c50000000c0300000c034f300040000c00c0c00cc00041040103000030711000c000044001cc404001c140c007000f0300400d004040040301030100000003003c0000004003010003c3000040004000dfd01304c000000c4313c304010313c00300c000000100c001030c000000d3ccc3c30000000700c00351704170400150c34100010001c000000c00f00d00c100001c040c0c4034000040000043401c000010004500000140c3c1401d4303d04000c00300010003030000030000000703c040004d0000f0c0000043c1030300003343010300c0030000000040004f0300010073004000000000000000c005000000c000010000c300c04100f743001d0103030004c3000c03c0d000f30040100304400000330000c00100c000c000000000c3cfc101cc00c000000003c3000000000c00c0000040000000304300010000034c4001c00004010044000007000000100300001000070001000031405001d100c000c1dc4c00014c00400041c010004d000000030101c707c0000041004304430001010010c00c00000041010000f340c31c0c0000c3411103000740100000030101011c31f1c00001c30001f000004f030c00031000c430c000401340340017000033030000400045c043000041c0033101000404c3cf1c00c04003c0040004010044011043004005704d000c04dc1300400c0c0734010003014340014033000d1c000fc03000100100435000130700000f0000004dc105700001057c00004000004140034300000000300000000430001041500700c1cf000040cd40003000000000c40043044040000100000030101040400000040530070705510010103c0074000000000c50c4c000001c00000700;
rom_uints[525] = 8192'hc10c3300c1c007d0cdc4c000f37031dd010c00004040400000011c400000035000f0d0430030004c03510040cc400d43c010c30000c0c0430000c0430101c4c000000d304000c3c00000c3f04c000c10c000431140c0000010c0400040400000003070031000000033d04030d0010340cc00c03f00c0d00000300040000510c030103000300010c0000000000100440000000000001000c01000c000cd1171010000010000cc7131c00c41d0000310300043400300004143000031030cc30000104504000c00300300f40104004050004dc000010000c000010070c001010030030030033cc10100c04004400040c1f010335003d0c4030001cc40c30100010cc0c00013300c0c04c04400310000c1000340c5301043f3003303c0331c4303000000c00010d0cc03005000f04cd3c0f0003700c00000030000070301c111704c40c0404c1001cc0001410cc03400d00341c7ccc000001000d0700003c0c030300001330103103101cc1301033f000003c1000000fcc04700c370340c30c0c7000001400d10f0c340c50300030000000d0300c1f0410cc50000f000d0300040304041003300c40101000ccc30004043c00007c041f00341c0c0003f0140c01d35c3c0d001007c40d0000030010000c001403300c0c100f00c00f01000005d7cc000c0c3f0030003100c0000d300ddc03000034ff0c0cf40c0700103c01c01700c44004000c0c00000400df00301331c01c1100000c3003413c333000134030d500d43404d0dc010300040c4d4c100c0d00033c3100040c00100004d10400000cc130040c03cd00d0041cfc13300100101c0014000401000cc0000c0400111300410100000c10000dd4300c3c30f003c401041000c01c0003730c140001f3300c1f030f00d11401033f0000100034110000c10d011000f07000050d011f0004130c1c0010c7103435104000140310050004c00c04f3003c31130c0ccc0c01101000c00030100000000cc4740000000001040400000c330010c70d0c0011041d0104d0000030c330300000c00f4003400003007007303000c000034413001c000c410301000340040000001d0030310c0c75d0110000000d000400dc0007740301051001040c17110304100400040034000000000711300031100400034003000f330f0f0c0c0704000014001000d50c040c013000050040300307c00000131c3010040f1f05070004d010000031c01c000400300433300505144c300000001cc4001d04503c00030f3110001405100304001c4c1100c004140f0000100400f00c1f070f003001c01100130400440c300c000400000c500000000000d004c41c3d0cc05c000310cf40040304500004001c001ccc04001d041cd0c000f350003001001100c000101003c00c3000300000001454130c000004c0100c310301d000003;
rom_uints[526] = 8192'h401000110d0310074dc0005010000130014050330000040001000333c000c0000104c3cc503000cc31030310300304300430140c40101c000c300cf4dccf0000000000300000400000343010010c0c0c000030c017400140d1f70341c714000000300c04000000001430d00333c4cc0040001440171730000d4073103100013014cc0c00044000004040d003000c000d014014003430c13430010030f0f000c0d0004c00000c4000c001001c01000300d3d00000f44003c410003030500000041c0040003000c34000004004030ccc0500050303d03070330013c0003001100001033014004000000300ff0c00003d300030d340cc005c3001001000010001c0c000400000c33c10037c30000300c01000300330d303005d100034c4310030c10040003040000c00100000004cc10f4003000003000000030c00300330c00030d000301000310003c030400300033400c00417103400037d01c3c7000c10413030003d4050f3003c1f110040000000000130011d33400730000000c00d00405f0744007cdf000001c30400cf00dc3c0c003400c000d4004c1114131cc000400c7cf4000c3c411100f111df044fcc0075c110c110400430c000dc0001c010c0000c0c035443031c00cd0000f000c3003300000041004fc10043330010f00040000c7c01c0050c3310003c10300000311c0cc0c0303c45013300003000c00f35001fd00500000310cc004cc00c0004040c0001003411000c00004100030003003d4cc07c40003410007043000cc0c1004d40004310000050c000740d3c00c11c3331000000100000000111013031013403c03174c000700003cc00004c0011c00cf0000033f000f053d030107c0000030440d0c0000074000340d440c400c01440cc04003000c033003440000f0111f41f40f10010c44cd00034c10c0c10000034f0405040000070030000003073307014d31000300fc00004000d3104340000d310700000000c003000c003100cc44000034010040c304ccd4000c030504c10300050000000100000044304400c30000f1000c310300c103300100001400000410001c0054100cc0cc0040000c50010c10cd00f010530cc000040c0000040f0cc0040c03100740c103d0000c00441410004c0d0004101000041100000c0501c403ccc00c010501030334000050010000300003c3140000000040000335131004050303c00100040cc7c03d00404704700000040003003301113000300c0000034f03c0473000c4c010003403f0470313000000730000c4013c000003c00000dc053c000000000f70040005cc4003030003c430c0000500010341000413cc43000030c47111034030013400004000000c00010100347000c10030c0034c0104101340c0140000700044c0300cc00013001000c10c030c01d040cc0403500300c;
rom_uints[527] = 8192'hf004000c1c0c04c0000c0004100c00f0cc00c00004c00000000c004030f0100000100014c40000d0170030030404341c0000c00133001c0000d0040000301c530c7004000310010c0000000100071400c400111070c000000000c000000004c0f0f000cd0030050c0000c00005103000003cc41014050c004100044c10040040003c00c001403000401403040000044500000000010100500004400003303430000004c000007030040c0c10701000400c0c000000444c0000000001000c00000010100c000000303f00c000c0041000fc0113010c00f0000cc4c0100000000000000130710000000c301040130d0434000c0004c4000040c05c4000040400c00000000400000000330c301004043c000c000400000c0004003c7d50400000000000000001404040010c0030003c040000fccf3004d0c034000000c0c704041500d03004000404f0000c0cc040100c0c0c4010c40f040c500330f0c0000c005044000340c0c03040143c3c3004000000403040004d10003030c013004c0cc0c004144014333c3d041400003c0030033c000c100100343dfc0c0300040000c0411001000010173c0000000404cc0c3013000040070414404c300050003004c0101d00c33c05001430110000d000c4401d000c0d000330c000c4c00014f000c0030314000000c0000000003d44300c0c34000c0030005000c0d031041400001c0400000f0430c0c00001000cd00000100c400c004005030000300030f01c040050d01c40007c0040001fc11c3c0044c000000000000c00c3040000430400541cc00c3040100c0c010033030c030000100014010000cccf30000d4c4000010c0104040000c310004100d0cc0c0dff1400400000001007040cf010c00010030004301c0003000400c4003034300c00cc4000010c400001400000030105100004405c540005c004400004c44000040c003400000100000c00770c4404001c0cc000000101100000000001100000003f00000004dc30c00000400c040014f3140413010030000003004400c0001c10040000c00000010c00000cc00001000000d0004014400d000c0001000010f340700000d4004004000000004c000010000000100c000000430700c0c00c04c0100030000430c4030014040c551000003c0cc4f0403000400300000000010304dc303001c13f00031034007413100100140004cc041300030003004c33040c3c0c0004340010301c0440c4500f00000000100d010f10c570001004001000000f5000040000100400d33040003030100040000c000cc4500cc300100030000000c73000c000c400000000001000001c0040000cc000733cc4071ccd0700c0000000410010001000700c1c0005030010cc14100040401014110c0cc003007100c4001c0014300000040c00005c00411000400c3004;
rom_uints[528] = 8192'h100000014c0001000000000f04f10c04c000040304000000004c0000005000000c000001040000000c000000040f0340110c00010005c4c000000017c000400100010c040000400000000400c0005ccc0000c01f3003000000c1cf0000410c0003c0fc4000104c005cc000404100300000000c0000004001033000440000000035fd000007010c000c000c0004c4c3003100000014030010101300400c0c10c0c3000000300404000004000000000003000001003400c5c0000010431f00004000000c0000500300c000001c0000c0040c40000000004000000740000d0cc0000c0c0030700000000000140d400000000045000000000004100301040000010000003dc40000d1f00300410000000000c00014000004000c0400cf0c00010000000c004141000440c0040400040000500000000f14c00004004400334c04404400000c0400100043c03c04c00000000004000c00000c0c0cc1c4c30071c00003000000404030144cc3000000314c303000410cc40301040007c700c3004000040c5f5040003001000043003c4005c00000400f000043400cc40c330005004c314f0cc000000000000c30c040c0010000040cc4cc100040000000c001d00407010340f5000f00000c300400d0c0030404c00c0030043311000c0040c30d00000c00cc000035c00501cc004cc00100000000130043000400c30c30000000000404000c0c0100150400040030040f00c40404c14411c00000000000f0330000000000043043300c00000041040c0005000000010000140403c000400c04000001030c0c4000030f00040c00000c000c04440c0c00010004000005403000100c0400114000400c000c000c000100140000100c003140040000000f00c00c0c0f000cc70000040000c30f00030000040000c3010c01001c0000000c100530040c0010000c400cc00c01000000303400000c00c4000000004005c1000c0c10000000430003004000000040000003000cc00c001000004c070000c400110c0c050000400000400100c404000c00000304001000000000005c00000c0000004000000000000000cc4c0004d000000000110003000400430c0104040001000404000c00030000043100400c5f00000c100000003cf00400404003010001c00c050003c004000c0000c400000c334334c40400000c0000000340400010cd010040c01400000001000c30000c000004001000044c30000c4000c4c0040553000400005000c0000f10700c0343040c000300004000c00cc0010000c40040000300040000040430c14043001113000034000400040f0000000d40000101c140000031c0001003300c1c0c4040f00cc300004431040000c00400004000000040000411c0000cc00400000300030c04c000004c040130100000000c0c0c000c14040000000000;
rom_uints[529] = 8192'h300f0000000d04040c010c03c00500030d00000d040c00010d0403000f0c0c0300000d0500170000040c00040000050100000c0000030004000101010d000c0000031f0f00010431010003000100050304100004300000011100000004010037000d04000c000c03000c0c300c03000000000c040300001d043100000000010001000f00010d000300000000040003011100000000000c00150000010d000c1f03100f30000c05000f000014340101370000000000000103000304001d010c0304040304300d010c040100340004030f0104040c010d3400040407100030030300050300050f0700003400040300030100330003000000000c0c0f071000000c350c3033003000041303040f0cc400000f030f340c0403000300000d01000c0f03000d00300104040000100330030d400004000c0001010100000f010400011c00010d0001010d00003c070c0403000003010107030f04000f010311040c00000130043d1d07030c030400010003000f0c000004000c000101300003010000010401c00000000c050d1500004303030d0c00000d00000300000c300001040101070003000400100d000c3501040500000301073004040c00000003000c00001007033c0f040404d0010103010f000005000c01000501c10300031000050004cd000007c300300c030405040040000000130304100f00000c0001000c040000030501400d000003070431030c07410001000c0300300000003700010107330404000003000f330f010000000003030100030c030305010c0300000c00100c3d0f0000000000030c0001330d0c0c0c03050d3015000100030c00000300000015050003010f003f000305000c0c3d001031000501100c1d00000f0c0f040331010c010003300d340040000c040003050c0c0d4d00300014070000070c01000f0d030c03031307000c0007030cc4000003030000000300070c00000100000f000004330701c30c0000000c0300000c1000050007000c0000030c33000c0c10070d00000000043d000403030000000cc500050400004d003101073300040000000300000c00300000030311001001003c00004300000c0f000d03000f0c050d00000f0001000004010004070305000010000104000135000000000c04030d01000500c110010004000503033500010d000c000300033c00000c0101c10000050301010004000f0003000400010133000000040700010404010003000100000000000000030f000000030000030030050c0c0300000c00340c00000c000304033c00003c0504030030001005040501030003100000040f01010003330d0000040100000c00340700030c4300010000000c000301000c00030f04040505310c03000001050d00050000000d0001011c010c0d010100040c0f00000701410c00040f0c0c;
rom_uints[530] = 8192'hc03c00033310101010001cc0000303414030010f041cc00000c30004353000c3333410100c00000310f0001000c500433000000474030000001030004000000000f10000f0c370c000334030000031110550111070c031011001011003000030c013554300001c04f0c000dcc1c15030333010c33434f0000c4001f050000400401000033c000001401370000110c1104000c0000000c00043000030003c10000c101003413443c0331301004130303000071000f3004400d100344100000000001010c3001341435331040301000130c1c003000c007031c040040f51400000c00010100013000050103051c00000300cfdd031d400104000103d40000040c01003c0f0c140c01003070001404000000f0134304303101134000340133000f0043f00307173400000040030010d34404300034040c03030d01104034103330310300030f000034400000003410000300170170c0405540033c0c41c030000c0700333400c11410101f3340000100030000000cc30c3c3c0c5c1c7c50004001010534031000400007044034000431100c0011000004000031d4031403033101350d1c0030001c000007340c0700004c0d340400000303040053033000000104011110033510001003c00730000000043105000000000cc0101104005300c3c0030410130d01000c4000304030500000001701000c00000103c00c04d00033f004030c10030004500d0330000404c03c300104c01005000303003c354000010c1001000f330c33f0030051113c1c100d00751300010c1c04401034001104c300410034f7000c30010443030334000000410df0100303c00043000400000400c1cdf700dd00100d030d34043000304414000703330051010c10340000440003cf300044000040305c0c0f0001040103135043f3100f0441100341540031c713000c14000033000311100404053c05003f000f001033cf00403f033d0040300f0000010c00300000c3003030000d0034c001033c404100010c0447000c30031c0c0001013003c01001003101003dd000000fd507c00033004001000d0d000f0c01cc000000cf3001400000400403004104cc0001030c007c00050003300000fc13000003000004014100001300030001333041133001f0100000000133003001030c0430330000000003cf3001300341070300313c0100dc03044f000000cf14010c0400400300000131103000133f0304030000040c0403430300301004c030010005d30f000c0031c00300000700c010504f0c03000130034000330030030c0030715005000401040040001f30000c4001c04d0000030c004340000400fc04000c0373c003003114c0411c0001034007005d010000010f00434c000c130c1d000000000433004cc0010d010101c01300040030011000000110040400103c310;
rom_uints[531] = 8192'h3070000010c10010140cc004000400d73400343100000040004c000f300f4004540003541150040400000040317c4c40d4400130343040f31000100cc014000c000c100000000030d0010ccc300300034004001001040000304043c015c700000cc3410c30000cc000000c000c0003c00000300400404000c031c070000000c3c543c050ccc0000000000100f000d07004000400004c003c0c0104004010d1100c50400c314f3500c100003001c0000400d10000000050c0fc30c0010003400c134400100000000130000030400070c03c11040000030401471001c0400001d0050c00c0400000c00cf00d30c30044cc30010cf300000331700c41c0000000c00000040d73311c005c00004010000000500001000c003541d070c01c001030400030000011c14030101003050003003000d03fd0c03c0030340400c4c411043000c000507001000f30401c00d000401003c500c04074030f0541400000c304504001c005034c4000c0000030300301303c10c0500000107300c040000000c10100004004000300cc00c0c0cf0c07540030c000001400c13017303cc40050000010331c030f00000000400c00557000c050031030c4c43004d000c0000000400cc003073000c400040414300040033001000c10440cc404000f3cc0040403017003001c0000c0c730fc1030c003700300000003000000010fd170010130d34400403040c014000cc01f0c40c00070c0403000d0400010003003000003130cc0000c414010700140300004c007510103000004000c01f140350c0030400004c000300440000003cc00c0c3010004c0c00c0310114010f57070040300030000000c0400044000070f5c00c40000c400000c000113c1003000000140cccc0540073000d00030040c300f01003f0f1007017cc4c450f30ccc03000030000440c47500031cc14013f00000413c0dc14040c4000000c000c0c0c0441000041c0050004040030c000000000100004040070000d0000400100c0304001d30cc700140300000030001f400000c001300343c400000000c30030c0000030f0403400500000030401c341000100011044c0000000013c3004370c003000000304403c005dc50103050400004cc0c000004140d100040010c4171340f0001d513001410c007c030d7c41000c043100030c005c00431000000040f430000100cf330000430001c4c40c30440c0040440000000000130711000400100007053cd0000300300300333c040000000530150033000c000703140c00310044c300130010000c00003000070d00000000d500cf0400413000c00033047d3000400300040000044c000c03000000000430103000000c035104000003000000f3c10c0005f300f0007c0103000c00010d044f403c0f0c4000370000000cd03d003c30c04004134000c300;
rom_uints[532] = 8192'hc01c0001000000001cc0010d03431c1f0000c0000340113001000000f4000cc4000407404c1c30004c0c040004c0307031c0003d00c00d0001003000000040c040001400100000c0300c4c4450010c130c5000dc34000004c0035030010000f050f433004001c030cc0300000c30001003143000004440000c371c40010300043fd3033300301f00303140300004c037005033000c147d00104443c003c0c0130000c3300440fcc033040017400005700400000000c0700014400c470030c1434c0c0101000100001c0000000c5f030c07c040000101304300300c0004f0000c703130ccf4dc0000000001f0c0f00cf0c3070f31000000033400000c000001c10f01c000013cd0c00c05000311c0000000404010c4300000c340133000c4c0dc43010007030001c001c00c07031c303704000c000c300d00030301cc30005350d4000dc01433000000001030400003044c50c1000151c03c1003c1003c0c0000d140440330740303c000340100f3001f034c000034400100000d510003f30130344c30005000000c00400100f100031cf000000d00000001400c07370c50343cc4374030cfc3c700030104f0000f04007340310c004050304003300d3000003c530131c70c3004410f100014104cc3005040040cfc05ff033c00d4031070c000000010d01001110c4c01c57f0001010f500103403040c044011c000cf100d500000c00043c400054cd4134ccd0fc00501530000cc300d10000013f310d01c00c1110d0004340103100d300174303000c3043001040fc500c04c4c0c11003cd00400d0514000340035c3c304000f0cf1c04001030000cc0030000c40cd340740c1f143030f01c071133400000f000100110f40330c00004030c01c000034030000403000000010c030000c04000045013404400014000ff0000c01001dc000300030100013c1301040000030450000041400150c00031000000310405130d000fc00d3000300300c00000c4300c3004f1000433300c341004301300c03c10cc0c00003c540f00000014300c003cc00f0000113440300000114303cc40f000000fd100f34301340f03400300c0040000000c14000fc403033c00c1cd10710003df0cf00c0000c0c74400300d43000000000c4333030c0c000c400043c404043000344550300034310000c3c104c00f1c040444c330c1cf0030c0070000000000004000c11001c00104000010040100c0c3000000cc0c10501c10000004c304034010100c04f00c00004c313100530c1f0003c3001d30015004004c00000000000f100305c0c0350300cc000453700130c00cf10540000030100000c0000430101c003000c400f030df001cc1f101130c000cc0404000503f000040000c110001033c00004044300d300730304005c0c00344000704f700f10c30301c0cc0c1000;
rom_uints[533] = 8192'h37c3c300000003cc000104344000c10000000f0110d07000073c00001100c0c70c0107f0f4001c030c00c00040400011000100017000010c01400004100300001c01d1040c0030011004f0003000410c04001011540000cc0400040001000c00c00040000000110000f0050030401d000d000f00300004d00300d0d00010000ccd33cc401000000001100301000300010000000000010c003001000000030100f1030c0d04c000000d3000400c40301000c70c0000cc4d0c00000101000c40000cf04c04cc0c400100000c000c0044000c000c3004004001700005000c10030001400000000040000d0004001c4100003c00040cd0000000000c00300000040000001c0407110c444c0000c133000401400000010d01000d3000c1100c00303301303000c1c01041101000000000400000000045001000c004c100400004c01d440c0c0c000000010100010131101000c1431000311c4c0c0c00f00101000400400150c0000004010044000c403c04f031410037010c004dc500cc4c000d0400110c00300001040430f00040000f000000014c0000403000000c00031c000c00010dc1100c000000000d00037c000103341c0000d0000000011300000010000c3140004c01010000100000033000cc0100c005f4000404fc0040c400000f013fc1cc7010fc1004303000404f1cc0040130000c03c000050130f0100d7030370c10000030000300041310ccc01c1000040c1c400cc000c0043000040c0001c0000c04013430130010030304040100d00545500004400000000000003000000c010c4c1000d30000000044040000010c00000c3c00c1405000000000d0100c4000c00100f11c130c100000054154003000130004440400000700040c0d400004000000430000000014c000ffc05f40730000000c00003000000f710400407001000d01c1040003dc00300d043c000004c0c0100030c000004004043030000400f400004000000710050030303000c000300701001004000c433501314043000400c0000c00410044c000000000030000c0c0cd05d00040303400c0c30040040400000300d004f00c00000f00000000000cd0000000000000700040500cc110c0000c0c000000040000c4000000000d101000013000c034fc1130100c00001403c00000c000000f0c000010004c0007cf04300003df33000010c000c00c00000c0300300030000000000000010000004000710c014000000000014000300004003430d50003000301000000001113c0d4c000340f0100d000014100000000100440c003001104000ccfc0000400300003500c443704400c3430041dc000000cf00143c013c001c5f000000c0440041007000c440150110c040000001c403000307c0013140430c0c300c3347130004cc000000000000001000c100c00000013000;
rom_uints[534] = 8192'hd000504000000000100c00100c0c00700000c000c01c000003047000000c30c401000403030043c0000000400f3c0c00000000c00305c3000000100504cc003010c0c044000f000c03040d70040c000105101000000000000c03c0000c70c0010000040000ccc001c10004040c544c000c010700001f0cc00000300d0003c0d0000004000100000070040c000400010000c0003cc03030000c00f0010d00300f004cc400000000c003000100100c3000000400c3003003010cc00100000001000000100010000003030c3500000000300c00400100cc00000050001c0f10003305404000000040c000000c00000c1000700000c500cc00400300000000c0004c010c0c01300000ccc40740004401400f00000000f00004340c30004c0c00000c0c00100c051000c00000014010000401c00000000104100000000000c53000103c004004000c03f01040c000000004c0cc030f1c003cccc000003c01100d50000c00050c0c00140100c300000d0043034140040300030001000010010044cf10c00104041000000d400c1c1000000000000400030000000000d0000001400c030400000001000000000cc00c000cc003300c0040150145040005d4030000400101000000001c00040001c0054c0100400c0010100030400000100c000303040400c04000010c700043340000000c0c000000000c000c010f0c0c10c0000f003c4000c00f050400400c5c000c000c0c0f010c000440300400300c00c010050c0540c00c0000000004f00001040c04c000010000040000000000030cf10040003000040c0303000000c50c0005000000010c00000100000040c00304030c40404f004f00000000004003cc30000c01c00303f00040000130003c13400c0030040000c031000000044004c00f340000400010000c000c03000c100305400c0000cc000c0040003d000000c0001c0cc40c000400033000004011c000300000000401c000000000c0004c0c00001000400000c0000000000c0c30300c40ccc00314c03c000050c000010000010010cf0c0f500c000004c0040003310010000000040400000104000004000000c0140cc0000c300000300070000001703000000000104c0040c1000f0c1003054c40000000400c0003000c030403000c400000f0000000000cc04f400c04000fc1c00001c04000100c1f1000000000000400004040000c000c101010050440000001100c000000000f040c3000001011000030004040300c0000004005000c0c00003300000000404001000000014c0c0c0000000004000c000000000103000c000000100004000300004303000c4503000004000f0c0000000c00c40000004000010000000000003f0c0dd004003c000400100c0001430000100c400030140f000000300c01000c0300304400c00c40000;
rom_uints[535] = 8192'hc400000000000013c00140003000001010000040c000c01000104040c003000000404010304000c000000040700000101003014310300303000000000000c0003000030000c001c0400c00103000f00000010000030004c3f0000c033100000003c1000041c0001003100000000140d0c0c001400c40004000f1005441c050003f01730040000c000000000300001c4000000010030000400100000c10c400400c00000040c30300304000004040f000c40000c00010004010000000f000000000000000400000050000010c0000c030004040000040000000404050c0c000314d4000400000000000d0030001d3000003f0c00000000000c0c0c000000004110001005c00400003000070030dd0000000c000003c004000000000c000f00444400000000011013001074001400000c3c0010000000440c000c0c001c0c00000000003001000c000500003c140c040c31051c044300010000000000010c00030300140cc300030c3000000000070c0104074530000c000030100000030000000015000dc30004000404010000000c0c00000000300004040000040c000000000000400005000c000c010400030307000c34100c000c000c30040c040000c700010f00300000040d071400304f000100c000310c00144000000001000300000f04000000030400000c0c0c04000100143c000c01000c0c30010000030000000000000430cc00030001000f1c3fc0000c000c000c00000100001d07000010100c0000040c0010000d000000000404040007c0000c00040c0c3f3c00003000004000c00c0c1d3004000c00000004003c000000100c10000c0c000c00000c00001d0003000c01000c000014000330000d073c000c001d0c0000030d0c0031000400000f041000000304000003c0050c0400040c0000003100040c01000d000000003d10000c0c010c04c0c3007c00c0000c07040000010c00000400000c040c00001000330c00001c0000000000040d000000003440050303030c000d00301f00000000000000000f0c00000000000004000c0000040000000000003300c40c000030003c0c0c00000404000004000c0000c00c00000c000100000000040700070c3001000004300c00010703000300000000043710001f03010114000c414015000c000c000c0c0000001000000000010004000000003c0c03fc3c000010000c0c001005430001043c00000007000000014000300f03000403300000013c0000004004000c000000003c00043307000000000cc30c0030030030000000000c040c00310c10000003c10000040004000c0d00003013f1003c3000010c001c000d000010c4040c3001000c00040c0c0c00000000000c00000000c5010c400000000c00010000114c00c4070310003c000d000000000000000400010300003c010c10;
rom_uints[536] = 8192'h100c040003433000c1030000c330303f000310c13c300c0d00cc7003143014000300013100000000001f30311c3000c01301000101144314000000400000000004c00171000001103000003300001001010400c1c043000000000134c00004030000000330400d0040004100010f000000cf10400003c0030450031c00cc00000003500000000040007300003100c0100400003c000d0000010000003010040140c01004030f11430300f0040301c00110000410000313013030000130050400001c00030300010030400040c0f0400073014d40474330000100001010101010003000010c00031000300000045f000c0143003300110000000000010010000000003003501143d0000045000030000000330015003400cf0000100f000330c00010030003034340000000004000043001307000001000000000010100003300c003001000f33c034030300000cc000303c1030010031334d00001c3000010000037003c403cf00011000c703400c10f00000003000c070005430f0704000c030c30040c41000001c100003033010403110000c0050004000011007003000000304301040104c3000043103500000103040000c00010004303c03010c0030c133c51000014003c130c000003c5f030c0001100001000000001c5004013f0300d0000000c0011c00300000000430000140004000003c0030003c00000000d000340300c4c0f5000c430000003c04343330c03100c01103340010000300c44304000100001c04400030000030034000000135010004435c100045000011000030700c000000000c000d00f3140c000400300d40f4cc00000000000000300d005f0c00c000c4d00000373c00c734011040cf0c0c04f431000000353050007000f0030c010c0000000030001030000000c0003140000304300140000010413003000001034100300003c0100003301003100030100000130300000000000043000034c00f000500003103c04f0cc0000030003003001040000000c000f00330000000000c3000030014301f000304010c0c00c0c40313d4000000300400011030400c3100003030000101100c000000c030000041f007000001031443014103000c11011100403030100010000030c000100000c01700103d1003003c0035004010401014303010430000c704300404010100000500c01010dc001c43c000ccc1003000304c00000010cd110f0310000000043030040100130030000000100000000000033003004000010000013010c43100313d0c00003f0704030d00030000010f0330040100000c304143310c100103000040033c7000c00f437000003c0d000000303730c4073010000c373403c0c1000c1c3040010000000c0040110c01003d0031003000c03310311015c00c0c00003000000000301033400030353000301;
rom_uints[537] = 8192'h100030030000000001100000300d0cc0cc4c004000c043c000030000013401c140000001c0c00000031400ccc10c44333043000001400c43c030004004074000c400c000f300131c000010c145001000530331d0040440030400c0f403f013c030404c5ccc00c1400000334140c0070004030440044303354005030d7400010c05c701c050400005043000071c000034004040330000000001054f04c433fc4f0c00000cc107400c40000c000dcc00c0c001000d00ccd3fd000000c5003400c10c04000c00000dc01000000c40c0300400470f00005001400447000c010c00040003000100010001013c0015c140404404000000c04300c003d010c14000000140010cc10014c0010d0c4043c00c0000c0c101410f4c4c00c007003c14fd0104f004030000430000c100000070c0001400003d01540030000c00cdcc13d014041000c1030003c100440c0c0c031000030000c14443c0d00f0c01d4004f0040f303c10000f00041000140c30c0001fc3000003c3303c00c14fc0100d04004300c47c3030010c74000110c00cc30003cc40300401310001400037005074010300cfc31f100c040000400000c40000c004c030147000c00c000cdc0070003d04400dc0d10000003c3000103000001000001cc04c003c40070400401ccc150c0c1410040011c40c0c43040035000ccc000143003000cf000c30d00403403100c000c100017c43c07c00c00c10c33430730c0430fcd00f0c00c011000c0dc0c1000000530300f0340c143000043144000c00004030400414d0400dccd0c00400044c100000c0040030000ccc1040041300010000c3d00f100c4c0001c0d000700cc0c4fd3300001c700d0400f10c000004400c0f343c4c05400c00111f3070000000003cc4cd10400010340004340c00000c004c0733000030470000cc4d00401400c0057c04070003004144000d01d30c0c3fc407c0cc04300573d000100110c0000440f001010000004410d00000030004300030ff00d0000100c003001000c470000000300414c5004c10000400000c000000071431000034001c004c0430710001d70c040444c340f700003040000000cc400dc040400c0000c40104005004f3c40c000c01400001c34c50730c1044700040000c0000c05c0000d3040cc7d00c740c4cc00f00343000c0301000d344000400010f4c00305c5034f400c00004050430d3101470f00000044cc0dd00040171c474001104d07d00700000300300d4054cd7c44000007001f0045c0c7140000003003c30c0414000c0c0100d4c000c04c0310c0070050d3404c0344f437c4c0000303c0430003000104000004cccc0f01c4570143044d1d3044300c00c40000c4cd00030000030700cc000fd1c144004000c104cc3000c4000440014cc030403c004c040040440300c00c0300c00004;
rom_uints[538] = 8192'h400c000405c013400000c1000c40c71100000000001001c130c10040c0130c0100003c00444000c001000304c0701f30cd00c00004103043304300f1004c1d130000000000004534000454c350001030131040044000134000330f04c10d00044f3c03400c7000000dff4c01c300c040d000f010f000000140000000c0300500000dd000000044000000000100c0003f343000f0070000f7400300000c0cc0f01304c0034001074001000000003030100cc340000007130c000000005dc000000130470c00010300410000403304505001cc114c001c3001000c1474000000000730000301cc40140d50045c4300750000404053103004001104030034400143c34014c000d00330000410004c500c1000d4c0d003c03103730010341333505000340003000004104f0410c3c0c1dc4000dd3110100c000000000005055c400ccd4054000c07000c1c3307c00000034001101013c501c0310100c0cc0001f333000001f0340010cc01c4040700100c5000404000c00030500c0000c00103000c0354f00c0040c001d0000030d01001000004003000c301c430040c00040c0047470c3001c0400004c0d400d05040403d0000c41d3305500c500c00000310400400004010f00704510c00c04040001c050000000c0000033000010c1c400014000cc4030110404000cd30014441c4501c044000c00037040c044000044c0001dc4001f411cc10001c4001d0010d43400d0c00f41300c341010cc77070400c33103000000010c0f00000315001d003400040c00300015000c003140001c00010f00030010400d013000010c1013010c040000400c0000051000000c3d0c0c001f1005550c140010010c1013000000003d00303c0040040405f044c0003cc000000000700c0c034c1001013d01450c41000100cd0c4fc3000300041f000701030300030c01cc00c007140c0305130010100f0c4d401c35cc05003d0d01044c000f0141444000000000100f00c41001000100c00c00d001311cccf50c03c54407100000110000f5000101001d0300303f01c0c000f0040030300110103000130300440c100c03003037c000000100001c00000100c0440000c00c134040710040c03410703010d00430104c340003340f04004000c30100c0c101430c0c00cd00000511000ff7040c00330010034301d310000c01c000070303100043000d0c03000103d00cc17f00f000c030f0c70040003100100040031033c000000000003000c34104000c0030314134005030000034c7c004d0031c00011d01c01c34cc00c30410041f40cc0c041030000034003404004c5531c000dc31001100000003fc004101cc0003100000c0003400014000d4040c05030000140cc00100104fc00d050010000c00001013000000011040d0000c1000dc000334170440004f03000100;
rom_uints[539] = 8192'h304310010030440c0d300307040000003070004c011c000031003000f00000004000341044401c000040c0000000c004710003c00041014010003d0cf00000000001c0001c34000000000030000c30004003010030000c0000000c1000314030c0301140400c070000103000301c0010f003041000100000010030550000303100c0c0030000000010000c00300000c100000000010c00003000314c00000330101000003030077000c4014001f0301100000000030c0000004000340001001000000000000000050000044010d1001103310030000430410303103031100411140000030001000000000cc130010030c01404014000003140300101000001000000000c0fc0300010114300040007000010044000000c00000000303c3004004001300031000000f31003005330030000c00103400003000300413070030000c001c00c1011000000c441c0510000c00400c004500000003004d31000400530c0040d3144101000034000c411003000f0140000100c04c004001133000030c04330004033004005000000fc030110000000003c10000103400000d001d000001740c0c10000c00041000010047100000cc30c00330140100100c0f010011001300400c00300040401c4000150030001c10300004cc44140000331000c0c140040303700003000400303f04ccc000c04000c000340000033c00000c1c300d00000003031000010140cf04000030000c00000010c014300047cc40410010400100010010100003300000010000c0100003300100404030c4510c340001000311340c010010003f0010430000c00000001000000100101000001030100000030fc00c0000cf00c0cc34034410031043c5010c0100000330300c0301100000000000400113000030000000013130c410000c040000000300400070c0100000000040cf001704c00f000013031300030030001c04003010001f000d1700001014010400fc0000001300c01010000003010700411401000101d7000300130304300003000000d040001000000440034d00014701344d4040d00000301104000401005001001000030011c003001100000000c00c01000140c33c000000041000030300c00000030c0000c0100130100004000030305c07430000c34301300c000c00430003001f030031000c030303c3003101000000004030fc000300000010100001044cc1103000c000000035c000030155c00c10310cc01c11300003c03140000330330114000c13040000300c03c310530f0f00000001004400000130d10003030000030400110000030000000c0000000300000000004300c01c001010000404c00c03031104000100010340010000110010000300003f00351f30037000030001031044d300100001400400c0c000c0000000100000003003101300001000;
rom_uints[540] = 8192'h3300140010000cd1003073dcc0001000400030c0100c000d170003400f1310c1cc0001050070c04400c000c00f003d31c0f0403101f7001c00005f00001000c0c3004000040050003c330c0030d304300c004c01c030f000034f04f0007000000dc01000cc00004c0000dc4300000370300c1430130c00ccf0001000c000cc01f100000000c000000304d00000000000000000000334400cfc4c0c400300c04300f4040c4000000001050030300c4000040000000404301330031001c00000300010000f0cc0c0340010040000033014c0c30010c10010f0f00030400010300003300110000000d30037c10030d0400013330004000041100030004000000d105cc0f000c005d04304000ccc0000040100cc3000ccc00133cdc04c050040c0000000300000030150c0c300015010110c00000cc30001c30110100dc00c00d0011034344d0c0000ccc114710d004170010004c0c000c443ccc03037c0403101104033100c300c0003000c000000100040000d400f1100000003d003f1c341c034030c0000c000000300003f0000000c10000000300000c4f0305cf34000000110c000f3000300000d00c401c100000154c00033c10441c1000300440c40c00c031c03740c000000c3c03000c3000110007731700001c0000707d0c0c3000c340c00001f0134403034c40d400340000030310003700ccc0003000330c0300c03330c0c40000004001c0040f05c30100c00c501004000001c0c0d07030300003100c0c040410307040071c00100010001c30000001400011000030000000dc30c144710ff01300300007dcc004c00504030100c0c010fc343d1f0344000c71c03501003dcc40c0000300cd0100500cd3030c04000f3001cf0000100040d100300f10000030c330c0c400c03d4004c0073040100000150003053c040cc00c0c3c0000300f000c40014c30001c4430041f3c7d00003030310c04c4c0c0f0330c04000000000000d010c04010000f030fc0110c114c10c00c73d0041070403f104300040000cc0070d10c10400313704703c01dcc00f500d000c30140d0300000041000500013130050000004400000000043000000001101000d3c007c000f00330100000340410c1404100301000030430400400517340004cc0000001c103000c07cc400300000100000000300000000030033003400c4030c400000d300c07730300c000030001c0c00c100d03007cc5c0cc014010f003701c00c000c01dc7000403310000c0011500000013c01c001401c000000354001000c30010c10000c0700011c10c17470000c0c0000300d000c0c0300d000000c310c000300000041030f400c1301cc70c0040c0000100d000c00004030300f33000500040003040301003000d0c000c0001100000dc0c4000f003030000c3300051c03f000c4300;
rom_uints[541] = 8192'h400000000040030700301030040c003033000400010c000c0330c00c0c0000000c0010030330000000c00404000000c4301cf01c70330037c004300d0000000000000000000000c000000c3c3000003000745030103dc41000410d4030433030040400003c0000c00000003000001c000030330000300000700000d110403c3310d0c100f00000100040000000044054003000000c00c0000c000000101504c000001c0000001c003cc00000011000000004101000000000030001301c000003043010000000400cf003004300303c0000000c400c7c40333f000c0000133010300000c05100000000000c70000c34000000000001000000300c0300005000005140001004000570000004f00c3000f01000003037030000c000137c0c1000003c0300000ff07000000c703003c00c30003000000400400000000004537034d1dc0110103000f0301c0c00d0003444003c00740000705030301c00003030301003003010c00311000130300c1c0000000031f03000014043000c104000003013100044000300003c00300050001031001000100c0010000010d00c040000c40040000004cc400010003330040f1130005034f010003c3cf0000001000033007030131cc004f000004c50300c000c00104000000400404c0030100000403000c0010c0f1017101c000c700c3307f04000303004050c0030300030100f001000004030400410001004c01c00000040304433400003300040c334c010004300000010340030040014000000000030300040440c400000030404013000000000300c3c50c00300000c30143003000c30000c00040c005000000cc0301300f03404c07000001140140c000000303010103010c00030000d0010001c4410c0401004000050030c0400000000003000440100c1703c301000c00010030404007c0000ccc0f00c300004c05030c0000300400030f01000f000300030000300300000400000005040000000cc3000000104000030003031001001c1c00030c05034000174c000503c00003000000c1000103000000030011000100000114000001403103010105030300004c13010003010043040d100104073000000d140017c003c1000001001300000000010100c000000004000c0c044c00010c03c50004000c00000000005f0000000f0000030001005040c040c0051005401433c100004000030330401001c00000400101000005000000310003c00400040001010000c031000000004000010000c3400000000cc00c40010004cc0000040000130300c00000030340334003100000003304003500000c03740001c00000000003c100001543cc00030f0c0000040100400043000d00343001000300c3003c030407c10300001400000003c0034004c100010000000c330c00000000430100005cc00000000000;
rom_uints[542] = 8192'h134000004100c0400d30000400373400503d000c3010c01001c1400040300004003c77534100f3030c00030000001c304c0c00c0cc144f0001040010000000000000007000c00010000010101000c0000000040300010105130413c000c00013100010004d3014f10005410030105c000030003c0007404c00100c00300030005c13501004c00c00117000001017c0c00300003000400400035000401017130470dcc00d001dc0103000000400c004c003005c000004d00f104cd10d0003034430c000400000000030000100040043000300311441400400c00c10300f0000011400003303f0000400404cc11d003014000c300010000000000100001000003004130000031073c1503c0d041f4001000000040004004001010070d3041c00104004100034701001301045fc7d0c10c000004010c0d0300c3000001400003d11037404000f0cc030000031030000000000c03f01cd410310fc0000701031000410440031407c00000100050c00400000000004000404000c331410100400300000047c0d40d030000000400740030c00c0000f33101d00100410470040300103013004c30000cc00000f00001c10100004700100c0d040370433000004000c10010c0010305403000700100330300c040000303300003d300000300003c0d501013010001c4010110330355c3013000cc03c0404000000000cc0300d10035c0fcc0c005010401c0003000c11f0004000100400c040000004000014040c10544cc1100004000c000000f31311400c0000c100000000000c0040000c0c000c00034cc4001c0050300004dd34f00f3003004403300f300c101700004400c0040000134130000c30500003307070001c0000000734000ccc030c050f301d0040000400c0334300400000000000d31000ff44740f3c00000300700030400010c001cd00004d01000c0010cdc7011c0400000140340c0700000c1c00403000700c30000000d0cc3003107040000c000050000d5104140100cc0c4cd400003c0cc01c040000000030000d400c00cd01001030300301700c00000000000cc01000c00c0c100014403030c40030000014000000c015d101007033700000430100000031343cf00000001040074000c40000003000c00000107300001070001730000c00103100400cf00003c00c11c00ff040004040004c00034400010c10000c00cdf3300100c03c30c044c1cc000001000000010cc00104c0000001f0330c030050043c000d0c044000010004511310003d00141154100c43d00001000c13d3c0133c0030c0004113001c040104400303300070035c041f0000dc0400701000100c40410c10110001107f00404010003f101c0003d050000c0c0c0c00000c00301000001000000001c04043400cf0003000500c00003004403370c03400004c0050000;
rom_uints[543] = 8192'h400100040500140370000101400404010030334dcc0c000300c340000c0c400000033cc314400000c070cd100c0d4d0003000d0000000c40004300013000000000004f00c1c001710001003f030c030743033c0c50c0ccc0f3030c04400314000040c1000c014004c404000c10504100000c004000004c4440c03c40047030c007430000400000dc0c0040c00040007c03400c000303040c3043000f14053001c101000300d344000cc0c0000c30c00000001040000f450140430000c003000300c0c40c0c07400c00d00104c00c0c01000304c04000c303070c03400103000334414f0c000000000c000c44f1f30000303f0c00400000000007000000400300c43104000f4004000c000310000040c3c10000000100000440c3000000001f000004300300450104040007000003d003030c0003c0000c00000c00003301c00c4303440000c0f0cc0c00c040040c40110301030d000441034401dd00cf04c000010004044000000334400303000003c0000510030c044100010cc50040000100033d4073c0004c0007004030000c000c43004041100300000c4000000100044400c3004044c000c00f03040000030103001100c503005104c000c440c10c001030000040704d0340400040030000c00354000ccc00043cc0070c030000c0cc4501040003c1004004000500415040410300c00cc400000001000040004300003d4000c034c1000cc00050c003014030c00034000f4401004d404440c0cc0d00c00000030f004000000000000310c073000513400003000c01d0c40143700304cc0404050300c0030c0403cf000f00404cc40400440c0f000c03c000000c00014000c40000430001410f4004007000004c0000000d00033010f03c0400700440c0030300104000415f03000004014300000c50004c00444000004740000300300700c1010001000343130033c4c44400c4010047000c01004030c0c330030000cc00001000000100000003c1000300c44c0543104400000040c0000730010030030000030c034003000037130401000c010cc30100c0000000050c040300330000400400300000001f1cc00000400000001000c000300040000c0000c3003400000c000c00000400cc03000003003c41000000d00f03c0000305744040000000000300c0d003500000c13400030004c103c00001300c0344433403000cc7030c00310530300000000cc000000470040d0404033000004d00030040c301000303cc504000010c000000003000000004430c1400000043405003030330030000400000c7c040000c010300010003000000500c0004013000cc0dc04c0000010000004c01000000cd044000cc050041cc0000330c00c000410040300013c400030400700040071000000000300000034040000000030303c034c034503c400000000;
rom_uints[544] = 8192'hc03400014c04000d04000100004000003700ccc0400030c400440000004d0c01000c0c0d00c100cc04300041014000c30303c0c040c00300c0300000030003000007010300010001410000003c0001430c04300000000c0340070c4000000000c01101000000004104c0030c000101c00000c300340cc440000050fc43143100c004040c30c000d4075000034000004000f0000400cc04503c000000000000310040000c0000310c000c0000d30c000c000dc0000000000d0c0000c0fc00034000050000000000c00cf30c1c303133400c000f03004013c3000c0f0f000f000000070004000010100030005d0401f1040ff00304c101000000c0c0100c3004c74c001000000040010730cd04c3400c031405c000300c0fc400040300110f03010133cf00300c41510c4410004d010000000c00400000c10000c0c000040000c04c0ccf010003c000700c001000c10000303f000440040400000d4000000c0000000c00013f010d03c33000030c000000030c0440070033d03c40050c4f004d0040000c00c0003000003300400000030103000c0300000f000400400300030c0701010d00040040000c000c0000400000c3030040c003000c0000000101d30000c0cf00003d4d000000550440c300000cc0000c00034073030000003000030403c4003100c330f0c70c000d400401070003004100040403c30003043000000004000044cfc507c00c040c0c00cf3700000010cc03c100030004010700301d45030030043cc03c00000000cf00010051141014c000000300c00fc0c000000c0c1d070300003103c00000034003400300004000fc0c001303c300400d0c010c003d000300040300000d40000300000c00000c033f040101c00c00c3050c10400400000003010000010400f01c00c001d0c0000c0f00004001040000040000030000370c000c0000f040000300030c00c000440d0440c1000000d00001c3030004000000400000004d00000000003004c30c004443c400403c03304000c4000d43000c0004c0010c01c0000304c0cc010000000004045700000440000000030400000c00100100000003cc00c003000dc1034107c4431000c0000000010c000f0d00030f0c001100000404c3000c03c00d0031004c410003000c4301c40000c0100140c00000cc030c01c04043000d00030400300cc001000413c70d730c0000000c00000011000440c3c14000000c0033000000cf000c0d4c0000040001cc034303c10c044000000440030500403dc000044cc00c0c40c450031c1c3d01000000000c000d04c300c000c400000d0000000300034c0103001030010100000001c0cc30451100040300c5440403400101000003000f0001300d70c300dd400c0013100c00c400010105430cc700c004c331ccf300000000000d004c0700000cc44104;
rom_uints[545] = 8192'h1000000000100004041c000403040c00040010cc10c001000007fc010370000000c0010004000000cc000c30f00c003044040101570c0133c0c0304c000c0000100c0001000d00100001c0100003000100000c0130000c000040cc000c010000000400004000c14010040000004000504000c030033c0f4000000000c040c00f00030030000004d00000400003000030000000c000001000000000100c003004c04400140cc00400000001001cc0000000114000000330003300000c0c0000400c31040000040c00000007100301c1140000f044003000000000400400500010030040000004000000040d000c403000304300400410000000000010700001c0001000c00c00440030004c000000030030100cc00000003004000cc00740d400c40330000000c001004d00174c0000071003c0030c0c000c0000140411cc0000000014003c30000c003c00000014003c00c11c700c31403330070300070000000403040c300000c00034000403c0fc003c0c40003c0701000c4004000000004310c010c0f0004000000004000000c0c0300000000000010043040104110f030c0000c000000003000c34c4004500000000000f3003c00313031c000100000f0c00000140003010f001040001d000cc0010000c003c0c00000400cc000cc0400000000c0c0000043030c40c01000c0c0000300c70004000c00c0040300040c30114004c0000c0c0c00100004000400c00c0040c00c00000010333030c444c7000004400004030000000000000000000005700c000001007500c0000040000030030400c3c0c000000000100040dc0400040000c00007d100000100000c0c7303000f0100ccc3030003001c00c00000c00003000331c01001107100c070000000000040000c000400c07034f0010041035004cf0c04004100004f0310d3015000ccc0440400ccf3004001000c44040c10773001000fd10000000c000c003000040010034c00000040041100c0000000c000073350400100000030004f100103c00000000000004000dc00d0004140040c0000000c10000c300400d000330d03000000000c0c00003000000000000300100403000050000000000004000000010c03000000c0c700310d040c40003044430047f30000140000c37000410044c300000f0c00c000000300000004410000000300510000050053c0404000c4000004c0300c30c0310003410400000000400030000000000000c0000c00000004300000c0c00040000000300000070401311044410000400004003d00c000c0030014400000c0000100400300040d010000103040030105000c0041000c000044030030c0040000030c00000000c01100000010400000003300040c304570100000100cc00c00000000c0404c00c30001cc03cc0000c0c3c0c300c740031040c04000;
rom_uints[546] = 8192'h70cd4040100000c040300d0001000430304c400003100000014010040011d00003c400c00c00100000000000d00010000000c00c0c301df1303000c340c000001304d3c04000010c00003f0030000000c01c34000c0300300c04c0030c101c00000c0010003c00f3000fd0000010003004400c00000030c00c40c010d170c00003030c00000000d003c113000000000000000000001040d000c00004c003000070401300003c1003000100003030301c503010000d001000003000374030000033100010000c1000300c0c104053c400003030003011c0c05030043cc000c0000000033cc5f01000c40000400c0c7000100040000000400000000cc0f00000001001000101c40040010c00000100c13d00400c000040041300000000031000c003c3000150030000300030f0000034307c3d0010003000003034f0ccf0003737c4c01010cc40300004040c1c0030104001c00cc040d013010000103007c0c00c104003130d000047c30c13f000000000c000f07040500100c07010100000300000131003d00000c040100014010c431150010340000170000010f004000041000030c0c30004c11001f040004040137001f0013300101044370000d0004c0000c30003cc41c030000c0010000000000000d4044c0001100000d430300340000c1000c1300300c05000003104c00000c0000c700010c1300c730000005004000000c410001000500140310030000c10004c003003030400c130010031c0040000000c14c10c0004700300c0003007000000c40c0c303010c30c00034c00000310c001c004330000000df1000cc7300000041400c0c010001404f0c404040015001000000cf3000400400004400150f4350000000073c000000c03c00c100000c00010000030000040001001003003c3c0c404000070000fc00c10d4030004077310001010100300c40004c0440003c4000c53c01010f00000f00443301030d0303c0000101000010c00005040000000000300c3cc00300300340450f000004300d001c0000130003000003c0301000340000c4431003000010000c100c0cc00013c005404f010100c0000100000c00c30130000141000100004013300d1c0c3c00000031c0001f051530004040004001000003c400c000004d1cf0771301000c10030c0c3001c440034001000c413cc000c40dc403030000000cdd00040304430cc1004040c000c7011000000000000000c0040f00003f3cc410000030141400330000003c000310401040d5000c000f0c00110001000c00430f400043000003c70c0c0110000c040c000004c00000100031134c070000000cc001000c00c4000000c1c70cc0013c0f000100c00f000030c0010040cd1d0000c100cc0011c001001001030300c0c01d34034303000f00474c000c400300000c040100000c010c;
rom_uints[547] = 8192'h10000004d000000004c000d310c0c000000000300c0030004470000470410000070c1050170000c00c3011000c00001001400030440030000040000c300000000000030c44000000000000350000010c01400010340c000000057100040000000003000000c100fc0c4400000043c00033003cc00000010045d00001c044003000003000000000410300000c0100f440c1000000400c000c73007074003003103c04400000000000c0003000c0034004003c000000f4f0c00c000000400000001100c3000000001000010400000040004007000301030000010c7000c0000104040000000000000000000730010000014501000000000041000100010000301004cc000001cc0030c0040300d000103041c400003c130001cd00000040130d0000c000c14000c0000c000300004070100000c4000040003c0000000300000003c000c73003300030f00074030c07c10310330000110300d0c00003040304001103000331ccc04400c303cc50004000040c00010000c00040dc041000004030000304017000000000dc00c00c0030000100000c40000103c000d0010c000000000040c00c00000c00000000000005000c40cc00c0000000004330030000000000000c0400001101000414000000000c00000c010c00c30c0000000c00000cd00114c000014c71053000c300300400400f04c14c030000c03000300130000000000003350071000000401300003d333000400000010000000330071100100f41030000000c0d100000c0300100000c4000f4010000030000300000030700010700000100100040000fc00070074100000000400004030c00401000100000041c13100c030100000004001f00003000100100000100300c04c40430000040cc00030000040500000c41010c0401400c31403300010030000000030030300003400100c3300c0c70000c01d304000000c000004300003c0131070007704000c3c00013c000c0000044f010000000000000000003000000c0340c0004000000c5000000000007cc4001000f710000000303030000f01000000000003c00000300004001300cfc0300300003400070000c004100c031005000000030000400f0c0440030040000300000030000000000440000003c1440cc000030d00400c0000300413100c03000c0000000cc0033300000030300f000000000c0c0400000000c0c101007c430000001030000400000040c14f00000c000c00003300c100c01130000d03001030040000000c0400000014030fc0000ff0001003000fd0001050000030d000c1400000030000304000c0000000430001c00000000010000013401400004300003400300003000cc0c000000030304000000000c0000104000001030300030000003c0400447003c000c000003f003000cc000000401000001000000;
rom_uints[548] = 8192'hf1000040504110410030003c430003413513010000c40c01000340000403300100034043c0c3003053100043000c01c00514010c00000c0370000004c00000010400cc00100003f1c000034400000000000043d100c00000014003c740004433004030d0013031450d1100000100cc000003c00000000411d00103c0000dd007f00c000040c000c30005000000c0c00c033300030040733011000000050000004003030010f00300300003c3000333f030c3400000003004100040cdfc00100001001073001040001003c000c0c040c100003c01500073c110300001c000000f00400010c0c00000401400cc01c1133100000001000000000011f0010700000100c0010000014000010040c04300034104003003c0300c00034003c004010001c0d300004050400000000004400001c030004110c00003004330cc00c11103c001104100d4c00303040c0350030130130300d031413001030003030041030033000010100140c000f04d01c0030100000013014cf0000040000c3c00000000000f0044300000001335014040c001c000cc0000130400000040cf400400000031407d1400c103000d00f11344010f003331040f3343c300004004300314000cc00430c10013000304010001030404333c01c0140030c1c3c001c3010100c04c0c000013010000440110d400c110c1000100000350400000013cc30010c041000500430cf10030030310057010000d40d0dcc003001100c401000030704015014003ccc04104c0c110000017001c30004100431000011100c0033110000100ccc3710070011000003104000000001001000010000d0303010110d41040000000150000000cf101c10141433000005010c011010f0000c0014103f133030100000000330010c0000030041003041100c000c4c00010040500700050d1140030d3c3d00350000300010fc0003000003100304c043014000010110700c1c1543c3001300070003000c040010003004501000c010000004473c0010001c30011c3f004000030000c371000d03040133003030300304d01404100000100053101c000c0000110c4c3000300000010c00010047000300c0000c10400400000033001130043c003030040743300c00c40c0000000000033f3c10000001000010003c0450303c00040c00c0030001c010003301400003004fc1130c0c1c01410c0c10fc300000100403070000d4c001000010040c0430c000c3000000c0040000130010100c0003d0030043000c031310000003d010c0c0c10400f000001010003c301c0c00001040131100000034000130340004100450010c50000000715030004c0151001c3103343007d1f00000041041c00010000030001c70001c0000103140030100304000007300500403300c0c0fd0103c000400004c051300401101001300300;
rom_uints[549] = 8192'hc44070001c0c00000010000000001c005000c00070001000001030001030000000000300c01c04004404003c00007000c3000003410010400000004034300030104400c000000000040040d003000000c30030003010043443000000700000c040007000c30000000000130c0010331000c000c0400c04c000000c00700140000f13400000000033301400f00000304000d0000000500000c300d00000f000000031c50010f0c010c0000000c0f000300070c0000000001000f0003444000000000c000000d000330000001330000000100000c0d0c0000470500cf0c0051000000001000300000000301040c1c030c0f00000c0f040000000000000403000100001c0f000513c10cc031c4c000100003035c053430000f0307350c00001010000c300000300f00dc0c05010330310c1400c0010c0001010000040d0c3030010000000d0100000300101001004f003f4000010cc005003cc301053c000c000000000c0105000c004c0c000c013000c001000403000301c41003100dc000040003310c40040dcc00010f000c000c00013040000104000dc004c00f100c040000004c000c00000000000cc000c300040040100f0310000100003c0300000c04000c034315100f000c000430f0000000000f0400450100004470000000000400000100001307000105000170107cc0000c07000c00030d400100000704c030340dcc00000000070100100000100003010110010103000c34000100110000000c00000300030000000c0100050007300c03000401030c01c003000405000d00003100000c0cc0000000000c0003000343010000000300000000000000000300040000400303000000000c0301000001010303010031dcc41d30001d000000003300cc07000100400000130330c001004034004003003404040000030c010c100c300003010000c0000004040000c0c00403000503000010000101100011000000040c00001c03000f0004f000070004010001000000100f0f0003000c0c041000010000000c0104000330000000100d10c000000c3c330c040000010030070c00000c30000c030407000140000000030003303400030fc00004040c01110000000003000004010400000301070000000040000100010100c4000f01c01041000100040003003400034000000cc000040400030f01c30003130c400dc0000f0104004031310f130000000000010c0f300cc00cf40100030c0000000c00003c0000003001000330000003000000001700003400010cc310030c00013403003c00000100000c003c000c004c00410f41340003010100011d000000000000000001010000011003f00f000c00000053c40c0000000000010000000c010ccc1030000c00000110000c000000f1c470070c000f000340000003003000000c0003000000100;
rom_uints[550] = 8192'hc300000310f00700d350000537305457005300c00004300004140000c3100000101c00f1c010000003000030500301403d10c000431000000d0c0001c001c330c0010001331000010005104000031c034053100c30013111c400004cc00f3000c1c3010c000c0530003100f0cc4c0003001d00301c00f0030040100013073003001f10c04d700010054003103335f04c000100000c0044030300501c0700f004c00c1104300f0710d504c0003c3100c003330000000000f00c00003d31000103301000c0030000100003005c000140334013001c000000003f000043c0700003145001014110c00014300340040d04107c00440330103c40000d0404000000030003030043100331000310c1d7000331005014013d00000000f0000310330700f10000034440030000c000d05033050103030c4100340001010c0000d0c10000010300d004f30005040750c041051040447010d000010c03f700410134010000cc14531c7530c504fc33d104430300335000300c0030001030ff03000100050c14c1040334c00030f000000704000031400000310011c0400000053c04037000f000000cc03700c100301003301c440cfd0000110c100741d001c0d0300011d03c010300004000c001400000c0c000000340000000344013030400000c00c040000000000730140c3433157d03040f00404043ccc0c43030010300003f00c437101010f003103001cd01111cf00000000031300f0d00c007ff000110c1000000100010c04f00c04003003000004310000c0c00003040cf001c01131f40030d400101333001c3c000f407005c1300130c0000030000400030014300003f000f30311003031d0c31c030340041704030073fc1f0c307301400051000000004040001c00310000100c001100105f000303001330f03304315c003cc000154331c00c3043c00040d3703f000d3c10f0400404c410c43f4043303000051cc4001010000307100100330007000103000f0000000304c0014733c00f00413070350003f1005300304000014000c004c10c010010c0400450003330401c10003000ccc010c00310010f3014c100f0c000300c00f0c000c0000f3c0030700101f5100500c41c00000101010c00c10000040005000401c341c04fc0741044c000000c01053d114011005330000051030c01310c00c50300d0ccc1c0d013f0050003010000033f40cd001c00010100c3001300410071000133100f5010034003370f004f000c001d01d1000300c00000c0ccc501000c0c00000000d0010c000cc0401001000110010f10040003000001110155ccc0f10c00001f000f71013000000111c3040071315300d0400140003003c0c501cd0430040000c3003000310330f00030ff000033040400300001140000030c33c01f0030130300041054300304010c0000;
rom_uints[551] = 8192'h40010015d00400000510c0310300001c00010c40010c00c0050c13c0031000c0c1000300050000100000031303cc00d1370010300d0470c0000000100500c0000000000000400100000404000000010000004430010000000030c0100330c040cc0030c000007c4c300c000000dc4007c003734031cc0530f3c04140140700c040c00040f004c10030c100000440c00004003000f0c0c13fd00000d00f0000010c3030040c00c1000000404d00c00d000f50040003001403440003030c00c000c000c1c30000003010000100403404000000f400010c00303c4300001100003c100004500404040000003030c01003043074001040000040c40430000000000000dc00100ff000000f0004c000f00001400c01034c0cf0d00000c010dc44400050c00030000c5cc04c000d0c34c00c0330d0040ccc03001000040001050013000100c00030f44000c040c71340c10f5000000c0300000dfc0c041003cc000c0000003403003f44f0c0000004040000004000cc00131d0303d004010f0000c000000d03f4c30007c500001d100040d40c000000400005001400000c0004c00000fc430010c40074033001400010010f1000c00ddc30c4c400114003000004304040433700000000c0c0000040001c0340c0000f00c40c73014404030004130c1000700c0cc0040404000c00170310c00000ccc3104030f40c00103334000c0111000cc00700c040034001000113000700000000d0001044c003000140c0c000044c4000c1000303000300000300c40001d004000043000141c0c4004400340110000004004c00000400c0c0100300001c01000300cc04000030300c0000004300000030cc00030400c0c000f044c00c33d04c0300001c0d40c500300000c0c003000c34030000100003340001000503000730040130504c00c0c000c101c0c044004d00c10033007100cc0501c0001410040d34100300c00000c0c500c0c40103011000c4000c00cc000000000004fc0000c0100000f3c0c3400304c04000c001000c0001004030041f0030010000000040cc4000010030ccd040000300000070001550f0c10c000300034010c010010000000030c003040c000001c05300c0c00030003500401c4cc4000000c303100300040c00c40000cc11000c001c50000030c4c04000cc00001cc4d00003044c1d000550404000100f0c0003300c30004cc00043005104cd04000000c300c10d4000c0c000430140c01c0c0000000030040401300c0040003400d05c400cc74c10010500100000000000c30c00001000c35131d03041170000000c010000c00c000003040d000070501cc000011003000011d5c4cc400c047c0307d000400010000001700c003001000c01007d0330c5f0500400400013c0010034343000cf0043c00c00303f7f0c0cc4000037100000;
rom_uints[552] = 8192'h3c04000000001000410000004003c040010030c05030300003004000040100000010350f010000030000103000000c0003001001110474330100000000000100000c3000000000400000111001001f0100004303330c3c0f3000011d000000100c0000000400000c00c0100000300500040c100000010000003c0030c044100301041400000c0004010300000000014c043c000000300000cc043c004404f000c01f30c300c04300000134040040003cc031074400104004050000333010000000000107000074c1c0300000c3003000034df03030000001003c0001000100000c000001014d700000040011040c03000000000c000000000000003d00000000000000010c50000000c00410004030c01c4300100000000040c0000300c4003000000000003c10410040110000000c10c0703417303001001c000104ccc1003000c00041000cc0031003c0030000410013c000003014010400300d001134030101000004513c000cc0003031000004000000010c000011000c010c0705004c0c10c3000d04000000c030004000c010070000000300000c0011c0000004003307300f00540007403400f0100000011430d0104040400c000005040f030400000004c000401000000101010000c700c000f41003100010d0cc000c0400010f300c0000010030c40000001f430100100000030c1300000000cc1f000000030000c0040000cd0410040000500701103030401d0011c000001300005030500000000700001000c050300000000000000030000c1001000c0000c300004000c000010010000000310003c0034100000500400404030101041403000c1d304400000004103d003040c1000333c0c004003010013340034003030c0000005000040040cc00301100400100150000000c44030c01010530010000400130403100410000000300070fc0001001000300130401010c47130000040300700c00dc00100000000300500000000000000400f00010103004031040030f4010c00400000f400d1003000c0c00000c0c010c0300f10c04c3054140000040c0000c10c0000000c000001c10003000001000000000040c000000100000c00004000000400010000004c0010c000000400703340c010000004000000c04003000000104043041044c013300304003030c003c00c050040015c0010000cc037c0c41c0340c00030cc003c0001407000c000cc0f10000000000c00010100100040000031000000c30000303043300c400000700000403470031c300410003030440000c00310001000004001c034030003100000f00000000000000100000030000001000c00040c000c0001c500100c3c445c0100c00c040000000040430040f330c1c000003c00000003000000000330001050c1c010c0000000300300010005c1f0c7c043000000000;
rom_uints[553] = 8192'h740c00000031410c05313c40140f01310410000fc0c4000041c0400000cc10000001cf1c0d010010f004104c0c1004400400740f0004040440f00c004303101000c04031dc00004400000cf00000140070d3017040dcf000100c3c1c0030110130440004104740400010050000400104c3fd000004001044000c40070041c0015d103010000000440c054030c00030000030040c00040000f30c0000014c03c00403130000d1c0400d0000f010005c001cc30330000cd4030044c43300d0001000cd000130003d13100c00000c004013000c0007000141f0100c1c000000003040417030d04c1100044000cf00300d0100c01c0013c000000000c000440000003c004000000410c1010c0005001340404c130fc00c04405070c3000d400313c0004c0d000c0000030004c374d004400cc013fcd3000c0400000c301004000004c43cd04000007104101c0130c001404c0d03d0040404531000c31304100035c100000c004013131033f4c00400c0d000000d400100d0c4174c110004100c000000005440040004c3000300040c30d1341c0004c00010001000cc5050100010403c35710004000400000350300000000c03400030f004030001003007104c101cfc044000c4100c00004c04c0c33014000000300c5300c0c40007301001d0144c00030300000030d033c4d000400c00311400cc4c30311000041340000f0c0d300c00100f01100c0710000570c4411c00c0334000c30000070000004000445000000000051f410300000000004d003000003430103040c0c4d4005c00c0000cfc304000030c0000000001103c0c00710400004c000c00004000350030310c407fc31c040040301070c7003c013cc000cc4c01c0cc040003001f0407c00741000470030003000130c17170d47070000440034071000044c4c500140c10300c100c0000044400f0740cc00730d4130340c100c004700000005070d0c074041000041d0104000000001cdc301c0c0004304000003c0000040f0033040c0004031c0c00000000c30000d0031c10000410000c01d1ccc1300013c054f05401300cc0044c041400710000003c00000c000c0034500cc00f0d0010344c044c0404004040cc1341c030044040107c1040c300700000ccc43c034100404c30303d0c0030300c040c053704c430410014004000300413000000030330400c10ff0ccc0cc4001f04c0000000c00c14c000003010d010c400cc00d0f3c44cd03110c40411000000c4350c00c001c003100003300c70000000d440040c1001040047003c5f0034ccd100701000000c010450c0c30c00100040104044000fc3f4c100001c000c00070c01470003c04c0c000041143000000300000c00103004c100c40000041010c000d04001c0d00f010000000c300c100f00300c4030300c7300300000035000;
rom_uints[554] = 8192'h43100c0330001f30004030fc30044000c4d000c430041700001fdccc03005c4d00cccc1c1000400001000c04c0d00c040000c0dd0cc3dc17144004003100000c300c431400130003000030041c00cc4c34070c00fccc0c000000400003000c000000c300100c0d170c037500500004303c0cccc03dcf10c0000c05c4000000001cd1040c040c000c000c0004cc00400010000000000ccc000000cc00000004001017530014f17f3103001007100030103c30040000c034c401100c144503100c040000c4300c1c040d3c00cc040403030fc14c301c10cc044f00004400040c31005103140000000330140000000c5c040c0140c31340000000104c00040000040000000100c40d07100c304030c001041044c4300003d000044000f100d000c04000000000330cc010c040000c30cc144030cd0ccf34000030001cd0f3544001000001000400303304cd305ff31300000dc7ccc0030c10c430cc0c040410300d300cc00040f3370dc5d70040401c50140003150003031004c0c003003300c100340000015300cc0073040f0c00c00c100100000000003f0c0d000c0c0140001030d4000c13000413000cc0370cc1040c0004cc00f100530c300404000030000c004c0c04000004400c44010043300c01000c05000404d74c00f70010350c001c007003c40c4c30cc00f1ff1001000c0c3c000003400c00401300100d33130c30430000000c000c04c500c00503d5100030d3000c003000040c0001300c100cd00300d440003c50001000c4040f14010c0c01040000170cf0005c00100400404c00140c00c10c400017c00300001cc000c000541030cc4103040030010c470c01101c00051d500175c0040010d000040040044c34335433c000700000131c00000c00c430400cccd400013f34141007010004700400c00c0000c0d1000d03003040000c333c40c5c1000fcc00100040000040040000300c04dc331c4033000c3000c034030c00c0103003000c0c4100f0000400300cc3f40c0c10c510000000001c00c0041f00333c00d400040000003c3c0c1c34c0d00000c00cc70c1c01030c430403000d0c00000000300f003c040304001000cc10000444151073000000400000000f30011410033c00f13c04141000c1403d100040040001001400c400050d50011c0c0330130cdd40d4004005c4003047310c0301050cf000000070cf07001000cc0c1040050c000cd0110030ccc00c303cfc00004d0c0f00d0401410007000100ccc004c0c540103f0040441041d0c0000cc310000d00000c0040cc0004c007c1000000c470003c0340dc000c30010003001004007f005cc0005100314003c3c01003c101500c1000003310c3d0000c000000c041003c30c000c30070004044000030d011c00304004001501000000c000440c000014150005010c3000;
rom_uints[555] = 8192'h4041c000033010077c0000000f54c3c00003700c0400704330774001434c0000300050000001001c03f01004110000c0341000001301701c004000010c01c00300033500007100330100c0c400000c10001301031040f040400000dc0cc100310031403003c04105304000003100300f00f0000010d100c40030c00700c00c3000044000004c0011010001454400040044c30100000cc040000000035c70c03510010c100000c0c00003404310c000304000010c0000d000c140003040440010013000d0000050040400001000000dd1c040f0000000003030cdd0051fc33310c301000001010330c031c0034f4001003040030043f00040403c3000010000c040040010044030c307d0c004f00000404dc3c00331c04003c00000cd40130c0000443000c004710000503ff00004410045c0540001330d0010005000c1c30400c00000001050cc0010000543010000c0c044401d040303d4fc031400033cc000000f04c0400c0c033000003400431100c00101307000440300150300307013011001dc044010000000310004000000030c0030c050100001f4000c000100c1403f0030000400015000000c004304033000000d10c0030330d000051300d30c01c30c400c1050c00000f4040000c303004374c100110153043000c004c0c00000103000400040dcc30013cf4003034040000c1053331000f037000100000031300001c0004303031c000011100000304cf070103004100400030034c0d000415101000030003101000000034000c00040500000004014013dc0001000c300c010000c3c0000405030403040700ff00103404040000100f0001003030031f0007d0000000070043003c04c00c30c1004010cf100c0300000000f0311000001c10000415310000030c34101f000c000c330c010c3c00110404000c073100303c0043333000d0000410050c4371451cc30f3d3105003c000405cd0000373133000c0000cd30110003000c00003000031c0f0003440dc00000d0f005000001034000341000000dfc4300000001000f03f0000000000f74441c110c10715434103430053c0030001330d140000ccccc000c0005c00000030743341100c5f3003d1c0300303000040d10050400000001434034cc000001540c04004fc04c03000c1d113304c0300c314cc010001000dd013c351c100c3d10c4300c04000500ccd0101f1000073330f00400100c001005c00000054100000c0f1c0d003400000400053c0c0d0f4130100004341c0011301000410150030003000d00c0100cc000000003c73c003033f1340f3c0030100101000000000c0033c40014c00f30000c1100000c411c704004034c00000c030c30000000313530340c001c1040d300c00c0304fc00303000300c341103c0000000337c0c100f03030300101c000c30010000343;
rom_uints[556] = 8192'h5010010010133340404c0000001033401c3c10c00d1004300040c30cc4c400100c013000300c3001cfd0c000f10cc4104d00040404015c0c014041110000c00030c0f4440010001103000c00c000c5c0f710010403010444110007f400ccfc04014073301013400001c010000000705004f000001013100c004400100d03f000501000040c3100c031c001003c000034700c10000010300000000400c004000040c4440440c0c31f07014c000c003030001c3f30000001000c0c00c7114500c10400330c30000cc000000001000000c414445c100010300c13d70d0c000110040c4cc30001000010301040d4001400300004c0c10c3300c01c04040c100000001400000c00c010000fc107100300c05000310000130c5c304703000005403000c00c0d00c0d030c44c110400f7000d010000400110040000c000007c4c001010c0400000110334001c003c04004c3c701c0c005c00cc00ccc004030d01017c00000300c340003400c334c010f0303500c0030c4300300c10000d3d030040f170c403310c04fcc000101300f001010170304013010c015001100110000000007c043030c0c30000040c1000004441d3d0075c0000c30c0000010000f43034c3000c1410c40000c0d030040400443001404c733330001d0d10003500d000c00c0000100470440000c0f0f0300d0c0c0530c4c03c00f330000540d001c04000311d0000f0044c00f000004000d000540f0430113d444c004cd3c000400d0dc0dc0507171005d1530100c000373030f00c00041474c0000c04101c44c134c40000cc0c400130c000c4004000c04c31c400005d0744100470d000c000000c04373d031741010043c34010dc00c00031c00301d00cc1ccc00310304414c000c340001030040dc00003040c105c10005c041700c40c441c101c030f000c3000040133c014c4c1c1c013300107d73c0c10d13501030001000cc0cc000000c14440700c011100010014000c40100000001010000040534d0000113cd0371030c3c0c00cc314003d00d41c00003040040040730c01404cc00c003d000400041c05141c1c0051000000403434403700000000000050c0f00cc400001c0030d304c00001003003c11000f7c000470033004303030470010c040010003010000301715c40003004340110040003011000d0707f17ff1c013c1034044400700300000000040f40c4000433140004510c00000040c10c0c400437004030c1c0310d00004047010c030c03003000304100000c010450100f010fc0100000c4000000c00ccc700073100dc4000000c03000004c400000004000c401043400c300041c00000130400110d1c41030010f0300100003104000030001100000dc00d0000f0003000000043301c0000d001c3c0c70c00001304fd0c4300c03004000001030f0c00cc0c104;
rom_uints[557] = 8192'hc0100000000c1043040c00004c400f400c0300c00c050000001014301c000000cc070000004f00000c003c0040000005d00000000c0c034c00000000c540c00004c00400400000c000007f4700000f0443c500c500100000c004c00400303300400000004000c40000d0c5030400c50000000cc4030c00c3c00043c000040100c470cf043400000000000000430cc004103300000000000400040c0404c4050000004044403cc40d00400c00c0000c001740000000100c004040000d00d4c00030000004000404004000001c0004403003c0c40040000c0000000c44cc004040340300400cc000000004400c0c01d00c04000c000700000c100000404000000307c00003cc0c40cc4c00044c0040000c04c001400000c0000310030031004340000000000c4c010d0000000300004000003010440c000400c40cc000030400033000040440000100c1007010010004000440000313710fc0c40c3304000300c4304c40c3f00c001000004c0000000310000001000300c031004c30001000044330054000370c0030c0000003000000000c0000440000004c04cc4c00000000c0300004030300001000070c4000000100c0040031001404d00000c0000001400144c00d0d107c700c00310c00d03000c04030040c00000c0c0040740000c0c0000c00003000c704c14041c010031400170c004000c00003000370000300c000d0004030040305004000c4000004cf40004d0f0000130005030c00000d340c0700000000000c0300474c0c3401003004000070000c030c0cc430c0000c00000000c00004300010c5000400300c004003000004000000000c00340100030000411014c7000cc50004040004000c0c00400004000cf0cc4d34044000070010c40040000001000140000c00040c300004c00031300000000c0c0d0010074000030700040c00000040c0000030000c033030000c141000043c4000c100ccc5000000c00c0000040000000c0c00000000070100000ccfc114300000cc000c400000000c04000030004c300c0004000000300004003c030043c30000000000c0c3104000000c000003000003c50014040c04000307000c00430000c00000400030000105000c0003304007004704f000000c00040c00034c00c30000040004000000440000f00004000001000c3000007030000330c000f00010c0050040000000000f4004df10c4c00c00c0030010c0000000c00c0c043040300cc0035400000c005000104000000c000c1c040000010400000c0003001040003000000c0000000c00000c0004000c0043540301000004000c10000c70c401004000001c000000001410003c0c400c0c0c400c01140c4c4c3000000300300004054304030c050440c4044c0c00000c0c0cc40004003004cc13000300004300000003410004700f000040;
rom_uints[558] = 8192'h40000000101310140010010300c4000410040000f00001500fd03000010400001301010414000000000101010000300f0344010103000014000c0000300031000c0150d030110000000000000010c0004c0303100cc130cc000000c400c040000330001100013000000f3000003d1000000001300000c00300d01100140000073410100300340700000000000000000c001001c0014c001010310004c0c000000c000c040c0c3400000004000500004000000000000004000d40050003000000000000000000041000100d1d05100c30c00d4300000000010c00014310000311411000007c30000010000d103100340040000c044010001000000140000004cc00000400710003c000101030040040004c13000c4c0100011000003000c505c00005000c100000000300100145304c0c03010070000000030004370c000cc03cc00050140730000c3004144300401030c0503041030000000001000c004010000000000030030030300000004004c0040030300c4130100075c100030003000fc4411100334030000000000c0500c401400000300000404003c01030c00030301000703003100c0041300f4044044007c000030000000003c4c0000c0000c00440340000015d00c301c00000000004f44000030c31000cc03030000003f030440c0410000004000073700001310000034000103003000c0004cc0c00104040000001004040300300040000c0303013f0007044000430000310303300001d4000c000100140310c0000c30004000000100003000c04000000000404c0000c00000034330500000010341c0c00000143003f0000300000004fc3044310000f05c10cc00010c400040f0c00034130000003000f03000004c000004100000100000003c0410030053101304c0c071f00100d00330000c10400c0000001030005000001fc0c0c000c45000c011000c10000001f300003300030000d000000000000000000000000001c000300013c0000031303073c00000000c0c000040c341000100000000cc003000004000000100003003000000000000001000c000cc00000001000000100000000c000030010001f00c000003340000000000000110070130013c14c044337000c00c0000300510000050300c03300140000100c000001401010005000cc0300000003000fd0c0303c100000c00001000034000000300c000000000000c01000314004300030001103d0000000000dc0fc3c0001404001f00004000004000000330013000c341130c0000c004c33003000400c1040303000fc3c03100000000d040001003000000c000c170000300ff00011c040043fc00c0000c005000300041001000001053000004103000000330c700000100400000c031000000d001000001c000000c404000300000000400c000030cc01104000000;
rom_uints[559] = 8192'h700d0000504105c0000c0c0c01010cc0c00000101000040c0010d4000cdc001000c300103300000c00000011400010c04c00000cc40c000014001300d0000c00040c033300033040070000d41c000c050ccc0c1300030d00030c04cc0c00cf0000345c00044400c004040700343c03050000000300cc001000d00c0300340000007c0c0000cc00431000000404000000000d00000000003c1000301000c3c3303100300001005300c30d000004c300c010c00000000051d01000000001030300000f3c4000004400003c0c30f0c0300ccc0700400411440000cc0c03133000000f0000000c400000005401c0001410000c50103d1000000000000400040c00040c1041007c0004c0dc0070f004010000040001030000c000004300f0001400cc000c300010cf000107000004c300000404d41404000c00c010004400400404304700504030100000c0000004f00000004000040100c11303cc003000000030000100d0c34014001004d05044004000040010000000115401c001f0000300100000040cd0d0100c00000010003000101f0f0400000000f030103c0c0100001c401330c4400c0000034000300040031cc01c50c000000f00404000130000004f00d403043d040300400cc33f000000c400c400100c53c30c0c100044010c0c000c100014000710c0100000000000d3003c0c0010c004000010c00c000c5340001d0c00c3101c031401011341010c040c10cc5013101300000041dc00410001c010304c0c0c570c04000000000030101f4c417c4400007c0070140000c00300001c00144c30c00414001400403c0f1c3c0000000430000000003030100000000c1c305400301400030010040010135000c3cc4c00cc00001040c04400001000703cc0c0000c000400f0000000f1050074ccd000c4cf40c340c0004400000c00cf0c544f01031003c0c034307050004004003010cc000000001c0000001000000000cc3004404500cc0300340c100000001000c0d0415001c003100003400100c4104f000000ccc0030c10000034400c000c00fc07fc0105100040100300100040c0d40050c03d031c400c50000000c00300c3c05000c00c0400040530033c415004000c0040010000000430001000d000c0c0500001004100c0040d4000100cc00000000053d400000010cc400c43000c00c03040d000750000cf0003000c0000001c40c030004100507ff010000000400c40000c000000030001000000051014003000c0000300340c4011300d0000440017470c044100d0004000100010c000c00000c004001011cf00000c005c01c01300303cc031000400000ff100400cd00040f13cc40040000c0d30040014300c033000000000cd000f00505104c05c3c140000043f040c00140c004000c400d3103c3030c000c0d040f14100c000000000;
rom_uints[560] = 8192'h300c004010c40110c00000730300401c0000c050030000c00001030410170000003005000c030013c400010001410030000000100100100003cd010340010103c000c000c000000000100000c0404000700040c3437f100340170c000010001c00013400001030130000003000c0400000c03c00000005000c0d000c0f400ccf00c0c10c0000cc0100000400001330c000001000040c0000040c01313101c0400041304011403c00c000004100000300004030000001c0114100c0f30c000004c4000000000300110000c10f000033000001003400040000034dc000010033110c0400014000010004001c3407404f00c3403001c000000000004100000000000500001041000f43010510c04431000154c000001c040070000033007411100001cc0030700010000f0100c10000033471c5043c01000040033000330c00000003040410011100444000440000000c1007000c0103003000404c0c0030030c0f00c000f70100400400000337050047c000000003000050040000400300000c0d000d4104040c010003000000001000010034010000ff00100c004030000c0513cf4443d73300c400000d0f0003000000030100000c000c00000300000c00335dc00041003000100cfc3001d0101f0007000000000005c4c00000003c01140100010003077c33004100404700d050c74000430001030071030c00001430134f0000c040c040000044c40030c0d3004000c04d0014f01c004011f03f1300000004001c04c1c004430000c000c500000031cc300003004001c00730000c00cd0000001300410c4c000d014000000400000400043c30010000004c354000c30d00c300000054ff10004030f30001000c0d30c3c000004001000400403101037c00003c1001400000c30410714004f0c5000000f005000014130040c00040000c0373007c0c0113030003c00330f40104d03000010f10403c4401040100c4100000c1c0003300000c00f00000010413007c0000010004300cc1c004100741500040c0000d10410c4c3100c10103301fc00c005fc3d030cc00000110f3013400c00004000104030400c10000000d000c0700c00070030000d0000400510001007030054030000100000430c00300000000004300c000010d0044000000f301040103004071c000000d400000cc003100500c0000003cc04c0003133030000000003100010004040000013040000000003010010c013100004000cc000030003040300c4c005000030000c013004030c5c0000003300340514000cc003001400100c0041040c0d1000013000c00403340000400d140100000414110140100000311c0034c03010100f74c101001010d1030000c0001c000000700c0410c0000030c0170c001000500103c00cc030000041400430000300010470003cc0cc004100010;
rom_uints[561] = 8192'hc00000c00000cc001010000101310c303f3c30030c4ccf00004c000000040c000030c7f00d71000010710030100003440f0040340d4301d00300000c4f1000000000030000000000000031c10c00400000000c04031f01d00341c000004000010004000f14000001d403010010301fc3030c0f1000030c30004c013140c11c000f00004c0043000400000cd30400000000c00000000000003403c0007043730004c00c100000053003c000030000000104000300000333003410013d301c00000c1f00400c00040000000010003110c003400004034000700000c00c0340c0000000001010130000003c00000010000000f0010c300000000c000031040d00300130040000040444000000010d0c30f04000030000000f00c110c00cc4430c40000f3000c1c001f030000000030100d000000413f0400040001c40400c01303000c030000431740c4304000000c00000040000403c45000c0cf03400300014000040000303000f4c0001f00004100c0000004110000010040000040404033003df0014f000f0003cf0300010c000000d000004d4000400033140010c0c30000c0d03004033c00007000000c00174010041000c05140000c00030df000304103c010300300010011c04300c000c000044030004000c00030001400100504c30010500013000c000300104071034300000100000004011010c0401003c01c0043001040000404d4010c00c30071c050100000c404cc010100001000400c0034700503c010c3000000304000c00c000350010140d0001000050c3c043000f00c0044001430100000000434c0000030c0300031031040c440004030034001f10003310003030d305cc03003441003404000037000f300cc400c01310000404000000004130000c10300c000f000040000c30404c00000030001000441f00011000005003040c0000c041c10c030000d0013003cc000030c0003134000c40000f0c00f00000c0040033c000030000000c000c14003c03c40c000c40000040000d03c030000f00ccf110000c000300101000000000000000450c00001403000c003003130004c00c0000000c000030c407000c4311300030003301000003100303c4301c03400001050c0010410044303404030005c0310c000000040000cf000f0000400000000010000030c10c4007004500cf00004003d04040000400004c0c0c071c0100370000000000030000410043010c04014000001f300710000d0000c00000310d0003000100110000000000010003c0041300001000003031000107000033c0c0011c0000c40c01010c010c40c0004d0003c300000c00f40400000ff0c000c013000000c30400000000f303010033074003000004010010103405000c04410740000103c04c04000c00000cc0500c00004f00001c10000d441400000400;
rom_uints[562] = 8192'h40d01003370c300413f000000c101c303100403014001100010100fcc115c0000430f111c1300c000f7011d00c0c07c00000010c1400c100010040000003003330d100c40130003000000c000040004c3034010030c0d00000c01310300c0040c0011c00c300d130000001150c370c30cc00004407030000300030d000700001f0f1d000040004300000000d30010d004000011000c000c010c34000010c0540101c300c000043000000004dc0000010000f00c000d03c0c013000300100001410000330100000cc04003004000100f001d3000030400001073cc33c0cdc04c040c03001c0cd40000d303d1c3074033511d1704003c0103c110c03004100003c1c00000d00c0033c40033500100340003313000c030100304500077031c000000c0400044004000f00f0f300000330041f4113040303000c100c01000331c33000cc1cc00f0400300c000d00140000c001f000c1403c40f0334c10d000300350c030434ff01000003c41301001040c000044c4000000c00c0100d00c30c073c71c40f0000300310c300300070300dcf100003030000000030103c31000d00100c03100110c3003100030304001030404c03000004040300c50000c3030000003740430001170d4300cc0000c3000d000040c7000c00cc4010130040f000c34443000130304cc0c00413340000040014110300cf03c00003010c004000000130c3033030000010000143330003c300c1c01100100c0100c00c010070030011007c0010d03030cc0300cd0000400003030330c30000c70c40fc010003000000c0fc0030303410000300c00340c00303030c1003000030f3000303040053030111100330001003401001000cc7c0000401000033300013330c10c0140403000030300c00000f00c030004030c40344440cf03f030000300ccd00041300cf000f304c0cc0c73100000003311310c00100440300430303040cc030c014033c310001000300000c000c000c34000000000c3403000100000300330103000400c0130313003c000d00003400100003000004010f000030c0000000300000011000300c3000f301433101000c044d010c4100c00c00143cc0000c00000000f0310034c0c0cf00000400001010001000300003104004d0cd0030003433c004001000040040100003000c0110010003c0103c00400c41f0c0150f00c111c30040000104001014c004300c1000040000c01d01030104f03003300000c10540000000001d0033c3030030000000100000001000c000d0000000f473f00033000300c0110000d0c10403000013010104c0010f00f0000043003003000000000c0c0030001110003c0c0100300110000133003001cc03cc000c130073003310000307c004040400030333004001030f1d0300000304040000040f1040d00c0f0130c3c7003000;
rom_uints[563] = 8192'h10010000000f4700c00100001300300c003d00000000003000000c000d003400000030000330000c0f300043040c0003001003003331000401033001c0040000010c3cc0300100000000000001000003000000333400030015040300000d0103101000000001010000003c3300337c00130000330500000000cc403000530f01f0004110041000050c0005400000130f3033000000010030f3300c0030000c0c000000003013310100100310100434400010070000004030330c030040000000f000001100010010000000300040351100000c000c0000fc30103000011500040140000005000100300001340000fc0000300000300000f0000c010d040400c3c00040013c30300c00044c000401000f0010000301300003100300040000fc000000f100c110104000040030400c01100001000d00003c001310010111031300c314040000030c011400033c1c00c11000030c0003300400c301031c1000c0001030401c11030c10c00c300010300000007004033103f000310f3c00003030004703050300c03001300400000100c040d000000010000f0c030030000400000c0000000c0310040f0001cc400301010000010074c30c003c33300c03030cc100000000cc0c001000301400030f030004300d000000d114003c000700000014c0400003d00034170c000303000433c13f00000300030000001c0004003cf30d311000f000300030000030cc500000350fc00c01003005000000001511d0000001000000010035000004030300030074c0005107000300300d04040c000f00450c3000013000011000300000000010013000001134043000000100000011100000340c00c030000c5401071300000000010c3c1300000030740001300000003000005000300000010000000c101700003f04100000c00c700701007300033c00010310010000c70c30f00430f1000000c033400c000300c0310c01fc0330010010010040110000000000c0000000000300001000100c15005133330000f0311000310000000100000100303004010000000000c04304040000000304300c00f0004010030414011c0510000f300013000340000c00304000000010040c31001100100000004c04050001300000040100030101044d00340000c074000130000010c0040000000000011045300303010351000001000000001430013100000c0030040c1cc0001000000c131000000111000000000d330007000003003000040400333000000100003000030000410034030030000030c053000f130300003c0003330c00370000101310000000033000c00015040f0c000cf0000f000030400c00004110110001003005000000004c0400300030000010011dc03c310010000000000000500401000400000300000333000003000100000c000400300000001000;
rom_uints[564] = 8192'h40c10030000c0f000f04003400000c00c00300000c040c04303040000000c0000070003c000300000c000070c001010f00000000000100c0030c00c007000004000c30300c0010000f000000004011d00c140003c030010000030c410c7003cc00c0c01c000030040054cc00000f10cc1040300000f0004000c0000000000000c0007c000c00000000300000000004011344007000040f00001c4004500043003400000000c0d0c4000030001040000010c0d00c0000000f0330000c0c00c030004004400c0000000010001c041c31050f3003000000103c0044d010400c00444c7000c00000000000cc001400cc000d315003003003000000010400030c000c305c00f40d1d000000c0000cc40140007040004000c0c0104c00000000cf0140330c3000000400000c040040400030000400c30001040c0010001c00440400000dc00c30403c0000000000cc0010f0400000c000d30000034000400000014c0f100c03004c3040440c1030c0040c10c00000400004c0100100cc0c00c00070700d100400000c000004040000010c304c00001000040001c040c0003130f3000003c33c0007000041007030c400c00030000040004010001030000f0c004cc0c75000c00d03004000f0040040004001000fcc000000000004004cc3040070c0300c000c0400c00c0f0047dc0404c3010000000fc34000443000003000c00c03330000070003004014c000000000dd34cd300c4300f0000101000040040000d400000c0000c0304400000001040010000001001c000004400100c00440cc003003000347c003040c00404d34f00cd03010000030000000c0fc0073c00043000c0f04440000300cc34000030400f00000000103440c1004003001510c00030300700c0110c00c00c000c330cc4000007c00045c00030040100300404704c00000c000000001003043404000001c0c400f413c03344300c100000004c00f00300030c004100000000000040000c0040040700c00fc4d00c500c00c00400f31cc0003c0000300c0000444000341c111c503011004c00104c300000100040000300000c4000c0400304cc30cc0504d00001c344100ccc000000000000000000c044030000040004c004000040c00400030c0000c401f03040000c040000077400c0000c50000000c0000470000010c100040040033340c000c004000407000000140c00100001000f10000000000031004c40100c10c0c3010c10cc0000000004010011c00c000c004c00040000000400404cc000c44100ccc0000304000030030000300010000cd0404500010001000f0000000c0c4007c000cc01000f00000030fc3010100304030c407001c010000cd00c00c0040300c000001004c014044000034001f0004c070103340031100400c03004300000c10400c00304040c300000c00;
rom_uints[565] = 8192'hc31000014403c00010000000004c4000410030000003c0c00000c0000100100000dd00701410000c0040000170000c443001c03c0043100440c0300070000c3050301300f00000c7100df33f3004f00d0100300000f0000000000fc00110000033c10c03300107c000c01000cc40000000303c0000303000004c00405131300f310000000110c40000004301100341000c03000000c1c00c0010300c0057041000d400c1343000c0c000000d30000c00000401000003c04c0f00010010000300c05000300010000004400c00004003fc700100c000304000c030030d0dc003400c000fc3001000000d400353c330c00100ccc0cfc0000040400003c000000010400c00304044f4003f050410c0000001000000000c035000003030cc40c01c000d000000037cc040c300000c000430030ff00c433000000044010004c0344033d001010003404000303000c03000103340c0c00000003031c0407040004050000001f000000c010110010330111c00050000400010c1040cc04000f0c0c03c0310700000d040000050c0014c0c0000001000c0340005f04043100000000400000ccc10330f04141003c130c300110000014700c344004140000cc1100171c4c0f4d030040c0004400073c000000340df00100104034743100c101070f3314000000103301cc0314003f13ffc30513c0030dc00004c43000c0030000dd030033014030070104010000c03400010000030c44030c0100047103c04040030431400404504004700c000000df003300010003101c0c00010050071c0004040000f3c0c0000004001c0d01141000c4334c03003100300100070000c30000700c1f04000400041c0000c00c3d00030300430f0104000074000000011c400cdf0c0000334c0704000000000010730ccf04d0c0c30003000000d40000130100f701c0003013037c300400c0100000310100310400100f0304330cc0c000c7030030000c04331f40000034000004000c0041043f043033051c03000c300000100f0041444000c0c0c431000000cd0030000c00300d00100c00000000c3307c044d071c03cc00100c300041111010c101c00400103c0c100c4c000410013dc0c000000c0040c40c003040000131000cc0c00000c10014f004300001004cd000000001300005fc00440030c0703000030000000400000000040010041100cc10000040400400040004c004c010140300cfcc000300300000000000003430dc001001030300043f400c0000040c4c0304134c0005c4d01f000c0304000440ccccf041cc031400070d3144004004000c00001000001c00050c100400300000140c000300c00400370730307f3000c003040330c000c0c0100001300000400c00d00010100003001740300070043f30010c00001f0544040000000d00fd010011c0000c0c0000;
rom_uints[566] = 8192'h10000000c414c0c0f0030400c40030f1d00300403c0100050c00c403c040040000103141ddc0000000c0c0010100400c041cc000040045440000c00d0c000000003030c14d10000c3000d0d013000000000113c01000001c0001001000401300cc133001000011340401030404c0c0000001404fd01000000000000330f3040003c33473c31c0310010401d3c0000000100c030000000004000000004ccf00700030340000005003f3000400000000004d1cc00000000c30cc04000000507c100000c10000003c000c000000000c4404000345430007c00053003dc000400000c0c0000404000000c00f000430c330c3c00043000000400000001000cc1000c0d0001c0010cc040071403404533c00044c300011404100001405005000004c000041000003401c03c0300000300050d04c400004c0003c0000000310dc007000700300c00c0d0c004130310000cd0150030000010044c4150c03c400c430c00c1040000003300013c0c0374400000470304000000000340c000000c0033030c041400d000301044300010c00000c407030000000300000007070041c0001000000f0c30404c00003001c4071003c303c0f00c00cc11c1003000100014001440d11000c300c03013d330040303dc0c00000c0f000df10000300f030700000300f0010f00c0c10d030c1c1004001c000004400001030014300400c04003430c000fc0114010cc00005714c3100001701010300c14cc300000350000004c0000030043d000c0000c01000700f104400100010c4c340074040400000410000000435410003003c001300c010140c04330000000c3c30000030000007c43dd300700fc0004000ff000c1444c00101400c5130cc00010340000c0100140010045c00041c04300c000000000f010010000f010301d43c034c0000040000f101c100003c740c010000031310007700300000c03004d400000030003000100010000cd10403010700000040000301003d03c7003300c401000cc30f104c004304013c0c04030010107cc043030310000010c4004101000430011c000010c45000c700003000000000c30400c000000c400003000013000004c1030003005030f4003cc0300400000cc403ff010d1013c00000f000003053c0401f13d03cc4000c104000c003040010000040c003030700030305c030410440030cc000501d03000030430c3000003c3c3000003000400004000300001000041c000130010c00000000104010c3f4030000c1000300100c404313c00010c000c0cc04000007c040000c00cc0c0100c0c000011000000010100c000000c03c35cc000df00100000000301c0314001004000cc03000014310003c00000000c00c000400c3010c0500c0000000140c0000c0c300100000100003040f100c010400f0033400c0443010f0000000;
rom_uints[567] = 8192'h3cc00000c0031d0040304030050503004000000130013c000000304000d14300033000740d10000000000334400004001000c00434300310000000030c0000033c0c503c0010300c00000f07000f0000c00f000c0303c0f1cd0000530050c3c400c5040300434000000340004003701f113c0c0403cf004c103010434010500c4c004c0010c00040c00000d0010000310003c00400303000c04c0030434141404030410007c307003c0f05c30003c0cc00c110c00000c04000000000dd0000430400000000404000070c00003cc003000340401003004ccc00f4c41000030000040300400003030000c0113310f003d103cc00170000000004000c04040c0013f0004007c0304001c403035010000700043c70034c0300d0c4100c0c70c00001400f0c001c0030c50300000030040f0c0c000017400504000c000c04ff00c0500300c4d7c0c510001f03cc0400000100331cc00c004104003c00170c1330334000c000431034010040001000c07340100000430000cc30c530040134000033f330053330d4130f000310000340000f1505004300040000400c01030013000cc501fc01034c0c01010003001000430400c00400c013031c33044c0000000443d0430001000700700c43410704cd003cc010c000cc0050cff00000500f03030003100000310043d004100fc0500100300f130c0f00403000c0000c0000c3c4300300d040c0000704d4d0050fc1c000c0d700c007f1c300000043030000c043403103c001c0335f101c000000000000fc43f403dc0000010c0cc0c10400010303473000005c1c004c3001c40f000030c00030001140f0c310000333003001010c103c0000007040004044144c030000104300000343c010040031cc3000040cc5000000334303403051330700104107c300430c74004340304400170000c3000cc00f3f30c03040400c004730d4141f11401004c000403000100030cf010000c0004000710c000000300c00c00030500c0410d0303004c40000f0c00c1000000003410040030f10300000040001000100000c03400d003c00c0000c00347100030c0000c4003cf0c00440c4104c000c00c03000c40730cd13c040100400c000001c00100000151044044c30c10000003cc10004000310c440c4c000003c000010000000cc0000000741004f0c040100000000000000030d00c4c01700400030c4030004003100000004c40000330000d70003005f300070130004000404010c51300000103c00107000d5010103010d03444730c0004401c4040c00100004cf40c3f4d310400303c01c10d00000040300c300dc103c000010000013000003f3c0d0004c0307ccc03cd40c000104000d00030c030101400c00000c100311040003041410000003f0004fd03c00110010dc00c00c00000c010f030304140c0c404000;
rom_uints[568] = 8192'hc000013c5000100c0cc7f04000503cc00000014510000040133c00100001003c00000440000000c1000304000c43030700c3c4000cc0003c5c003f01003400005d00011f010c030040034100300c00000011f400001f40001040001700004c0ff4410000000030010d00310c000130000f000fd0044d30331c0401fc1100fc0700000c0f000c0034004c4101c47f4000001000000f30000103000354015cc013000000cc40c3c000040004cc10c700c1000c00300f00100d00001c40000440c00430fc00c403100000341014014000fc0c004004003c0c0c0440040300c000000000c04c1005037100c7403c410c0c005f30003100000004100710000001c04000c04000ccc44004304000401001400f034010070000c051303f40f00d030d500000004000030004f0000001000040133c013403c100c0c00c0030050010110c50401403df030000040c0740001fc504c030400dc4300cc00f0c000100d101003311003045000005010c030001410c007c103c44700cc10c3000000001304314f4034100cc00040400000c000011c70c000004000c04c13130400cc4004c004dd50c01314000c0100304c0133100f030700c1034400c0c403c013400703304314014c000d031c0c4c0000100f3000030d503374034100010013cc000010c300010c3103dd50045140000d414303431400f03c3000300001300c0144140010400070c0400310000004c4d70330000010d0403c000004c4400303c043150040053105cc30c001f0044004cf0010100307f0d0034040050043ccc0431000041000304003c000003000c0030c0c51f00034154c00040c1000000014041003c0c404000cc4c4c0c1dc003340034004004543044f000100f305c4c00030c4403fd00f0f0400000c3f01c1400003003000c34310310000000cc001503053000d3104d0070000cc10c4340000c40000040c00c34000ccc0401400100f100c00f000300c430003000000000f100c0004c0c004c003c00313043000041030100004c001000f0000000440300030000000401140040c04f34304000370004c3001030401030000010f10c0400051101000c0034570001000411c10c00404005fc041311000000001c00300000ff4f0011501c00400001044000001700010100040c0300003010004c4013100c000d03c33d3df03000c500310f000c4c101000034303100400100130000010000000c540c303005300103034013113043f0000033000c000005d033000c000530f0000000c000c01405310310c04004c3000040010000300c0400c0c004511c000c300cc00c0000c00000d0f00100101000000c3c40010014000c00343f010000010fcfd1000f004100040000f1010007330cf00013001040d0104440000033c003001003014000701004051c00d00434104c010000000;
rom_uints[569] = 8192'hc0404003c0000000010c0033000031104030c0c00c0010000c04f043c00dc41440304f034074000001100c030000c000017000fcc030c033f0000044000000000000001000000010c0000cc1c0000000500000104014c010100fdc00000c00f100c0404040000047c00510000140010430000041303353c1000000cd0104c13053400c0700c0103000104010430071100000000000130001d31000c00000107000333010c040c0c00070001001c000c0003c4000000010f0000000010000100000c0004040007c01c00d005c03000300000c500010c40101c3c07040c001003d030000000c0001c0000000f00041000f001fd0034401000c00400000000d40c013101000d1513c047700003c00050010004444000344034031c000300010c0030003c000c33303000010400100000c5003c05010010010000100100000c100011300d04000d0c100004f00c0030401c0313c0030c37031c03430cf14000005004300c3301f000004c104100000d0000001004503300000530c0040000100000003004300f37030003004000050004000010000c3000030000000040040000000c35000000100000040000030004dc000011000100dc000d3c0003044001400400140003000300300403100000001300003001003000c00100400000001c000c0f0c3cc31100c0030301430100004000030c030100000300cc0004300000f400100c100010c440000131043003030c000000031c30c0000100000004153004040000c30500f0103000000f00400000004d3300c0410000cc100dc0031c100c0f1000330303003000004000040010400000000000cd001017044000c00c11000c00340c03001413110f0c0403000003000d7000330000000000000c030c430400040d00c10410000310c000040c100c0300d50000003c41c013000000040003004043c00330001000000c0101c4000d040413304f401000413000001104400000c00001000000001c000510073000000030c340c401110040000030101000300051300000f0001300fc0000010007004004430dcc40000c3d00040f000c30100000000c40003c00f0001400000000cf100c00043004000010000f300f10004f01100000000040110c030c0000c100011000000cc40133304000000011000104000000c00c300c004010770310030003d004010c0000010000000300c0100c0f0110000f031040d0000000030d000403c0107c000100001001010000000043010000000c0340c007d0013040010030d100c400000030003030000d0340000000000c30d00003450044430030dc40300000400400113c100040011010000407404c00040c0cc300f0c000001100003334071030d00000000d000c10400000100c400000001000000704000dc4300c0c00000f0000000000040004410700000000000;
rom_uints[570] = 8192'hc0000000c3c000000c001344f000001043c000300100004000430003f0100300000010100101000001000050540030003001005003f00c30410000000300000004000d00000000000c0000000300000100300040030300500c00110400c3000000f00cf0c00040c10000110404400010000040c101cc0033c040001010f00300001000300000005140000000300000703004005d000c300053c30000300c3cc03030303100f0300000010c003413000000c0c000003004004010c0000000000010001000030000000cc10000000001f5c000c0f000000000000000000300000c0000000000030c000001c0074d0030301003000410c00000400101100000003007300411503410000000111110000030014004c300f00000140c00300003004000000000c1c1005010010000000030c100d010c40100000033300c0030010001040000f300004000c0030fcc1300000000000000004100c000133f030030f01c010f00cc3001c00010300d00000000c0035003030000d70001010300c01000330000004053003c01c0300010c5004070500000000000000004f04030c00000401001010031000000004300f10050300c0000034400440503030300030030340110350400330c50f00403c000c00000000000005044c003c00f1000100300010541005130010004010001c0c7410054f00004040040cc40043310000050c4000700000010304000050000f00004404c30300004401100103403000000c4f005000000030000000010010131013000434003000dc0c0f40000c1330100c00000cf000000f0100000000040100003300c00c0f0010000003030010410d100300300001100400300003030003000000000501030c00c000010c000c40000f34000030300000c000017003050c00c0000400130f10000400c0c0c000040004f005001000000c00000005300f0103100c31d710ff4300000000033c000c330f00000f00000343010000300cc00034cc01000010000043000f0743000000003000030004d0030000300f04000000004c4000010f000000000100000040c3100430005004004040000c00c100f000001c1000000540000000000300300cf00c0c410d01100f3000040100cc03503400000033c000000c00001404030c010000000f30c010d04050003003300100c000c00305001d000c4000311504010c10c0070c03030100033000c0300040000000c4301301005000011013001dc000000003041100030010000c0000000704033450100410103c00f03305c0100000051040450003033c0c400400011000cc03000130000f3000cf000030001100c4001000000000000303f100001035000105030105d000cc01c0001c0c00001043cf00011c0373030300000000000430050c004000400c00000c030000000c003000d0c0c000040;
rom_uints[571] = 8192'h70700000000115010f01001000000c1c0100c0011c7f0cc30004010000000000c0c1004000040003c00c10101000004c30000014f00000310c00003c000000000003004dc301000450001c1d700003010070400040000000410c000300443d40003130000c00004c0040040430c3c0030300440500700c0034040014000300303010c400000c0040151000000f000405c0000010004004c0000f3c00030000c00c000000007f000104000001411c030340013300000000c3c001310ccc3103000f0400030000005001000001300000030000c030000000300040044004040000001d000111030400000000d50005ff0000044003c10000040004005d3c0700000500031d1054c0c10c0334100c0400010010000c03330103cc300400433700000c010f007c3c40d000430000010c000c00000030000030400003003047c30100000000310c30d4004fc00c000040430cc0c0000740c0333c00001500400c040300c041444010c040033000000000000c000001000700c0000f0304f030000c034d003c0c011c040c000000d00c00030140000303400033000030000c0000c00000404c05000000040341000003150f4030000700c00003044c10000310140403dd0004d700311070100004003c03c040c7000000404cc00c04c0dc000407031014c01c01000044340103f7701fc0003000300003c0c0000100100000010400c11100c401c714073011030341300410000004000ccc000000000001044004133c0000030c00d0003000030344030c0f000040c400000d0044300100cc340005f4703000f0004300403c14030043d0440030ff0c15403304000000000c30003003000300040000c0007c00030000c03c1040043004c4000000100100013300c30400401040040000d30d03f44004000f00177ccc41000c0034000c0000100040403c0f3000c4dc4c00000400400c0d0010f000010c00004030000033003f0300f400030003040030010303031000c10000000100000f000000033100003340410004004d00c001c111000300050105100c3c0041300004000000c0000004040c000104f40330043000000303d01001103c000100000000cfc04c03c703071c004cc001000c000041004300000c0c14000000000c144d0f00010c1010401030100c0d010c0000000c044004f103000014030c00000300c3054100340400030000004000c0c00010000003000040730044004c04000000004f000001000000c40003001d0051040014f000470c040003550000f000cd330144000040c0000010000300100007140004000330003cc70004f0005030134000010000000c00030000f001c4f40100003d10001405010110001400c00401003300701c43f0050003043000000000040000410440300c1104c100000000034c0c0c0c4000000d01030410;
rom_uints[572] = 8192'h40c0030000013010cc0000003010000130cd030050c104000040050000ccc0401034ccdc0040000c30c5005c0d0000cc100100130300040140c001c010000040403301050c04000033000300cc000400003cd1000cf0f010c0c000cc000f000003000c315003c153cf0000304030dd103100301434c100c0000f000400c10000c0000000000000440411400000003000000c003000110d00f0000010000000041001100100340000000000040000000000003000000034f00043000f33300000c0c70304000c000c10100c05c10010000c040004010c01f03000000cf00700040003000000400000101000450004d104f0100000400000000000040000000000f040010400300704c53300770413001000000000c0c11105f0f00c01300c3f0000003400c01c0000000040371100401013100c00c000c00000004f30040c04004011400004d100000311110030500000007c4030c0c4300001003033030104c003cd10001c0f3400350000000c00000000010011103c34430c00003034d00100300000004d00311430304001c400c3010000400014000f11f0c00c00c110000003001cc0c00004000c00301003144c30030000014103004011000030404030000000000030510c3000dc0000000000001c0041110fc001c0043400100400100000330400c000f000717445000cc0c3f1c400003530000300c0300000100c0100cc070500040f0003504c0101c4031c30000f000c0000300040c0030300400010c10030110ccc000c003c1304dd00c10000011c30000c3031510000511c0000cd003010041d0000030331000f344c104300301004c00c000440d051dc10011c0d00000000c430c01110410c0031000403030701cd00000f10003703040cc0470d0031004c3c10ccff00cc000f0300300001401100f01005c300000101c13011c10001003000001000000301f0f0300131000d301000000c3000103301010101c01ccf333031000010c030c0000000000000d40030c0300003000531f000170301c0000f00000300c3000c00c03404001300c0031c40000300430100001c3533001000001c1034f0500c000030000100000003003001100071000400f7030001000005030c0004100040010301100000000034003c034000101001f0cd13000101dcf011000030100030d104003000010011005c01c0030003000003030003111d300100c4d0000000000000100000040400000501c0010000c4000000731f0000c500140000000cc01000300cd00050340033310c0000000c40c030100000030114000101010c00300400c01003c0000000310430c000010401000000130c0000000000134100530410000304031000100000000314301070000070333730cc4010f000004000000c300c000007f010303331003011d014040040001010000000;
rom_uints[573] = 8192'h10300000004041300100400031001c101303000100000410034000031033f3400000f034cc10000000000031000005c3303000cf30f300c330c0000003013030c0405ccc0c003110500030100000f140303330450047300130031c3301301004013d01410500c01000030d003013400000500301001c0040004000031c14400040c04005003000030010014c0000104040d00c0100303070340131007000070330000101d03c1330010c403000c0001030f4cc0000030d00130d00103301f030000101c00000d0010030130100070c001035c030100300f0c3c00300311000cf40000000310004d00010013741410000000c0040c100000004c3c03c030000d0400140f000f000001cc0410c0000030001070100130f31040c000033c0c00cc10013000030034134004400004000c0033c3c0c0130c0c000c0300310ccd340171d00c00011040500000000100050040000f00001015017030003c700001c10003003705c003111030003031f03c1331000101001330cc1c003001000c100000001c031c000033300cc34010030000351300000c31000cc30cc0000133c033305c11d000003304130c0c33c0c001c3030fd03010c100c10033034030300444403cf01c0d03000c03030774010cc010c031300d001013010000cc100f30c0707cc0340fd31c004000000c00310501004031c003300310000c00000000003f30c30c00007c00007000100010007505304034f00cf3cc000000003000400000310c000d11c1dc000f3000000c0004c0075c00044cc0000c00001100c340030000333c304c4f0000034010000030f003710000145c000303c00004710013c01000c0000c0c0000000005471000003c03040300040030300043073110015000010000c00c130c000000040100300405001d000040010c3c03001400003501340c0301fc030100c01100c10c100004cc0000c10513030000c03030400000c450f030000000031003000704033cfc0300010003010400010033cc043003d330c070c40c400003000c0cf00030030ccc0c14003544140f3503000f30030011c010000330014030010103100353000000c00000011470103030010c3000003000030d1c01074c000cc34034000000300d10c00100100030d000c010003cd40c00dc1c0c0f00300c00100c0411000433100c5045300033cc0304105005001c0c00030003310310140c1000000030000000007000c000c00c13dc0001010030001cf0540000cf00353000000003c3040000011f00410c0103004c0000000ccc3c13030c3000030c03030010413100c700000f300000000c000100000010000043000001030040000443031330000000011c03010030000003000003000c000c07003c0033cc0000300400101000f30c00000400710101510000010003304334003401000c0c0;
rom_uints[574] = 8192'hc30000417c000110040000104100000030000000c03000000075c000f300400000cf4d304000401c0001415001c0d3000c00c301400440400040000300030c13000001030000000000c110f30010000c003030c431000000000103000300000c0100703d31000101000100301300001000004113c03000000030f03010c00c010003001003000300000000c00050c0000000000003c30104103000030004000003400004014c130000000000000003000000000001030000c000c07dc0c300c0000000c0000100714000010000010304000500000000003c1f0030c4d3010d000d00400000000000d00013c00d0000f000c04c00030000000000000c000004010001000010000404d00310001d0040134403410103f100c00d000307c00440000dc0000300c040000000c000c000000100310000001400000040000000053f073000001f330000000cf1040004001003310050400130000300c0003000000000c030070300c04000000000000ccc050400340003040011000100c040007cd04c1150003043400040c04400330c00f000000010040030700000000001c00300337dc400c030000400000c05001d0000000400df0303c0453000003000003000010311cf0001013101300000000000c03000400040c00030c0df000100c0c0010300f040000cdf03005d5f41c30000000000000f400100140000000003000cc000000d40000000004147100013c00000c307030cc44001005100310000404100041300cc1003d00c00c043014c00340003303000010400033030100c1300303400c300004030000cc0151330074441010040c01d0000000003000030c340004c00c1c000413100000000f00400000000100c40040011034000d00000c4314000000000500000001000000ccf030003c0474300c010000ccd000100000c04034c3100000010c0300004033000f00cc117003000001051000c0000300030400000000013030000400730400c000000000cc03070103400000c0030c701c041f140c000030007c14c0000000011c3000300000301c30d01c00000000011c40040000c003430c0c0dfc30000001403300034c300f0c031300030404010000310000040030030000100040007cc0004c4000000d00cc000000400c03100000003cccc01fc0500000d030000f00cdc0103c4d40041041000400407cd0300001f300300410000400c00000001100034f000c0004003033000000001510040000030010040000000400000c0000000131cc0300101c0c4f3c05003001000c04003000013010c0100000000000300004c0100003000531000440040c1000000000040000001100001000f010c000000000010004033130400000000d3c10000c0c0004340001040004000000000c7c1031003300000000c3100000000c1c0305034000000;
rom_uints[575] = 8192'h30001330100404000030c4003c130100004000101c000003c4005030340f0030c000000030301000004000000000043040000000000000300000010000001c30070000030cd0000030007000c04050000c000030100000343030301c0c3010003c001c003034000000000403001d0400300400700000300400007004040030c00000000000040410000c0000040004000000007000300c000004040400303000c40c14003000341000141c3c00400001030000143010000004040c0010000c00000000003400000100000c001c100331c31100000130003c10041c1d00000000001c073004000114130c101c0004700013000400001000100003003000040c00300004341103c00010400c103c10000000013c0030000c3f30ccc30c1054004c000000000000000000010003010040000010100040000001100000000c003731000000c0410130c030140c0000000040000010c0310c300c0000030031300000030030301000cc30000030004c10000000000030001030d0100010fc00001c430c40130430443c00000c0d00340400000010340040303f07000000300000001c040000011410000000041000300c0c00000c00540004300c3c0000003000003000000000033d00004300000000330000103030c015400010040001101050003010c01000000310ddd000354000405000000100000400c00c000014130c00c0000000c000001004341001000404003c0000f1430101140000c000c001c01430d000000030000000001114c000000010f0500c0004041c0100003c4000000c3010003100000430c01034300c103010c00004040000000000010400000030010ff0000c00000000003000000010010040c00c0004100c05101000000330340c00f00c100030000030300000dc0304100005031000003c30004c00000400cc0000000000000c010c5c0c3000c01c0000c000300040100c1313c000000030003000000004000001000c0c00000013000000300c500500003d0010000013100000c000f0001000000440031c0c00133000010c00c000f000000000001004000000510010303d0c03303000401000004100cc03000010170c000004d00000000c0003100003001c000030000330401000000000010044c07404301c000f00000cf0440001f4000030000000000031003d001030003010503001000100000040300c330c14003c000030001100304400f400d010001c0074100c030000001c00003040070300100034000400000c000000031cccc00c00030000110c130000040000000c01001400000c0000c1010000000300140010010010104c0000003100444010d0000c301000100c0013c04014000100000010000c1000000010304040000000110004011c0034003c00c0001404c00c000000343410310000001000001000;
rom_uints[576] = 8192'h71145045057040031000100330000cc353c410407430435c430d4341003cc0f003031c10000003000c7c0c0003040f00cf54cf004c01457c54000443c0303044c0000303003c3d30c00c313fc00430c0400001c0c0130543001c0cd1ccc0030000050174403f1304f04c4404104dd5440c4301c1304c31d413c03114510c1400c0100c3004cf40404f040537cf05f01003030f100f01f011010c00d0140340007c004c0350f5033030c3007040100000c04400000003c13c50300430f3533704110007c50000cf30c5001100c13037c430101030031c3407031043010c5000000000105014000300c5314f10f0110005107f7fdf45000000cc30004000f010f51c7140003cfcf1303f11130d303f33030030130fc4f1fc5013c00301f310310fc503100f304100c00f00445333c0c40f3034040303071000c0004514f0f4c0c4740c10303171d0030f10cd7054031cc40070000030fc731ff0cc00400c301c100f0114003fc070c5c073c4305403000140401c01d0f55030c4f405454010c4100144cc4c7000c0f43500010100004510c0c01c4300170050c7400ccc000cc01d07c0700c040003304f34c5010ff0c3050d0100f57000c410310400c0001c5c01ccf0c03cc700130f1c1f0004f505033430c10034401343310f5333043f10fcc040407f03ccd0d0414c01030c0000c014300d077101d007400c301c04401134000c0c5f1c7400750cf13000cc5f4f0c004c0f00fd0000100fc303441315104400003030300dcf000010400003400ccc3004010000c3343417004000d550000004f0c0100cccc0c41f3fc30411d443000003c00f0c30ff3c00417005350c34d4040c303fd0c0040ff37c4c003c5015c31f4500fc0f000dd4104c030404404013c100d45000003030000cd3007ffc007f03c40f30434f014400037c4403f303c033f0f430c501300fc7047707f0f57c3077cc03c03130704f3c34000c544000500fc3c350c0400c014005c303350010d1f573f3d01013cf0003043c005c70301033000cc13400341000403301c000413440011fc03c000300000445c0014cf0c0cc000505ff3fdf437df03103404c00700001403c00c304101000c00510d0707003c303400f30300130f05300003000000cdfd3ff047540114cc1d110cc413f00c3c0cc404447343c0f0c01c0df5030340f14013fc0f45cd0f7c4334003040f0d00c140001070c303cf10150c33c00310c0343d001000d34031c0c0c053c004c030c00c30401503c4303c4410d0cf3d3cffd0734044014cd343734fc00ccf00c00405340c33c0700010050403c0004ff05c0350cc43000000350530000f01110370c0713ccc43c1035034305f00c17301300440407d0430430010c00f750c5040335000301f33c57f1404c404334ffc04401c45c33007f47c0f00c340334140030;
rom_uints[577] = 8192'hc11000300000c304c10c00f1cc0143310400c00c410300300d10000c5f50000040001330114f30f333c3c70ff0004300103033fc05cd0c304100c104c31c047c00c40030ccc730000000313f1000cf307000cc000004000c0c303f04000070c001ddc40c300303070113c03d1004701001010c000f303530000344c045700000c474411003c3005030300301c00df3000000003003d301700d033c73140100530304400030c1007f000c030fc34001c005001000001fc17103030cf3d040c0301c700044430d00010c030150105070000c3000030f3d1f0d03101f1c0fc0c10c04400074f3c000300d040f3fc1f300143d4f1cd0030000c0dc0c1033d4000d0101300700f0cc00003fd113000c03303f00000dc0d415dc0440000f00010c41c0c0d40000135503000000303313d033c0cc000000dfc000051c0000010000000001000c4f00073000c30010310cc5000001003005dc1c0d430c0cc031003d04301c004d07740c50d00334340047c7040010004443000133c033c001d0130300311005004301004300cd30070fc030f473c00c1030030003c4300033c5400400707cc0400170700130100c3000040c0f3110703301100030317c03c4430c0005010cc003000000303035711305c100cf311000c0d1c33d00c000f0c3053f11cf000f003fc00704034300c05f0443d001003f03100110f01c300333040330dd37cc701314f043000003040507000c70700f0c0074300c00047d33cd044cc107c01000c0f1030500f3330c0001c1400740c07437103c0034010307c0700434033030d030410010c000040cc300cd10000140110000000300040f04370100431401c074017f0cf00113d34031700f01041f73440000000c07300c4c0303c4053c7303c1001cc0cd3005c014705f1f303c3300c000371c03440530000013f0cc003010d0c0110374370f10007c03011c000c1017140cc1003c0300000d740dc00440d401c300000003334f5cc00000143fd300100110351c0fd04130df10030c0100170000300d30000f100030dc0d0c00004dc30003410c30001c00013c004100000c10c440005033030c00000000031101034000003007cd003044f0304cf04070d7d00300030000fc00c0000100400040003370d0030f3004030144d0047007000f430d334004c40013034c3004330100030003013400c037003c0d0400cc30307c100135d040c004fd0c010400100410c317f331005135000033300014c01d13030003cc004100f0c3000113c400504003d340330f01300c00010cc01c0000000431c00d01170003c1700100400fc0140005f0c070c003000101c40003014030d00c4f57400fd03300000c000030300110003c0301000040d0fd00f04100010010c0c0c74c10c1013140f4fc00354010d10000030010d3c0704070010c0043003;
rom_uints[578] = 8192'h34104000d0140c40c400f13000040d34003010f0130f05300000400033000000c3014c41c710c00c00000c707443004f0c307014c41300040341c04370005100c000c0c1cc10f0d0c00030c440c34430c0c01f10f0534cf0040034400000104f00c0f00110037500c030f0c040010c100c303310034000403001c0c050035300c5d0c0c00c3043cc00000c0010010c50c0000d0000c30003050000cd0dd0ccc000040c000c3c1cc0030000c0c000000c0cf10000010304004040004f3003330340c5c0300001c0014010c00340533d04c00400c1c4d1c014000c14043c5000c0c00000004450000000000570ccd307300003004004d0c43030f4000f440000c003351c34004014f0ff4010f0400300400cf0307113501c00c130000403c3c0c000400003d5c0541000d034d1f000d10000d0301004000000c70c0004d0100100d00000d34370001400700c700c04c000010033130010fc00f5f0130f03c00040000c0ccc0030040010c00400044d000043101c044030103443c0cc00ccf0c43301c50030c003c4154401c011c3c3c3c1f001cc00d0004104140000030010f334c4f030c0c100000004dc30003cc440007430d30c0443cccf43cc303c1000103cc030030304c1000005c03000c0c1cc0400f0c0f01401c4c00cf4037000401fc004cc1040c04013c04d0c1001cc70111f4003fcd01304c400ccf500400d031004cc00c131000300cc01074300c40c0f03001c035c0000d7c5100010000001c0100013f314454071700101003c30c1410000004004040300541c334104000443d740400133c01c04c003407000401000c0c430d01cc04014000300c0d0c037f70300000c0700c00c73103103010000010070ffc01d037034d03030d01c4554c3003001c0c303c005c1004050300035303751c0100043304330007070cf1410c30370400300d0c40000c400031014130000400443f003dc0043000030c1c7000003d00100000000003141c030001c0130000c30000c00d004cc330cf33c41004400c000100044d0f40030013c003130c000d040c40001c0c3000105d04dc001000340011004d00300d4000047c11c70000dd40f330dc00040010cfd00c40d40d0c5007003130cc013005000c0101340f04040100300c3143000c01f34c044c010fcfc30c0c033434110c3141004c0030411c507d3700c000444cfc0c00350c3f0d00070ccf033c003333040c030400c104f1040c01404101c3c007000c570c0040cc003c03030100c0330300050d4003c0071cc0c7000305330703170031c7043c30300f343c0cfcc30c310d000704301c04430300140031fc0d04000000033303300c3ccd0300110c404400fc70040f3c1c0003000d3533110003000c3030135010000c1c4300031f00700c404043037033000004010c03300140010f30000000;
rom_uints[579] = 8192'h4c100030377104d3d04000470030403000104040304c003000cc030415d0301c000c03fc414cc4403c140000f0cf3cfc01d07f05101fd5c00000c004c3c5c05cc040c04031400370c000f30cfc040503c5c011001c040330d0f3f5c0033130410050c340734c1710031cc0c31cff3c000400cc00003000300d04310ccc07000c000d000404c00510010400000000074cc43140000c00100300fcc004fc0fcc0000cd334400c0f0104500c0cd00ff5d410410d0000c004100d0131cc7d050000d3110410fc00cc040c00ccc10c10044730c1fc05007c400cc0310000c00140c303c3c0000040000033000453d13403c50440f050010000001c44c505300000c010040075c00f04441f0fc0004c043030cf5c0070cc00c00530c300150300c003000304000000040000304c000501004df17300cc000140004c504001f1c0c44f045000404c004000013c0007004f0cc1cc305000010c0c1f400fd0f3304cf000c00dc4000c00000c3c00733700001c000ccc1d040cd003000330c3000000040001c0303101510014371000c07c300f10d0000c00000c7700040c010c0c0400000400c04000005040c0c00c033433cc00401f404f3c0713040013003c105fcc0400c0c0104f34300000c7c00074030030140000500d404030001000c4040c001400c043c4001c4ddc0d4c7133000d0000000c5c443003c114004f0040413d3c70cc03017300001c4104033041c1c30c4c00f003cc30104c3440000000fc4305001053d00c0031404300c033003310d04050304400304410c01330c44007000070001c030030c0f3f00c7004000c4c7000c00c0000c300030053443407c0c0000400cdf3344c00004c0100340cc00c533c30c130cc347030000000c0400c040010003f1334300000710f1f7c4c70000f0c03400375001d04c004310d0c00c4c001c003414134c00cf00000c040d073c001030c4c41004f0d3c13355004340107700400434000004400310011003c0c0070c0001c0fc107000041011d0d00c0414cc1000000533440c0010000c00000000000407153040c010034030010f340c0c0303000041400000f1f0d0011004c0000030000000001c000c0000c000fc004fd701300004c003d003000000300000540030c0cc301c0d000cd170c00c700c141003003303c034000f014040d0000c000c000334f70c4030403044d00c4404d00333100f04cc00003cc50c0000000f504c000c0745d034d07c3340cf005f11000d401cd0dc0003001dc10c0000004f73f0c1c000d1cf74f00440c40501c0c0c003000710071000c01c004c0c00c43000000704010040c0c3400000f0005000c0000530030030c07cf0043d04431c00003c0000cd0040300003fc144cc010c040c4c004040100c30c10147300c00400d00dcc004013dc05000301070f0010c0000;
rom_uints[580] = 8192'hc003000053031c0370000fc5c01074d004000d04c115004f33514c34377340000000fc0700531c033c04001733441dc30530001000305cc307440003410f13f0f30445cf0014151000070c5f0001c03dc0001c0cd303c40037471f00330040c40f305400100333010d47000001110d00330cc73c3dd0c0303c0307d01c3c7f3000044400150000330fc30410300100401f00070000f50c1c3c43004c051cf553c40033d340300c04113c1d3c57c0fc10f4004100014107000070070551700c0407141000c303130340f11041001f3003370c4f303004f000c410000c013000340010000004000030035003330000303043c300c0043000c4c30030c000000f0303041c0cd43f3d0f4cc0c00030001303453431051c00003c04000104533f0c00000c30070c04000400100043310cc1c0330343301f030030030000400c330c0c1c30c31100fd5105733d40130007057044f404004731031030170d503f04070c0f30435403c4f4f000cf10c10c101050401440f030301000343fcdd135030405111513373c4030030c03301010130050400030cc00000010c3cf03000c10745041d331313d050c00000401c000030730040515030131007713f303301300333c5fc4300033030f430c13ff04000d40143304c50030100f034c330cf7c3cf5c131f0d0f003c110700f0c43c4c0c0011037007c314301c333c0f00004fc3101f0000c017c3000f4c033147c3047103000034c010300f0c1c3304000303dc0114d000034050c4c1110003c5073300000303c40d30000713c1c3041f03cc003733d00431dcc010040403330047034445d001301310001f03333300d00d05400305550400300f4c307c0f0c10c350c04133071104d7cd030010000c05000037074fc003044313c0000d05c47fcc100310140301f1df0301c4040c000470c30f0300f134c001fcc15100000030137010000030dd100000340cc0073c344c310c300f0010cd000cc00c1403000f330c05d143c0cc04041043c4030700c10f730dc000455001c003031033000000403031014000f000030401c0033f000c13015400f0301f1c00050000170300014c40c00407dd01000310cc3143340477300f0510d44003330c0407105f0140c40410c0150010f74470174c303dc0711000d307300100000f10c3cc071014000330045304010c000fd3040100041c0f0040001c003000131347731c10000c403c5003f0003103053403000543130c0c400c00400c0f333007110c3103f005000c0d00003333000110cd1fc7f0d00c07130010173f43f41300044f1300cd00713c04f007c0033300c00037d00003000004300400dc4003c300003004fc3053040103300133033000c70110313301304040310044c1040ccd403cc403040f0000c003034ff07003c04c000450340000000f00103301330;
rom_uints[581] = 8192'hc40300113500cc03401003000cdcc1cc7d0044c000c444405c45c30cf1f00400d037c5d340037cc0cf3030400001001050003070501f0c3000000004c30000000c0c0740d40011c00033dc33003c4300f000c3331c00073c4f0cc105105041c0414d003044033300030c0340c1040c5330001dd70003c044003404401dcc403340013410440400c4c044000000070504df000000340c5dc00030c0040010403f000f0001044000443c0000043000300c034ccf000070c007304003f00740430c4141414000510f103c0007cff17cc0c00c40c10040c34c01100440001c00c3004100444f4c0c40400c0034f3d50fc000303cc00300000004c00033c4000c13c00c00000033f0503cc001030fcc0c00414c4f00103030000100401004017c0303040c00cc33003500000310440013cc00004440403450d0300c0341130170c0f10c004dc000d0c040001ccc03c01dc0030f030c0340454d0304040f700c1d40003004d07d330f00400000cf00003430410c4000407404000c05730103331000c30007c3c0d1d0000c0d0404004070dd7704040700000004014c40014d0710050304c04cc301d0d0c0c37000c0044c3cc401c1410c04101101fc300030303fc00fc40000c037004c00050c000f001f00c0c000000cc33c0f01f01c004c35000d00040ccf0370105100c0300405c34c0c44f0400c0503ccc303c000f001440d13110c040c0000010c00f50f001c054ccd03004000f30c04cff40c0c0d43c0103c0fc04f313d0500c30100c004dcf0c00001541000001ccc03c07101701000117070010d00f0c0c4104c55500c11c000500400c00400c00000cd10400ddd03400c0f340003c30ccc0000d0c03040400334c401cc0cc40c44043cd40c00050f00000c0040d00c40030403110004031500c0f0c0d4030004001f004000000c03300c4f4f030404c3c3f4040d410c4d3cc1c07010000000cf4f000c04401004f10000d500f1303100c0003403400c0c301c000007501040c0400dc03f054c0140040f0100030c30cf0c03c0100007c040450c0f34441c0c04000cc7c4141031d073001c4751c0cf10010c0f31c70d0000031034c101010c0c10d04f00c041430040000305003c4000400c03000001ccc0c401c05d0005030c04007c550ccc304c07c334f4cf11c3c044450c35c04d10c00c10370300013045004013c00010c400ccd0f47000c33004004c4004043cf40041d03d000c411410cfcccf04c0040034033c0000303040000f3070f10f710143c4034540000334c03d0000c034304c0cc00f340c00c10cd00dc337c3003010000345000c000c030030031c00cc0000010307c0f10fc4003007404c00c005c3cf000c0c41c0000301c0d00040004000404001340043103c040cd340c310000007cf00000c0004000cc34cc041030000000400;
rom_uints[582] = 8192'h4c00013434c31000300000100000d13c400000100cc30000c04c0c0d0000430c0000514010040000110000000000c34d510303010111103100400c001130030c0014100003000300001011cf00dc401f0c03c0033001017301110f003030001010000053000500004f100043137cc13000100300470300003000000033c1003d0307000041000c100000030044101400310010004030c3cc000403033110010d000000000510c34dd00003f1000033004c0c00000000301533403c1c30403001300010013000c00171c0334c33103c003050c003330d030000fc40c3d1401c00000dc0c00000101100003310c3553003c0113f403c0400400130105033003733c4330c0030dc0010001000030014701c7c330d110140004c1100030c030c0040513c0000004040003030f34c003c000005001d3dd50100010030000c40000003d0140ccc40c30000010c51f0c00d400010003013000341030405c4100c00010034c00100103d0c00000000100300d40001d407000130007103d040011010c3dc0d4341333030733c300300000000044004040100000000cc0000000031001130c31d00001300000000000103c00001033c30c3003f3000000000f4000041400003cc1cc000100fc03330100c0000003f0c170100303d00001d1001000df0500040d0cf0043003c05cd034073000000110c3cfd0000c0010000110303001007030d33030001103d11330c000c0c00d10003413101dcf7103031013c3c33304cf0d010d17d00007300103d0331000700000f330033500ccc0c0030013c005110c0003d0c4130100010300000771510034000010000030000013050c00d31107030fdd0043014000c07010014000000f00000100000d0f0300d03d1004311100010cf0337000c00004345030040400300007f0001cc00330c30407330000004d0fc0f1000500341400040110011331d410c413f010011531141404003404100103303100c0c0030c1000300f0103c001500104131143cc13013000c1110d0c000000000300300f000000301040c310001300000f003331140330001000c1c000c1033030c10401131c0004741000100003300000100000335301c00303000110003c00000030c73007c303030031500110004300c0013000014030000cd0d11315100fc3c100f000103000000500c4730004c03f003007000001d3000003c00303d33014c100c0015140c003000000f001000c0001033c0031d00000c730c3c00330014c040300c401730000c1c40010041330100100100400c00d541cd1100c00013000dcd403104000003110000005400cd3000030004c00074010000c0045cc3ccc14400405c13300041030f00000010000401004f14703007001040d74000053343033d4000cd0000000030cc0100010030400001dcc10f340530110050c0;
rom_uints[583] = 8192'hc10f0310c4c400c0701300000300f303c30310000c00d033000031f03c003000c003f40400f0001ccf4f034301014070070040000c00001d53010000040001c3c400410c005000004000c0043d000331000440c3000c000f4130303004000007300300d303010043d0c0c300044507d5430c4f00404d4c0000400705d0f440007c001c300343005300310011c10000311010000000004470d33003370310c00ddc0f0c00314c43004c000300f0c00040030140c00004504403034070c00040110403c00100000050c00010d3f0000130c031c03000c130000c000000f071c003f0c004c03400c000000001f300504130101000c0d01100010030000700000004f0cc0014400000c03130f444303c330031c000f3101fc343f4303430c0453c00003030000300c0c410d0c0000d0404c10c0f003140034100c0030dc110c10300d0f500f00cc01c00c1710c3010000040c0330000dc000053300cc0c0c700374000000030c003300f4000001103c1c0c3504000f7403cd443c3f303c3c44c00f1cf0400031c00405cc33000007cc0c0dd7100c0011311c500c5c0000c0001107044037c1040f0300030704010c400400011c11015c34400c00cf54d0100000034c07004004c40031100c0030c33000340730000c00310030f0034c30300301170c333d1033dd00440d303350017434000710000c334000030000c40c0000011c3010030c400d300cc0fcf000043c3c5000000145003310c134f03cc1700c3c3100113410c40d330c001000301430cd000f1d0c10030c01051dc0004400540f0c03c0153c00003c0c400310d0100cf4c000c03dc3000cc0c14f0d500c0400017c0f0d3c0043c3007c0130030cc300100c70f140300534004c0c000005c0d4f0d1000d001107dc141074cc303300000c40300310c1030c0d000040000001c0f30007f43cc0403001300d0c0010cd0001c300414d0001003cc4cc0400000001f044c100000030000c3013303c00c30c70430000103c1400001100000007d0cdd00004100c100000f001c00d033310000c00000010000fc40000c00c400f0400401300310d4300f10410c7000433103c003011700003031001000c04000c4c0003000c0310c40c010110040f54dc41c0043301c4d0c304030000c01c04733133344c0000c03400c00d050000000f000c0c340f01010c503c170c000f0000340f0100310c3c0370c100040013000110f0001c01c0300040110c33300400005d004c00540c43c0cc00000cc5110c04153f0c370f4d10000cd500100c1c0000f1df00001d3c300130003440730411110113d007001cc00f5c17000401d130000c0c1473330c3700f0340f300014070f7030040000001400103710c000300c1013000c043c3044000004013cc1003404000c003003300003cc0440c0334c00301ccc0c000;
rom_uints[584] = 8192'h1130d400310f4500cd7003031300c0437f13c0c0010cc01400153043000f0c01407307344515001001014000131031707f4c000c140100c50c30010c0000f0c4d40101051000000100000045dc000000c100313c0c1c037cc000300f00fc400000dcd0dc44300c040404c100371c03000c0400c0c110075cc0300031c1400d0f031400103d7c007050700070033cc4df00300040000053d033530f71c301751433f034f11003fd10074000151013c3040707c5c100100c00c000c031400f000007c7000d0ccc0143c0cf00c4c0c00007033017fcd7310304c0710031d303100cd0400053d00c00010330000703370c0f401c007334100104700000470000004c134111004d1003c5503c1040cf30310c400301f001c70313f000c0c340c3430000503c000cc4000340ccd0c41040f3343c01d340701040700470431005070341740000c3cc0054c040d03f30f40440ffc33350400001d04000d33c0300730001d3130fc07107300301000c40d000443400001d01c00cf300003f0030d01c15d0310100733c7004f3c00000000404c0001300140101001f5040c0040003001c4d40757cc401c330004043c03c00d1fc03c04c1001040040070330430000f0c0100003430df30010f40dffc0401fc00504c4c0c0430f40004040007000c37000410c33003dcc000c1c050ddfccc35007d004700357301c407c40031400500000ccc03ccc3d00c0c0107c40c03cd040400c004001c03303d07734015c3cd000050f40f0110004750000000f1310340c4dc00c01c00000470030c300f310c0003330c01d0cfc00000040001f341000d0011100f00cc1cc03050074cdf3cf3010c1c7f10340301d3c3cc0fc30005c111000d043010001470d35f340cf01041001170000cfc00dc50c00130d51c4f01010404c003735000073f0c300000f00d040c341c3cc1004fc313d01d504444014043f073340034f00d014c5c0c01301d43373003040d004c7000470d0140000c00103001c004050510c10cf007f735d413f00404000c3431401d110003400300cd01003c305c14407c00c00030470c05f44d34001ccc000117c000c0c1410401400c001f3c3131c4040d00330001cc0c00dc1c1c34f00000cc57f0000c001c0cd4c303030d10f0c703010054fd1c1710c1031f433c0304c00f00045033cc01c0c30073007403400c0034c4000cc00c04403130130100000103c0010d033c143ccc00f033400c03f0d3d01033c00004c073337000c41551333007d5ccd030ccc30304c410014f0c7507c4c000400c3430c5f000f031c10337334300000dc1033111003140045cc7310003c7cc0cc3c0031f5cf30003cc07d307d73d103c0507f3170cf03101031443030c14d411013cc00dcc30cc730450375000000c311c03004003300f3701400015f00003d030ccc00040300;
rom_uints[585] = 8192'hccf0014c3cf03044d30c00d1300134017c3051f11c0100f0000000c14d541030010c0ccc0f100010007400d5003fc0433c440040303007d1003040030037c30403004003005f0034000030033034c43cf5cf4344c3f33513f0c1f7dc0033030c107c00300003033f733cf1040f03c350c4340013d75c30d0004fcfc041100335cf0c000df053005101000c400001553c7000711003074c0d70f0310303500c3011cc40f103371003d310100d3c0037f0fd1f500001004cc7c070100f0005000c00530cfdf00331f0f13c0f30003003c00f1c30c00f04c3530340001005c74310313004c0d7700400c13f15f00457c030047401df330000403173040040000100f130331000f07770340301130103cc051d3015cf4f3ff00ccfdccf00f0f304133f10f003433441013340c1135f5703003440c5c0d405d000351300330300031c770030344f0100130430f035d171f70c34f0011d4df10c000c0dc0700707f0500c40310c1dc047c01040c1003c0d0000030c700300f50c33cd010130440c40004c05313c41145c400400c0001f000c51030f01000004030c007003ccc440700143300c00f37000c040340340f00dc330c01c5011070fc03c00d01c31317340c314c0143330c11303ccccf0c100c150033c0000703c143cfc01c00100cd414100100503000c13c7134c0030f010340005d5007d4000d3c5310000000c0c3104c074d10fc00ff010000704c31f0130c037407cd01130dc3c3100734040513350471740144033113c03030df0ccc0134300cfd010001ff3d353003ff004c00c003fd01300c003c00040f1f07c00c03c00c0300070c000c53003d3c00c30000c0fc030303004d1f0030f00c0c074300010d370000c004303033000c150000c0d000c04d0c00410f0c31f130f5330c73d3030f413034030dd30d100fc3c3304cc004300113010f05d1f434c0c37f0007131f00f10003001440033104c3c0030f5101f0004c3c000000000057d0f0000504f310c0f3d1c33140f1dc440444f0044000c7000c30500000300c0c030c00dc010f0f3003c4c03c043400100c0cc100ff3c0344cc1033df33f54d04031c004410f3f1400301d0171101c34c000ffcd5f3c457033000cfc0f40f0ccd03400010400c010cc53303d01d0007f3300300cf000c13300c000301ff30033003fccfcd00011d00035dc00000331c3cc7073050000f1104d01100c00070f74d10003c00f00304f007004c3d00101c30000037033cf331f0c7000c000d14d000104030ccc70c00cf00341053340353007300c5300131ff0d714c00034307cd010071cd4c003f015070103d0005370000000000140033005130c41030dfc0010c171304100c0cd3000003300d00311c305c04013430df0004403100131003035c334d013cf337731301300035405ff1003000030d1301;
rom_uints[586] = 8192'hc000400303d00304c0c0c105347004033f030d330000110000c070c000d5000cc0f03300373404f0c5c3100100c00410f04003300f341cc3f010400c0c301000ccc0400c0cc053f0000004c17004103c331000447d100d0c3037340ccfccf01000001c1d33003d0001433000070d100c1c0dc01c1105c1501c7cc00c0700100500c33c0c304000000504334010030051500c04100141c00440d1300040000041441410011000407003000c504f0c0000c0d173c0000c040f430301ccc0303c3400300473c044700f30000c0d0c104010007300cc0d4cc0fcc03003300110040f53404d700d000130c3000354130500015c40304ff40000030030c0cc03d0000c130010c0304c0c400c1c31300410003450f130f00000c00f400345570004033f3c033000003d14100110003700c003c4c0c3c0007c000003f400c00f0c000004c41f33f054c4310c000001033c14315001f0550003d0047c30cf43103d0c07d00c0050c4f4c40c00c00030307f040330140303cc0c1fc4103f03304001000000c44c3ffc0431044cc0100010000cc44440000400300c000fc300ccd054cc30400d70343d3000000000107030c3c400f004440353c4c0001100104cf00340c700014411cfd0000103cd0f30403000d3c150703c0030050101017034300cc310f0c30f010300131d0c01c05130d004010cc04404fc30d035004c10300003c0003f043c4370040010100d40c300cc140700d007000c3100ddc4c330743c003344714f34c34cccd03d3010cf0004340010c313cf113031f4dc0c0f3f0000100030f3045040c03c0500430f0dcc0c0000430d00c34004000000c7010c1010413cc04c040000c14f000cdcc435cc00100000c14004cfcc041d40300000030053307300045340f1c3000c1c1c40c101c0043c0c04cc500730001070034d4000c53cc30cf0050133c74c0c103cccccc003f70c3031000000000d1400f100f3710400ccf0003140100004dc010030030004300c0c0c333000400c10c40017444413cc01c070000403c0fc300004d074000031010dc00c7d143010300103cd04040d0c0003fc4c50110cf00000c0104701000431f1000300c010000c1430044c0344143130c00000c05734c4100f4103c0000d40004044cf0df53400045f103344007f70003c04f01c100000703c5c330430000100f0310c1c0013cf0133703000003c300003340c0003000000001404444030311330c034f0005330355c0cc3304c4034350c014000000ccd00731003544430c00cdcdf31304cd300303033d004c0000101000010104000cc40c0100103c000013000305400d003fcc01004000037004c4c0355fff33cfd0004030133f0171030cc00304000010030304005047003100cd0304d31c4c0c330f003403700040c3c3004003ccc00103051030f1040400010c;
rom_uints[587] = 8192'hf0000000c0fc040070003cc4000700c303043f04dc0470400440400003d40000070cc0047c310400c10400c000451cc0f0000cc0010373500d00041000000000f114000c0000103c000fc1000c043c03ccc00310d44004040000100f0f0070f304c07d014000c4440337c0007c00c010103444311d704004000c00c01c4404050c01300ffcc040530031000cc000473c003004000d0c00000000030c0100417c001c40000430f0c0400000004cd03f30f00c00c0000003001000401310f01cc030404000c0007000000c0373cc0000000034030d0c07033c7010ccd0330104000c000010074100147fc100d000c50000cc3440000c000000000003170000004cf0444000070000f00cc0000c14c103cc03400400413ccc0f000c0045c0cc001000c300030c30340f00000040f0c0d00400d070000317c000c03300054c43010011cc1d77c00000040043c000747333104304d0c0400c4d0404cd0030c0c0c0003cc0407ccf30f40f000c311cf03f001c000c1000cc00005000c0000004000333c000404030001500101040430041f003100040000043c1c0c440000cd000014c134c0004d0430400045000c3c0cdd0100c01050cc00c0370000400ccd30400c0c00004c030040477cc10d007c0c0310f00f5c3430f0d741030fc4000c40007dd00c300d33c0cc01c0410340000740000040400d3040070c044c34cf33000341071c0c70f45cc0ff0000c30c40f030400037c0000300030040003c30f04000000000140000d34030000cc100c0c0004000d0c30000000413c000cc0c0c00cc0c31d500cc0c0c0000133c4000000140c000030000f00c3df03c1000c0f30041f34ffc00005340030000c030c00c0000f045c30c01074cf00000040c0c1000300003c0030c043c000c44f4c3ccc703c14cdd0cf1000c0c034000040cc000cc0c0c1c74d004000011cd0f41035fcc1300c01c004000004103000d440414c43700400003c477c0004010d00300000000000040040c00d33f40dc574030444140404103003310c10d4344043c050304ccc0cc00c0000d4047334000000040740030000710d410410444cc0000040004031000010000000030541000404300c1000f00410c00403c0d030040100f3c115000001000ccfc000dcccf00000000001c0c3c30c00cf00000010000cf00c3540cc000ccc01030435030f307fc4400c04c400050c0000c410c003c100c00c0c0c003003fcc0c3c037341011f300003000000001c0c4014030c7f0010300c0c300000070d0300c300010c00040010001c3c0400cf4c40700f1f0034c000040c00444014003330c04000f0730c143c0040040530004f4f0c0ccf14000000d03c000c3c0c00f010c00003400030045c03310f701101c04000c4000477c30003cc44c00300f30000000040510c4100c0070c1c1000;
rom_uints[588] = 8192'h114300010010010003c10300c3303c1cd1c0103c300450130310cc0013373d010430031d00fd00103040f0010003407344071f0d5401c0c300413130c00104100300013010110c0d0c00d00c0104fcc0f00701311f04034f14005c07030ccd13030031c01033030011000c0340131f430003031000f3010010140f0034c3700f13c10100010c00c00003000040000403100110f000033cd30d130f0041041d0000340c00f3c0003f3030310040000740c4335d0000003100000100730144030001c010c00003000003100000000103100000c0100010133c000f30031744030cc0cc00533001000000400343014004d31300300400010030c0000330030100dc4300400330f000040030330c44337fc003f50f34f04c0000d30001003077c11400000000404c50f30033110014000157d3000344433cc000300034304115130f031c01d030410c00751300f070110f000013113031c313c43030f1c40003c3c104040c00dccf07003414cc1300030d4400303500033400cc0030f01340033d013d50c03000000001030300031f00d0c1030040430500d31c0c303c040010000c0c1c4000500000dc0c05f070003d7400543401305310d000003013000cfd01070010130034000133315033001003f03c11304f00d0d03310000c0000000003c0f33300fc000c30c401000047131330500000370d301705310c011100003003140043500007003310005130300410fc411100000103000030130011c4001c1001003033000050d00c004000034c000cc1c0301c004300300100530d0c03000304003000c073100f1100fc105053010d00440c01300c30030c033001500c013d401003010c10314300070f5300003040103304f0301c03100000010d0000d0d30c3371303c0000001001f130035d0c0f0000443c00003000c30cf450d0043ccc0d71314000c00001300400c0c130c1003cc33305f0001104040311070d400403013c0c043004000000405000414404000c030101c000000d0c141107030331070fd100000344f0d0c0100c4414d000300f45011c3c10000104000051cc0d0f3011c1300350110ff0cd310001cc500310110dc03704dc00000000301017f0343f300cd300303f00c4034c0003c0010100300030c37001cc330df4f0070000400c00001c4c000c0c040100400000330004004703d00c01431031f37000003100070d30c000701cc31035cc300001300035503d000dc7c30144030010000041541100c43d0c140050c303f1330131c130ccc300010d0000f371000340133005070313cd00100c0141040d0000013cc0000013007000031c0000305000030000700f1c103340000cc5503cff30000f0c3000001030f003003403141c011003000010170c00001dc03c051030055d001c0c4300401f0031050000c03404f31c04013000;
rom_uints[589] = 8192'hc14003c0030041000001f000c303330ccd7f0030730003010013c13000c00010c0f1d14100f300700000000340003c34c1cf003c30050000d003c3001c00010100404d4300010000c00000fcd1c0d0d033dc33037cc00303100070d00030c14c4c00730101000c11f3003c3050d531700000d3403000c1c000d070040004c0011374f140013010cc0000000000040033030443000010c0f3103033130171f0404440010303401030401f30c3f430103300404030000001000c4100c051c35c0141014000700fc33300344000105043010d1013c0010003003540000100c05030c000000300d1c04030400000030c10c11c0300000034400010c310c301000043c30040c000300d00000303f0031100000c4000c05140033037c3103f00c330001003cc0071710003ccc740fcc101010010f003c0c003400003d5c0f33011d0000101477cc0410000010033013400103001c4c304730f3113c000d030003c30030001330c0c1170d04c00004403054c430000035110c10400c00fd00fdc5c710070304300ddc070c010430000440000cd7000c40fc000113104c31311730000007453c0c37300010011400f33d0413343c0d73070f3d011034c01130040000134f3c01001cc0c0001004073003f30d0004500fcd31001c37c00300043174c334d033033d1c71133430dc310c000dc00f3331153000c33c14cf0030001d100000030c00300040100c010d00cf000c00c1100d43340c00dc0070030c0d030c00c0000033000110000d100c040d04000001000300030cc300170304000003000c1000043d0004c1000000333d100000d4007d01040003000030000d5f0300000705350107030cc30d0dc1030c4c00c3000711110304301c1004030c03000034000100c3000cd113000f30003d130314d30c0000d0001001004300131d001d00c3c305c0133c00003400035305300430101330c0300f03370100030d14c10014301031d000400c00000c0004340010000c31001c0c170c7c040000c1c00c01130d0130f00300c0cc30010004300f30000000000040340c000d3003300f000c1cc50c111000470713c3cf40040404040010003010010035000dc00403000f30001304000c0004f0f03d373d13000337c1440c0010371c0005d030043c30300c03033433c43f303303143035c3000c130010003000340f013040340c0f30100313c333c5003307040330040333003f31c00d03040c140c003c04300100300c01013500000c131c30d0000035413c0311033c440303111150033cd4300c003c0000000d1433330100300c000000001d0031001d1001000f000001fc0030000007071f30000c0011c7050c3f000f045001000000001130000700141c031f30030c00403d303d0c0005100d3d01033014330001001400033d101f04cc001000033c3000000;
rom_uints[590] = 8192'h30010001c5c00004130f00040005c0340004040d5d0737000d00000000c7700010030c03030c10c0d3004000000cc4100c340d00010001001330000f400c000cc1c013030004040f000070dc70000c400130034741414ccc010f0d743dcc4d0007cd005034000fc0014730cd7140c0ccc0cfc4340d4040000344c50d000c030c400000300f4003c30750010d0000dd4f0301000000404dcf3300d00fc0cfdf0d30c0c403734c070f0c0cdd404504000c0000030003437f0043410f0f7d403000d4c3401500011430000c35c0410c0c30030c04000c000c0c4300fc00ccf0c51c01000cc50000010300000fcc0030430c03f34000f3cc000000000f0443010c13000305c14374000000f037c33000c0000f0cdccc0d40c4400d0007470404104d0034000f04530404003005c40311cc0f0cc04c30030000030000c0053c03ff004c0100000000000000c00c400003cc4f0f0000410c0c0f40c51c4c700001c00c434c30130040cc0c0d0cd1c1010c44c30110d4405347034300c04001000034010347074c00c100400000040ccc0cc307400334410c014ccf00cc0c41f1000000335c0c00c040c310c30140c4074cc0044f1d0d0cc0304f0c0400c0cc0c0143c0c71003040304000000c4c00000cd0017300003444c0d0c10f7f00017c3cc0711100c7c1c04400d0d0300d00fc30030c400003c03c0c0050c40400040304d710c00c0530f417c400307cc3305cf400304cf4ddf0070001d3c0fc0c7dd000d010004ccc00043000141c0c0410300011305c03404000c0005cc0c3704cd04030dcc3c4fd0001c0300c005000503135543403c000000c104040c01c00cccc0c5c001cf0400c00f04c310000ccf0f000000c374030d010c0443c0f44f000c47c00c1003c044d0100f03310f404c4c401c1f0c0c0c0f000c440d40c040c3010d30004c0f400505005fc00ccd0c0d000000d004010c0c041c4d330c0014c7004c00cc0c0c04c3f0000dc0307400003100cc40c04d0c0d0041fc0003c0030c4f3041dc04400040c4c4cccc3303f0040401c041000d4f030c1f0c000c44c00043004040050d0500cc4fd33c000300710f000431cf01004c4c00104330c0c301c14014fd0dcd400d0f410004c1000c70dc1f0454000050d303c710410d0000c300c00003c77300cccccdc1cc03f044500c4f0c00000100030f0030140f050f040031cc0300011000d10443070d4000000f400c00310747043000c1c3cd00340d004f40cc00cd10cc733d00c0004f03c50c304540530c00300f000d0004000000cd3033710f3000003c00010c400101000f004007400f340cd000000f010001000c000330440cc0040cc044411040c405c0434404000040003400704d030045cc0440003300034300c0700073033003c000c430c300d0c1cd4c4f1f5c040f0c0f104c00000;
rom_uints[591] = 8192'hf440f00c705cc40dc4000301f100cc00c3100010c034c4c130f30c50007c1c4000035c43d4c7000dc05000000004c4400c01f0c301c3fcdd4c1310f33001000c0f005704040014c40400dc405400300414034050dff3003044c113300010c330c33d0010010344010c11130c34d45cc3003f000f0400007f00043010c030033030150fd0104100fd003dc0004310c04f4501000100000031505c04c3011c400401000d104030130000070040475c00f40f30c0d40000c31f100304040004000c5034110d4c00ccc40f30c4000014fd51f0c344130c0c0ff004000440c00740100300031d30c00c0000c40d5c11f773344c1ff00c40c0c00034000005310000001300cc00c4007d4005c30c34ccc0540ff01c00c3100013c000300ff410701fc000f000000500001c0f3100c030040fc03000430c34050f001cf3c430c0341f041143143cf0033403c301304c03fcfdcc401d0004030dc0010014013c03ff3303000040005f353f3c505103c0c00417c3400014300041300d53433040000c0f010403f07554300000c330000c4451f0c73c004100c000000d00040f40433100730fc431001100041d00c0c0c5c000130c14400d474cf4d4030d433d000cf3400000035031030414c30054030cc1000000c4c010cd30403fd1003504331c4131035c00c130f043c0c011001d3c00f53f3c03f000c14ccdc001710505007104f00057c5003cc40004010001f340dc1c010004044137343ff71dc30403fc44ccc53c3014c030c01f4000140cc4000040443c0c0cd0000fc55cc4c0d40000cc0700500c000d41c00c1100300f7f3000503dc10004c0c7440d1c00f40040000000530001c000c4031400005d041110c1000001c100c310000407c300c001f04c04c1000003cf14040010440434f0100400301043c043350345300000405c010c0f0007c0004c0040135001c00034ff045c140c4d400400400df0011c30cc3430c10f00c0017103000000004004cc04000c3004ffd00701333c045c0073014043d500000000c03c00d0c0400010d003031100013f0040411c100400004cc50c0c01004cc13500d3017ccc40d7c1d04f3d05c0c15140004c3004c0000c30c100043c10d40c00000050300340000fc44c11101001034f4c5f044103313c5001c0317c00c1c301100101f340001010400c104c1c010031100010030703cccc040407f01100f3001ddc104000313004303c41303cc014030c007143f31ccc440000f4073f700fd005003300cf0004000f131370430040014c304c0451403130d5411001033c03f30c570310003c000330300cfd110c00c0ff0cc4004d01c03fdc0030f03d0c0047304f01107d10f103404c073500003045cc3003144001000003f401c4004c40034401c310c30403070407300100040441000510310000044351c011405000;
rom_uints[592] = 8192'h300000004c010031104000307030010000150c34c0400d5030044d40c000400340017c110100104000040000c003003043100c00340004c44d700001433130400000100c001c340c0c0003c47c10c440c50fcc7700c1004003001c3030f00000f003f0f04d4010400300dc000031dc30000130c00010404035033000045403304305cc0003104100400c0030c31400000035000c004c14000053104c43f01300c0101004413cc4d00033c43400d4003000350cc00000c7304010000fc3c0000030110c1000000003400030000000c100040f5c40004300000145304000c501c0100c000c30041c0030c70004f31f000c0040053000070cc0000000007100c0cf3c13000000335cc3c0f430d00300403004050404d0c4c000050c0014300c310070c3000014310c04004011043000f5ffc000105133040100040070000f0f404055f40c4cc4011c00f700f0003000011131344c00f1000d4001d110cc4031c10030d003c14740301303055003107400c00031010c000000403010005d03443500f0f0500d4403003000c04c00c030c11f14304c00f0004440f010ccf030011c0130430000d00100004100c0c340c0cd10000000f70c00015c300000c0cc1001f4d0c100f10c3000c1c13dd0ccc0f070c040300300770c30000cfd0300c0000f3110003d040030f00404050040007530ccd43455f10c1003cc00c000004d3cc05000c0500d100010f4504004c00c031307c3033104dc01007030104130f000d37001c0c40070005340c40000300c004d00f03c030100000000340350c1c4001c11070400000400000cc0c001500010c04300340cc300010000333530f00c00dc44004c00c050000074000c0c00301000c000c001c04c0700300040c0c051df000c00f7cc30300000c7005c0cc040043c10003c500131400301000d41000300c40405f40c30101010c10704430734f1000d41040f04030000350130015051c04100000030430400100050d00010000c10730010f0f05c30000c003311000c000430400003303004c100401c05c034000400cff003033c401c354cc0070040030030400000035c0c0041cc0c40d04000c03c331101001c10313404c044040400010317030100f00c000000cd030c100c04047d03c410403d004d43c1040001f3cfc00000c14d0000c030313040000c00c00040c0000733330f0430d4c100000554000400ccf030c0004000c7c0400c004000c1001c3c0300f000c0000030000343303303004031c03400500000374c0c4c10f030313d1cf03000400044c003100c044cc0f00000000140000304404040005cc0330030400000f0003000000000110140c0305f01005fc100c0730000fd00c410010004c30104400003301410003cc00404004c3010001f00c33cc300430d0104033030001004c00100d5c0000c04c0;
rom_uints[593] = 8192'hff3000c30105000c31000330c4001110c430000f004d050100100000004f0c0400010fc703030034341c3030c00c043d010c10300cd03ffcc0030400cd000c000035331c0105040000000f070d00c401140c0d153dc0d4000cf0043c00700d00037c043000c700c1140c11300c4c4d4d01430303000c004f000d4d00c0403000400303c405400000040cc0003c040f41510700000000000d044c00100c00cf0fc0440c050003f1003c000000353104300c4cc0010000014c000700031c0cc13074430f030400fc30010f047c0345c3300003c70d0f0d030f340470d04c7001c7031133c100cc0c00017d430d0c00c30c3c0f0040333300000d0c0c00000100cf70c5413c00fcc403c53c00100c3400003cd000300c05304317000c4f0304f41c0c1cc1001003740d0c0100000300414c00070c0c000c0035c303fc0010100010310011003005c004c10030013000c1000cc004040434400c0d0c0311000c0000003073703f34033c00000010c30c41c10c0300050c0c0dc003cc033700000434340f0130000000000d5004415f00c007130000000100030dc1040d034104101401c110c5c130100000033000000100000400034004300000004000000007c00c044c000c303c110001410400c00043c0000c0400c04ff0c40000c030410f00c40c4001c0c0413c0c04047403100dfc40c70f00140f0100c50004003000c0031144004c0000cc0033040c0400300101014f04000400004500f4cdc4d3fc0c010030f533040f4c10040c0114dcc007540034333c030dc00cc3303c04014c0003301c10131000300030003c0c000013c3040c3315007534c40000340f4103071137040d0430cdd400004100c00f0c0c000d001c000c053c00000c1cc00f4000c40030030f343103000d0c4007430705cc000d7c0001c010010d00004100fc0df0110cc0030105131040070400d00103000f004c013400c000030c000c14000440c70030313ccf004d074004003500101f0500c0c504000dc10330000c0c100101c010000c030d05000000040d73000f47033500cc50c00004033d040103030f0c00100c5d03150104c40400040c000d14004030000003015f000001c40dcc040000030f000730d00100c03c00000414300000003f700cc303040c4100410000140c0c040cf704c30400014000011c0f0f0003c1003c00410004300300003107073505300f0c00c400d44f4c140103000004040300070c300435000304300c5000000300c01f043000c31540433d0703040ccd33030304300d00c3000c00000c0f31330c70000c3c05100c40300f3c00001100cd00033004000070400000110c1c03003f3ff405010704000003340700000f00030300330f00c0000071c300040c0013001c40043000ff0000010f00100c000700410c000fc00c0074030c00001000;
rom_uints[594] = 8192'hc3c00cfc3300000100001f100400001c0c301d0000c00000304f00370403040333745cc33104003dd00040003300dc734105f0d1410fd0fc0330001f013f03c30d140744c1030003000f00000030c00001d0f11040040d01c3141000f0314000d704c107300011c34fc700301005d1000070c03c30045000c0010003500004c71404013c3d003d000303000041c0040500000c0000031cf004001c03041040000c0040431000030740c300c0003010033cc000003001d540c0000401c100dc0c30c0710005400134f000044111c0c4c0c10300c00cd4000c00c740f0c000cc01011300c714000c04100c10c00000c304f00c00000700c0410000cc01033030f3001003c440030c103c04330c10000400c000f30411030c5c340004c0000c003c140c00cc44000307001000303001000c007004404c1300130303304040c00710143000315c1c0014330040470040000130703133c35431fff0c034135340133100f030444cc000441000044000341504c144cc0c050f0c00c0f407c40150040c15074c000043ccc40c4700400330d40d005414c000704154cc0303413000411131d1030405000f0000700003f40300c7c00c1c003d13300c0010300c0c0703100410000cc00c040311c00cdf00c0401c0000f0000d30dd0030c04c0030010c3100fd3d0000c10c01003700040500c0100c0037071000c0000c0d300000030f0000ddcc00c00cf1001c03c0c33040000f00001d043000001f0173f114c0c00000f0cc100030000500030051400101004034000004010440300130411010c1cc145133070140010001010030c4d7410335c1100400400403000f0f003c0c1d033d1f404c14000101015c00030f00001cccf03c0074400403cc00100044103f300c0310010400041000400331c0005d0011c07033000033c400730500cccf0000300400070000c1c4c010401000331f003f35000003d134000c003c10040000003330d0070700000430030313c0300001c000404040c0011103c1000f00c04f000000cc000301c00010130c1c40fd000cf3000030df0430000000d1c04044000001000cd0010f404400400003007d340c0d330330371c0c0000d00c3000040c0c0c00000000cd003041000000c5c010100334013314c3c340100300443000000c0c0c40f000c001000000c0031f3070310434000fc11c0c033000f401130c00741040000004c000c0010403104030cf007d0400007000303700400044000000c0070c10030300fcc47dc0c3c0450001c03004033c774c00007440cf0ccc0004300c0400444000310100c10070001000470013031d00003ccc04400c00fd33c100040300314071370d03001000430c00d71000130dc00341700d430740cc0fc011400c00104300041340c10001304301f00c103430340d11040003000400000000;
rom_uints[595] = 8192'h301c070004000c353000d7c5301500101c40000501070000f000c030103ccc31045700001c0100450304dc400f410003f5530cc0340001300c00c011700c0dc000d7401f000000d0410031004370003d330c00cc0400313c033f470c300c0444000004dd0c00403100007dcc0c3003301cc001000f340c010044003033141df000340043c0310010444004f700100011000001fc0cf1010000003d1c33c51010000000500700d00f000004f40404d11c00c4100dc04000000c04301c31340400700004c00c31000707354f43103400000030300000303341030c00113154030c0010000000c00c04cf530d44fc1c145f400f000013040740000010c0f410c1470430001401cf0f4000000c4c04f500f004030cc0510f0c14f3c0701730004300f00d00030400dd03404004045c3000f0f0103000003430001c40f010030c5400f0c04c0004c0410c00fc50cc00fc1010140c00437014c40c0030331440c0000f4c4030000d71010c100031c300f10310343400003340700cc0003c0110c0135011340000703000c3000130c11400c0f1c000130053041000101704c404174071411c50c3310104d003543004007400d3fd4040fcdcc000113c30c04011f300000001540c10404f0cc400f3105010c135c4440050003700007c30033440c7c0c0000c473301f104fc4134f005ff30f04435c00070000c000c1c0030404713f04cc70f14c0013030000c003000d34050c00f00c00c3037c170f0700c35001453f100dc00c43000004011401135000c13c000440c1c101000071300033d300c0400000300311c003170c41d0d10c03000000cc31c1001130c00000413c4c4331040cc5c7000300031c400011c017c040c0300000f003013100cfd1504030cc40c03000f0341000010f1c000001c00410c030400003f030d3c01c030041337000c134000540c00141034143103f13153403000cccccc40c7040c01070d000fc03013000030cc0430c000131d033c00304041c54300131fc13770001300f040000f00044c033500733000130044303cc043f47d10000300f0c0307c0100005f13c304143c10403514403000000031cd3000340c44000134dc104f4030003c00ff00c00f410c0010003405100c03033300441f00300500005040100400004d030c41001c30f30040000c101c400d1000070007000f0103431f075004044005cc45c101170f0010c4000434704000fc5000070c10007fc13fc30400000710103030d50000003331100130f34404570c00dd0c0c00400f0010011c300c000040c30c0c434c305c05130040000000003d0043f4310c340330003d3300c00000001034c5745407f050003c31354004c0330000dc003033000300c73c3c00004000c033400047c0000400340c40404c4000f5000100f130003400401c00440c1300;
rom_uints[596] = 8192'h45000041c040011c0c30c0c340440c0041000cc0f431c0003403400c710c00003044f0f00500c0cf30d0300114f1030fd000f400445f14003334000001c0001730c04d003400003400cccc743050103100401043c401034c0403c7100000c0041f400d70000c0000107d0005c0371d3c0cc41c30d1444300c101c4c05c4c3304f100c000300031030334fd40004310c011303000cd4713100454c00730c0f534c03c301401033000c040010130034400003400000c1510114000f0f1f310700444c003100040000103000401cdc0030300000040c003040113003441c00030c104003c00540404c041001cf031400cc00c040f000401000c003004000000c0500107000111f00cf00054cd301f30401030005301007300d1340130f0100c1000c0c000341110110103504030c00040303440100c0553000f00cc1334000cc5c0413500c1c00100c414001c4471031031c004103c4d30fcc001fd3100c0700541400040fc00c100c40035f0400dc04fc0f00c1d1033500000fc5d0010030c040fcd7300c040d0f300440050c0c00c05540014000000dd000410c34004040410d0400403f0c1007f00f0134550c0f0735003f0d4f0000cc03000cf30cc01045cc04003cc3000c140c0c43000f30001c34000000417407cf0c0c0f4503cc103c001f3013000f015d1c50d1033300d40c0d1107000ccc0033000c104ccdd4331470070f00c04004103f0c31c3c40f0103f30000005030440030700330350034000043444c50000000000c0d400c0cc300003301001704400d30100c3cc1300fc103304c31000c0000001d00343704f00014001330000100010c00c0070fcf41070113000f31f015ccd13f03351303000000d10cc00134000430c04f400c1fcc73000503d015000100c30001cc41743013100000f0134cc7cc000000d004734c0050c40400c00c035044f3031c3054131c310057070100c01030303130c41340404cc0013434000000077044303400c00c000c1f3005407c0f01f001c303c041f33c400f33f47040101c00000d0000000004300303733040000070fc400d30305030d001000f1040430f405011d0000cc33f700c0300c10010030471c0040d0340530dcc400f0730040c71000003005d040010430403000041000510030c303010c50d0fdf0c100300041f1331073f03cc400043010c05c00000c00000d0407c3031004c00cf04000050513003033004300010f010300070f4cf00110c130c34c34d0c0f50000001013040013d3c44031f111000c0d31c107017000f403340300504cc0007c000343010040014403040000004350d0cc10f0010c0d300034403100071c0030c0140335f40d3cdc41d5034cc0103c3000000dc0d11400403301c33c1501d4104c404d034c44031300400d0440c000000030f0040c00043c00301c00;
rom_uints[597] = 8192'hc3cc0c00030500cf03000c00471000003f0f00045f41d30000c3001044005c0000c440104343010300cc0c014c001103c4130403104304300101043305330000040c1310143000c0000010ff4003030000000d115304100c33071c4500dcc70000c3c77cf0000f5f0c0c7704003011cd11001c054c74404d400c0154300d40004010f000000100300010c340c00013c1c730035c0000c3c45c0010ccd10004030f035c0f05c353c5104c040444100005007077c0003034010030c31c1cfc333c010c0014c000070c007000510301c415130307c0000457035c4705403f000140300001d0004c00030300001401d00c0001013f000507300c0c000c0303f00001113f000170c000073710cf0311c00040344400030c301000075d0030c403f3004000c7000f5f0d30d00001330f0034430c071004c4013700000004143504d440c0004cc30fc5c0004000c0c00cc313000c13500010c00704400ff433cddf00010000151c51433040110330001733f5530c44040370100110f01c7f040003d000ccd3100c0f340c30304d001c11c00035000010d37000034003030d44000013c4cc505304134710c01031c3430c0430cc10450135fc3004ccd40d4c0c04c04000fc000003000f0d3c0005030433307c07003014430c0103404f33d0d0000c0cc33cfc17cc03c5f030335f00c3443ff0c003000c03005c003c1300004000044004c000000c0400f10410140f7c3370013000c4350d10444003100fcf3d3d300d300c43531440d5000c00c01400000041300404c0400007000c430c000040000c13004001040c00dc000004030430d71000030c4000010000010304c0cc0c00c101df1c14c0401f0043003310040400000d0000cc0c0007041c343c00c00003043c0401000f40103cc104c13300f0c000130540100c335c03400030004433c00c40000cd410c0304d1347131407c43103c10345f51f1154000000300f00030c0d430044c0100000d10c4104c004004c00030014170cc71503c1d0cc4c4cc04c00401300043cc540003c00d100000c00c34c003c1d0d0311030030c0540c14403d410701050c51d0007d0ff000301015f7043100f00c400030040c50004000c00c034cc50004f00744f0000400310c0c100340374f1003304cc01305705031c500030004c1c010c0000430007d001700c4400404440dd0cc000500c41f000c7313c3c00c15cc14030000c4401000c10c33040400030400443f100000c1103030004100c15f0c01000403440c0130100c0c0c50004107c0c30400070c100034401140dd00fcc3130cc4c3003000101453c010301f300cc500300f0171cc004f500c50030c30c0033c1c07003000d5007003005434004000404c4001fd0414033d0004f43004410fcf30030100044000400c301000c00c00005000137110df0c000000;
rom_uints[598] = 8192'h740c4c00fd3c0430cc00f0003104c00010003c740301fc4100d50c000435533030f0140c4c130000513330000000c503f0c010c47000505000004c000040c4304040c0005d0c00304000f3c4030c0c0c0345f03c7011c00000c174434cc501301000c430f000f41003f00140f03305c750c004c01010c53004c0000c100cd3000041fc4c00c5305c00000000040003c00010000000307f14f040c70101c0c0dc500017f0f0011f0144510331c03430d40cf04d00000043cc000c337000010040c4030c0000f0400031f000f430000151000ccd40c0c000300031107310f40104ffcc0070044fc4730c000471f00030f03100004cf50100000034043033fd14d0003c73000c50f0341000001cf5c070f140307000001030f0cc550c10741f00f7c053010000f730f030100f0c707044301000107010405c400000000cdc1000104c4341001030c0104cc4341310fc10430030001cf0c01cf0fc43d0dcc04000c000c0f034057144414030003cf3030000030710307077300040fc0fc0004c0000d030c0f4004050503130c0f0d300c00f300040330c000c5001c31050c441040030014c014d330040c00000544c3001700000cc0f07405100c1000014000cc05400545300137000c00404c1003c001000040040f00cc4c411c0c01f30f0f01c00dc00fc44503404000017f0004cf0007113c030cf070f0000f015100cf0c0fc31c010350cdfd01310004100300c101c1034f41c00f1c0d0307400c0000440d03c0011cf40f5c04cc00010c04040030c00f0cc4c00410013101113cc334300f0c75c03c1433000403000f00000403f400c000c10000110c0004d3007f40c05303430c430000453c1301c3071030300500400c0003c31000c33f07dd303d00001c403171c3400003700ff000f03f0fc3cc0c451303401c030340000000dc040005070cc007cc0c3130705fcf0cc40f000f4c3f05c0c0050c000730001fc40100340f4004c00100000000140040400cf400cf3c10010c04040fcdc00f0f0f3011000c00040403cf0cc110c000070f4000c0004c031c54400c03040105d00ff143004f0333c0010fdf000401030004cf4fc4d7d1cc700d3410030005000000f1300000c03004133ccc3c0104c100000fc101307c070c7110c44f400c400c040401700310f055c0c100c0f30c700040430001d300000443cf00000c0300000533c01003500043100c40030f550c00050000300113030c0501cc0304cc00010c0c0000c73cc4df00000044cf000034f50f4f001343c00f300115f34c0305c0100f043c0030000c051c1ccf0400034450310004d0050c3c04000c0c000000000f057c0f00037c7c3105cc0ccc000340cf1f0c0000cf0c0c5004c03300cc034340c0c0440c000305cf40c0001003031400150f500301000c0c3d04f0513f010c400043400;
rom_uints[599] = 8192'hc0000000343c134c700c1534000c0001cc5f30170c0030070001c1000114310c0010133443d300100f0004304400103dcc30001405cf340704c10000004407030003c41f0c100410100035d1f3103d0c040010c0417c04403734000404d3cf30303c10570c10300c03457330c10103d1000d0013c3c00cc1000000f434c1010c0007c030000f03c0710c100cc00010c10dcc0c0000330cc50104040100000d0433c04003310030170f0c0045010000d40355440000000c05340c0400ff0c0000d30144040010cc10100033100000430300c40500130c0003df7000c004f50c0010c40104030440040004004500cd310c40030f000004c00031000f000100004c1400130c00300000301c0400001c0340303c3000d0c00000050c00f300107c07403500000fc00c04001c770c140c030c0f1340451003700c300cd000d31000c4c50010310031c00c00000031100c100330050c034075451030143401040c0000034c11000c0d4c004437040000340c0004001000c4003c05c33f040c0c3c00c01c01000c30c4000f040c00c0070070d4040303004004100414004430144501cdd40f700c4744000d0c0fd30304070003107010cc104d000d0c143cc40010c301070c0000707c044c0714033077000100ccc0c04c333c0c4300340000433000003010340303010734000f00000041010570001d1400340f0f05040003041005f417044400c40d00700333031f0c310101001050cf5c00c400100c0c4c140c0f000000340040d4c00d04d07144c4000c04d30c000c0013cfd00f0c0cc7040ccc70dcc117c01040000300d470cc04740cc0300fc00313000400400c100401400c0dc33010014d033c00030010040c0001073c3000300c01c0c3431000003d0301300cdf01d30c10004711c1c0ccc013c53340003c0300300034100c344c733717400c00051300444c041003c03fd4000c030514f03f00440100f03030c100ff4000dc00f00c0000cc00f0300030044cc0330141fc7101130cc30000410431030c110d000cc014130f0c34000c0c00400540dc0003d304c30c0007003f10d00404010fc4c03f43300300100004f3004004031f3031040c000100003401043010c33043000c0314030001003400141f043c30000473104c0304003c040c0f0007001f00040011000c00100f130c000000404c04040c14403100030003d400d0400714000c34407304000005000340f100f0000f0c031f00100003330d0014cc030c0c3c00347000054c003d000004cc14cc70340c1071000cc70000003f00f0400431cf0407c00f3f0001000f073f350d300d001c00c13f140c03040100000c0000400000c53c10fc0107100400fc034107470004344c03fc1000c4d5cc340000050000354004cd4404c0c40c1f000cf00d3f13010c0c100c40000cdcc0140fc43000;
rom_uints[600] = 8192'h33400407404c0011000311f0f00303ccfd040d40007300c03017c00743014000f700331010d001030dd0ccdcc003c3f0010070fc40130d04041f0470c4014003043c1c040000001f0000d30d3000f0000c4303c033040110110007700f0403c0037343040400000004031c300f3cdc3050004c03000000300c00c1d10f3040010cc340f1c01004c0c0300f4300111c0051c000c000c350c34300131030343c144300c3070c00733c0100c43003cc0030cf3540000c0dc040c100101cd540003000c4044c40003cf0040c03700000740300110c300437f0000714cc303c3003d0c0c00c00c103c0000f000f04070fd30c000300300cc00400c501c3f0000000c0030f000030c5c034c433431c1000c0040f000443044c0001c0d00c53407d01c1c44500010300005f07c110030c01030014100544400c400300330003170043c00c30c100c333f7c14003000000003cddc40c3400441147c00c0000331030f0100033104c1cc30440043cc0070d710f01100d10f00d1040c50440344101500003c0430ff4f700000c40404f0010015f30d1003307000040004131040cc73300cf1c073001304f01f001c107033fc05f007007c330040073000c0d507100c10c030c0304c00300c000ff3dc00450c0030c1000000033c43133c0030000fc17011401043cf000413005340130030c00044d100011f1401d010300f000000004454337c533c03cc404c31d00330c30f4c04300000c03d0437134c0d134110c030440c01dd4033c0dc0c100040c00400300cc3771300140500f001d050c0c0003c10c3574c0c3000c000031c0111c001cd3f34d70c000c03cc00330c0034c000d534030dc30cfd00d000530c7f0c10314410cf1f700c30301c330fc04c000710300300330030001000070c0d130053fcc30044c33030c30f00143013014010030000d510040040300d353004c4f0cc0f00cc0440d400000104c14100d17c044c04407300c7000000f0710004c0c40033c04c0001343c71440dc070c430030c40d000cd000300f0000050013c103c00c3c140005004f003400030000047c0cc00f0003d43040440010030300c4013044330101703cc3f301cc104300030031c3c4401c3001c000311007300cc0c10703000c0ff0d414401cc1c3001700000400440cc300c00100004444ccf3d04033c305040c354400f10ccc01f5444040cdf001000310014cf0040010101030040cc400c704c34004004fc30033c0c0410d0000004cd4cc1003704cc34dcc0001400c04cfc00030f3c47401303043041404c300403c0743c40d40043cc0004c31040030000000333f0c30040403004000030c00140d07431700c0030000000c00fc0c0c0cc100030c000100c401cc0c4405440300000000c00c00500030c0cc00011d00010f000001c001101030d0c50040000030c;
rom_uints[601] = 8192'h101c3000f1010000411304133fc14c0f1f0cc0c34004001013040c0d00f03013c00000c04c0d0004010503004000c403334340f0005dc01031fc0c000711440311100f101400171c030000cc0400001014000000f4000c3104403343c030100c71331cccdf01070dc0030f000c04c704000f00337154c037004430c03000130004c0d3000c30007100cc1c0730004004003c70000010301cf0040c000474cc000000440c000043cc00450013100013030414000000303030c1300074700400c03c0c00c003ccc33001300000311430000c4ccf0cd00050400100404c300010105f01030140501013000c07d435440c7005c03035d00000d04710000000310014001f130053413fc35c403001330d105010030f01431100300f030433c1f00c3103300f003c1031f100511cc0300f1444c00d300c00040c300300501c5d130d301c0400cc0100034043003c00004503c00c5d0055703310034f001000010f0343040540cc03cf3c033c03c0000cc0000c030440013700cc0000c1c30c00307003513cf1001c44530013330c00770044041000c01010000004030c00173110c070c030c0030410433f00030c010710373ccf400704310014044c30000c1037010f0c3101000000000c10d40c000c0003030f43003334431f100430c03d030cc07d00c0c05110003104c00d433f00300017450000100303001c0034000cd010334fc30000c7cf34c00001130f0003000c0f531003370300135c1f33c03c0300400077300f304303004100000304d4033404000d00000051c011c1140c105c0074cf43c0031331370f40cc1007003144003004f0c300d10011c003103031070001000c3003001300000004cc101013000001c0300c404c110000700d17000f130cc040fd0c00400000034303cc05d00c000c0300033000c4003000100410041d00713545f141300c3000300c1340fc03000cc3000cff000100000f3703d310303003010014000d000005c70c00000103300d03435f4030011704cf3103430c31340003000000044c0070001050300c3703300000fd0413c03000003015030300c0000000f0051030300001000000c403000005330c030f00000c0c5c4c300030003f0c1c00340110540dd104043301000030704c30cd0c001410f0fd330c00001c0f3fcfd0311001d00700303f0013c307010000100500140334000cf103430c0f100c10333100033040c3740000c0014f0401000000015f53f3340300101007c50574000c34c000043000043034470101d0cd0010f0cc715300dc0f3001430000040f0c1dc00300110130000c00c0330413300001f00040c130010003000000fc433130033100145f0c00003000000503001000c3340040017c400c040c00000007003010104c3c00c4f03410030000303004100c34003c034000000c0000030004;
rom_uints[602] = 8192'h4d14000c30743004005401107100f44dc54f0000f40100d0003400000301100401c0cff13047100330c34000034011f1350c30dc7044074c0050c0d00dccc050d7300304040c04430000f157f50011701400c304433071c033cf35014c4413c10373f130010c10000cc3c0cc10f0c03300100fc103d3015150110110f34000c0c300c10040f40005100300f0000400500c3c000000000430010000101ccfcc030000c040004f50f70000f000c3c3400d044cc03300034cf010c01001fdc041c030d04050c300001001143005033131000010cc5000c0c0d04051110011f7000404040000040ff0400010f771f311d4454100300d1003004100405000cc3000300140010c01013043f0000c10000140303cff0701c330041c413031c03c334107c040010030141074000303000c1f10303000010c0d000000c000004015010445c000745500f0f114c30334f34d3c1103c05103040430c004440430cc034cd3c03033c110c0001100c3d1304c0470000c00c0c3000d1350444c00c00403530c00000001c1c300000010010010fd10c3c10c0000c30ccf71007cd3030400100004f44cc1c0100040510000300c4003f4f040c3113d100000104400c0f303f10010374f0070300c0070041515407d000c740100000f04007500c114031c10c001400001307130c340c34100430d11d041133c403c10f03300401300cc305c00c1ccc00c110103d00410000f000100d0c0c010340fc1d0c0001005d055041f100071443c434100cc011c0c00c37cd5c3c14071cc030000145c31004c40005430c1c3303c031100c00001303d40131033d30000fc01c004400010305c1c040cf7105f170441f40d031001011d450303000003f050313314010334c050c300c3d01117c041d304000000c31001300000003d3100c3d4304d000cc3d030d3000434304c041003411040dc0011414334410000cc301301034330033137d044011001000c00014c404000000010070010100c0d01103033c3f43dc00c00f07cc401c40333100000f07c0000c00007300040037307141003cc0010000011d010f00000c0c4444c7d0140000033f404c031c300c40ddc1037c004500340c0c000d000c34000c0c100004113c134143140300401430305040000c0005304044410403c101d00f41500cd0000310040c040330030f410cc00443d3c33c03c1d00000001103c500110f0c001100040003030300d4001c170131c4dcd00d1d1300c00004d1d3130cc1043131410cc303000c4101140c4f00c0f40d0c0f00c4141013400f10333c4d40000507cc714dcc00410c003030411004051303100003500c00300c000cc000071d0005c0014f0c310c74000c71010034007c30010400cc0c101c00c30d03040cc4cd04030d01000737030104dd040fcc0003000c0ccd00001001073f33300;
rom_uints[603] = 8192'hc51300043107007d4000cfc3c4c50f400040300000103f4007c13101d00dc0f00c03001374300000140c0f000000c004014c03f075f0013100c01c33c00cc03704c0cc404f303733c00f33f0000000000c00c304f3d3030300000c0f13f0073001f3d033037cc343000cf0400d300000f104007cc1c03000c07303300030ccfc3f40f003c00040300cc00c04f0440cf0c7100c00010f00070d0cf44cc1000000d3cc04340c00c3000c14004ccc3c300001011000000fcccc33700000c0c10000cfc04010000011d471d0040c0d01c05030fc500340457010c0c501030c30340f40000c507c00400001c04c31c00dc330004403404fc010034c000071000001033f33004c0c00130110000d00d40040dc00d04503001000433ff0c1100305140041c0000104010030c30000010001cc140f040d031c7c000300030c003f40f3cf1000110f14f3040c013400d450000030d4c0011410003d04c007030501001300d30701003031030cc00c0c17004011000000404040c303300430050100d10ff514c0f4003010100430d0000d5000d3c350c0c03cccc0307300001cd0000c0d00c31c70cd07003c4000000000137d00010c000ccc300033030c00043cc301d10340050c00c00000c343f4000550000070d0000c401f05d550100000d5cd000101000403305cf00000330000000d000111c01ccd1510741003cf0c40334310000730004f0000c444100cc01f0401300cc03400501c5000d0043dc4d4d100cc111033c43c100cc0030c0000d104110c00000ff030031c03fc10000330301000c40c5dc10000cc17f40000100011010c140104d030400d1f0301130040c00000c00cff33000d3351000043374003f000ff400f00d0c003f3c700107c0331070004f0071010040000010000100cc0c00cd37cdc00d000dc000c30033d3070100f31040cc0c0300fcc3037043003140030301c34c300000dc0cc00310147000010401400cd0040000c000010cc0004fdf11300c0041355c3004c373d01014d04300070c00300117473c3000c0101317fc0001500100314c033110040c0c000f400000733c0310100300c0110000d504c0103d34000c111004004c000cc00c003440c0c40c0011330cf01000131101c0c013c00c005143004fc033c14f14f0c0113c000c040001010c30c40330130344000c0304150043400330fd51101300004c04c003030c14100c330070104005000030c0410c33d4503f0000dd0000000030710103f4310170003c1030d010dccc0047c001fc03cd5f45cc5034c4f0000cd40303031c0004c13010c410105300003c4c1f0034c3cc7300d70011d01100004c105003001d570cc5c075c00110107000031c37c00004100c00d4f140107000004c00c00004005f03c0f4000330c14c04d4004c001001d00dd0357701104f00011000;
rom_uints[604] = 8192'h3f133700c0c500100c00300c001c1070c000000410c0c03c0010d4000c34dc4000f0c00d30004030004400010400c30d113cc03307040fd7000030c00c0400103cc0000c30f000c000000000d000c54700000dc00cc01000000310d004cc1c04050004f311000010001c13300040c034000c3040400010f0c040c1cc10300000d003300c00c0003400403434c00000c00440004100d0f040fcf3c04c0000040400030d70c401d0300104000440c404001004300000703430c00cc07cd0c03430003c0034300c700000cc00335010cc00c011c410c00c1f0010000140c4f3005030010cc03004440000dc00d300d00041c0c0c0c101140000404000c000000070dc001c041010cd0340c0007d305c40d1304070101cc7cc1c30df003350f47000c0dc0100f05cd0700010c4030500c0001cd0143431f0c400003000c74103d0005700c00041470c00000c1000f00d730c401c304c0100004003001134c00003550000d10000003cc0400434000c0400dc044404010000d00000d000c3c0f1c730f040c3401030f4d44c0000c00c107300c00000301000c00014330c10c4c0303000401000000000304c0000000700c0c03700300730c00000c400d4c0403cd0ccc3000d00d100040400100070300040345100070475304cc00030000c070040400100100050c0400f0104f000000040001403cc0d00c0000040c00cc000c44cccc000103c4340340711000c000f104050c704f40030000c101c30c0fc100c4300300c3c144c044010040c00000d00c13033f00404c0d4017414443000070000cc10073310403c0000c4cc0c05f040405040001c1d00c40cc000100000403004044000000ccc0001c000f11cc43000d0c030740c300c1100c030001000c70c000c003074000c0370004d43105c00c1700040004000000c000300343c0000403004114100f4f040411c13d3071c400d11743cf0cc000414dc01c44c00f001033000000c04f034001c005c0400f1003070c03010103030ccfc373000303045c0000071000c0ccf1003cd0004c00c704034000c4c00001d0004001c3040014043d40000000700000130110c04347000c100003400f0004c011404001300c30070c00044c0000404740c045030100410100000c04000c01070304100d43c00c0044c001c0d1004c354c34d30d0c0c034000040104040c000300c00103400000c0cc0000c000f001300100050c07000f0000110d4c500c43c44001c71d004100c40cc34cd004c3cc400130031000d004440110c04c0d45004cd0030000cc43003fc10c015100300f14010004000d0c0f440c0f400fd0000cc1c1000000004003c0cf0001c05001dcc015c330c0070343c4500c30035f4400004140053c0c03c00114044044040000cf0413ff7f40030d3f00000c300d05040000000cc30300c00010000;
rom_uints[605] = 8192'h3c4000cc01343000005c110cc4c1710070d003c0c05d55d0031c373c4cc0c0700cf010c00440000cc0fc0000000c40cd3cc00010c00f1c030054300110f0304c7d03100000100130c00d00304003003030044f30300c3410004dfc0410535cf30304c33c3cf10010001c30cc00f0c0c00034f3c400c300c00c00c01115400c7304c0010430000c400040301330447017d43000000000100c3c40d00cd045041400037c000c04cc04003500003cd004534d17140000c40000c3141c3cc300000c51300cccc004104c00000453040c4f0000311430007cf4033cc000010010000331500ccf1400400cc04000304413c400c37000c044d00305000c014c3000014051f1301077f000707300c3ccd0ccf00cc0070f4fc7c70001c00013cc0c5370700c000000cf7000103000504c00104300cc310cf0c001d04c3c000cc0500014cd00355c73fdfc33740c0c0cd0040040c4cf4c4414cc000f3df0f343000cf004533c43000040d3d040413c05000003500000c101c10c404c003dc30030c0d3c3040400fcc170f4300000300007c040340000001f0100c70400c0010c440070d4001011f035dc3000fc04733031000000c1400005dcc3001c00f00700300003000000d7d0c030c003c13340300fc030300003003011104f440000c170c03f010fc0005d33c440501d0d0330ffc000c0004d0000c5f0c3c454410004033f3000311170c0cd051c303c0c30d0000c3c7c01003000041fcc50410050c70104133014175404c03cf4d133000c001010c0303c0000110c00c1f31703c4003c01003cc130c003304c0c100010c35c17d00074507c000440134ccc300f01f010300005d0c070000014c034c331043c40cd10003c1cc1c3fd004c005000c07010c004000040374407737014c710051ccc3040010cf00730301001d1340040f0c0003c434003d3fc40fc0c30fc000004005030310f000001000030dc0030010111530140040310101300c005f00c430c400100c0c10c007430000040c0cd041f1700f45010f41000503c1c30c410410c00c000f40013440411000400000071c45c0444030000000000403c1014305037300c40c4004311c0000304c7c0c4d140304303ff0df10400004004c050c0004c414001303000cc0cc0500c33d0001044c544f0000c001330340000410300c0ccf0047cc00c50c0c04350331501507f3310c40003c430143c44d04030040017400070400d4010000c000000003c00044000000c5404103044c0130003c304104043100040f03c04c30c3c311c100001cc340040c0c33cc00c0400f17c40f003074330400043c00440c034f000c0d304fc0000c430ccc0c000fcfcc01dd0c00003c004070004303000c0f00c00f000105c300043100cc0f00074c33dc0c140434004000430c0001140f04070cc00f3310c0410001f003;
rom_uints[606] = 8192'h1344304400004f5c00000004300730500430031c74c4300000107c00030d3314c0000300414004007f5f001c340c0cc0d01c00034000cf4000003100c05fc0003130c130010000030001075cc0c303034000144f400f0005c0c04f31000c00104d0440443d00540000c400000330dcc0001001314c070c0013000ddf00013310f440c0104010001014000c10140004d0d07cc04000fc043000c0c303c31111c00030d00033410000303300030c140c4007110000000cff004c00000c10d003d000304050000010cc0c00300004030c300c01c5003c0030030d5000001fd40c0c00000000c001c003034c031c5c10f00410f3007040000040001013040000040c44300110f3310401c0cc3000037100000710c44d00300c0000330013c4cf000000341001f30004c1100cf1f0c0001c40c000310c071003000433c7040c0d0c00330004c3000c500cf403443340c00003c040c00c40300343fc00f00040000003100c400d10301000f004011c0003500c0f0000fcc305000c0030340f3031004040007300cd3000041040040c1f43cc3000000c033000000135003f0010c1f00304441004004c000007c041000cd3f30170000cc1000000c10000000c000c3c0041c000410300440000d0341714043fc0f0034400c014070107504c00400007003c077f100c00500c404770cc7740070cc403c7751040f41400000004000400c34040010004010c0030330c013030000c000330000004f0f43cc3100414c04000000000433ddd03004dff1053000d0041cccc7004307d3c1070051fd000001ccf0cc030cc40c0000434c0cd07070043f004433000100cc0f74c0c500000013374003c034c1c00004133403cc300003c3315330000000d100005d10010001400100cc003000003300c00100f504300c403f040c33003c00c30043c100c00c0011c10340100003014000cf31300003d30000c00d0c10003030133c4c144c400c5cc0104f00100030003c0340c3017530100c1001010d4fc0034000701c3007dd000f000000333040000403dcd10103034400c0044303104000401c0000cf4100c0c100130001404033f01000000400051c4010003000000303c04f000000f1441010fd0003c000ccc0305c4013c4400000003041c00053c0010c474445030cc40034147413000013c070c01003400000030c0040cc04010000c0c544c1307000700c101c31f000034c1cc0030cd5040c1100c0c0d01003000000c0400030c00150c005100030c0cf010004000dc33cc143700403304000cf0401f01404ff300400c3c005d344f0f03450004000c4030c540007c0333d00d5c40044c0004000470410c0dd1534d15fc4c3007040303100c00075133000c001c0c0300d1000d0003c3533000100100301000c4000000c744c300147f00000144c0030100474c03100;
rom_uints[607] = 8192'h33f00040444405033044f3c130010003c7175003d700003100dc0570004c3700000034c40d13cc30dc7010443031d05d33730400443700314030000cc104f001c00035077d13340301000310f3007ccc330d37d4d0c1c0007f3034cc54303c11c07000cc000440fc001f3004ddccd410000c031c3f14f0d00000f400071440c03430ff000011004000cc0d0030400443c10700f000c01144d4c004c3dd105c3000c430704000700400100113c31070100000f000001000f3040330c1fd0f300414dccc31f4003043040010d0301400c1c0004070001dc0f334404031d0d0c0f00c340004043d4f30400100110cd440c0dc00c0c000fc0030c07001013003300cd0ccc05003fd400371d3435dccc070c37cd0f00c03c5c40457370000f043c0c003003400004c130303f430c00c13f13cf114d17c343070c04330f074000c003c010f00401033c000c040c070540c041d50fc0043140f71100014d0c303c03c3001d0d040c0c010000341c0707177c4c440c00c404cd00431c1d00350004004c1d740d0c04011330cf0400004c0000fd00000c110f000740101c000fc04105044f4c3fd0040000040c0c0070000d443015c4140005003311033c00c00f04d00450050c34073f4013c05d14330f00cd0d005c3000c40d300c0007000404c4fd0304c5050f00cc417430c0c533010c3000100cf10dd4c00fdf0001450c043071c43500c0043cc4c11cc74f1ccd34cdc040ccfc044150f3cd700fc0c703001fcd10f0010305cc0c0000f0430cd000531d0300073d30c0131f0d4c00444001310cf500040100c00100f013c030d7500100301cc300404c033c100cc0054f04cc0740504d00470fc0000c044f4c04001d000d0cf44d000d30374c010003c045334f0c340001101000000c10314030c01f13100c1fc5c5f305c4000447070010c300730c0500c0400c00c30c0c54c33155000074301c40c5cc4104133c14c110100051cc0c031304000c3100d3c0400007010c50c03341040c003100dc35c7f30c34f30c000c300c1340c07300c303d401fcc1000cfc01dcd100000c04031003f33f0f1000053003300000c330c344301030031d14c030cc301034c0031f00030dc04ccff0030c01500033cc034c0000010010134000c57f0300005c054733c3000400c0cdd00001c31405000d4403070cc4313000000c400d0c4101f7f100007f040c0d44040c0d470003000c000c0040004d0470313431400c74cc1434c30d0ccc1c0c4d430df0500ff0033101010000440f041f1c0cc3c700030703040c030300100c4001f00c000401007cc3004473d033100c010c0f4004033cc0cc0003c14000000c4cc4704704174cc0c0c47c000000d0d40c010030c03d30310c00050f00c0d04d40c10003300101710303c10343340000c00030c4cf00c101040d3033010c0;
rom_uints[608] = 8192'hc04c03305140cc010c3c00054400c0303cc0001d330040c00304ccc07400c170040dd344cccc00c00433000500104fc31fdf01071ccc03030000000007004f00400341300f04c5000100c031000004013000100d10000c445444cf400001cc0d35cc00fc0c0d0f40c40cd3c10030110d3000034d3cc000350043000c3305450ff4030c1c30010c00044007d0cf00004dc1c0c004000cc0444d00010441f31705040c000dc0c00c00010040c0170f4c300311c70d00c3fc04c0c000330000c4340c0d4047000004053d3300303f7cc0740c33d400004440007c0d0cc0004c0d3003040433040407c4040f000d04c330070100d044c403000040030cc00dfc00077dc0331534f00100037cd0040c710c0710f0cc41c1ff3f0011c40ccf105dc00d04000000cc4c01400cd0c300c0c01d0300cc4c03c1d010010700dfccc0043000031dc4004d4c41001003103304500000f43c0433007c47170c0d4301d3c303340c10044c0df4cd403003f4c050c10010c704c00034305cc00c41371c01cccd003f300c01dc303001fc0d305144c4037c03000300cc00c10c30030443150fc07404c7c400040f4000304c01f013d051d310dc1034f0c30001cc413400134733c0cccfc000310c05cd00413300cd00c70f3f400cd40f4474d43407040003440c03c500500004dd004703741d0000c104073444c001c3f300d04403470dc31003150443730314f3cd0030d03f01cc3744003fc3c000d5404cc375f0001f570000100f0cc00304fd00c0000343c03001cdc05ccfc50000cf3f11c0c00001470c0f500013030401430030010040c3000c010300cc0301010f0fc00000114d0000c00cf30000070f0cc00d070170c00f01004c11c040c005010c0030c3f4cd000c3473040c00013100010514000343343100cf00001f110040c034000c03001310c4dd304543cc40f3c0030c7c44030c3000c0400c000cf0003c47d04f140d030c34040d040500c0000c70000c00000300c300400403c40750f0c54d400003c03c4000c40044000ccd400000c103cc1c010c337c0cd404340004007703030c03443c035c0051000cf400100000c0cf00c0c0075403030040c0f70c0034300c170f0d00431c000f1110df43340c00000c0c40000104c1ccd000c100cf4dc303f3c4c43113030004007300000103ff0005410f0000040001001c03c033110000300dc433453037c30c4440040041cc051400330ccdc0fcd0010c0c333f040003c0435014cf130030010000000334300337000cc3d010010c77f413c0c0c0cf0047d3000c0c0c0dc4cc0c4f00f00c700c05740ff700c400051c000cc34131ff0000ccc30c3341433d31c33cc340c4dc0c040100000f100cc004303d3140c50d000c034744c3300700310c044400cc010000c4c50c3cc10430033001030c40ff430c034004;
rom_uints[609] = 8192'h1d701c0000f14000c704f011cc704d10310c051031000510000370000133000c00300343c040401c0c03003f1350301300030100017c3c1003000000c31fc711110034411031dd0540000c43033003c40c130400500300f0d047f0d7c3f410c304757c1c5c000310c4c0c0003004c404c0c300c00033303c4df7043703040c3dc30071c0400000003000043c13001c0700040000000000403017070007d373745c034c0c140fc3334c3000d075f300440f3110c1000017000331003c30c10000c3100c40030040c00c13034413075cd0100140c110070104000473cf00c5000d033040c00003c31c0c4c04dd0031030cc3140f0310040010f000c1c00c00005c0071000d3cc001dd0c07044c3300033c571c301004033400f0cf303010f40c00f0f13c0003c010c4c01410414d0005c30c10700040001300cc0014404014c1047040307000340000c0030c3c00d140f0031c1c330df30070031ff0300c0304000310300cc0400c03c0c34f404001501c1f0030f107c0340c07f40070300000003c0c0cfc3710c4c011030004c703d3440300035c10043d10145303143050f374034d0000001f000d00044c03c1003cfd040433f70fcc00000df000ccd0340371130101101f300043c00c40101c000c0cc5030c0c0704c10c33030f000cc00731000003c1103304331f00c000000000001c041035cc40001d10f3c303c0040f31400704c4440c3c0000d00cc343d473f30c0004c31f00100350c373300440050343c30f34100400c0c00000010c000f03014001000c4d003410010d0c00003030003437100cd7ccc03033111003dc0c07047f00c3c147014c004d310000f3444004330000030700d0074c1cfc1d1004d3110700c0c14c10c510311c00003104c0104430010c0047110034c0001dc4300700000c0045c0010f0d0fc713c34d11cdd033104d305cf30405003c3f700c0c1100033c00c31dc31000c41d311037000430401701000000300010004000000033000f70000400d03c30cc0c001033373035000010114c030f100010c1c1d00c03000701d00000340001031400040cc3001030371c4c30003003c30c17140340400743c3305c0c0c4003c00003f30c4004d7f40003105c043100c004403cf0000c30370f33000000f3c0740041535403c0d103000410010cc300340c0f7c3000c403501107d0c500c3c3707c30f4110c030073cfc01c00000347033340371000077c0100010304710003c0000141040000c100000c00000300330433d73405f013301000c0c00c00303100c3030000034031000d30333033f30c3134700c100f1430430700c1003f0000003000405ccf0f3c37303f000301000030d0f010c104311000300005d303f40030014300c3c1dc03c4c0c04c0c031040c705030c00cf03004c3fc00300100f3430004c13000400;
rom_uints[610] = 8192'h3c01100400304c0cc01000300c00c30cc304003c00c1000400cd400c1c341c00003f41070d000400c4000330dc00c140003500f3c3000037cc00c10301033000d1c14c0d050d3303000030c041000d103c300300500f00df00d34341050000051040043f003c0100000cf000000c3430030c003010300f0100c00cc50c04000410403c000c4400cc004c10303400700d0c04000000010410110400c0413c03000c01400c0f3400000c0d300f470400410c33037700c00dc000c10c0074ccc0c0413100cc300011400fc0000c7705c0410001000300041c4314000c3f31011c1f301300030c10c00c0c300004c0300c0001010700f004000c00030ccc4f0000c401030031c0030c30004d0004300c0cc31c04100000000d030c0c00070c3cd31c000fc1000540000c0300030c4000df3000c041c30c13100001110300cc340d00f0400d3c40070710004c07035000c004040cf0c030f0300300410030cc0cc005004000053000d0043cf7f4000c0173000f3c1f0400001d0f00c3003000000300330f0d30030303040330100f4300c30c040040000000300005011d4070c004000530c00c074c00000003000504073d370d040c5d3f0301113340040000000300c00f0c0c3000030c14400000c000300014001c3001001003011c00000331111000c00417007040000c304000050f0c003c0070ff030314df03040000710c003c30d044013133040c3100c0010cc7c000000c0c0134c00000100713d7030000cc1400104040fd00050000000c004035000df1040c00304d0d74c1c1070d00c00c0c0013303c0040000ccc0313c147000503004c0000100000010000413c44c000001d030c3f010000c1001c33030040040c0133c00700000c000300000c1c10c0035103cc4fc30f000f01c04c3300030000733340004004fc0030300304dc0134f1000c0c3033f04355040cc041330c030d30000500730c0000d0140000130cc00403113d0100040c05c004040c33070c0d00030f0000030c0dc0751c0c011500cc00cdc0440300000000c0130d10000c1400c3701c0d100cc133c1c03f0040004f0005407ff00c4000003400044c03d074300f000100c401100310f0010f0c41370f00c1000030010d01000c04041000400074410ccf0c0c3d4cc00cc0c07d4003000fdc0300040ccf0107100c003f0140c0331103100030000c0100310000001000c003740000c001000000400100000c0347ff00701000d7d1010001000000000104f4c100c0c30c00100d0dc00c004070004cc0070dc30c0310003c34001003c0030003043c3300c0000001100000001000100000300c00330c00cc40f47f035134300cf5c0030d300000cc171000000c0c01004f4c3504310f0cd000c0041000d0041003f0d101d5c34c0041030c4100000c000730000d35010000000010;
rom_uints[611] = 8192'hc5100000c4d5105000f4c7c0df1010cd5403c00000400f3d330504c0c0430041c033cc544f100031100000500500110dc1304c0031d4047c5400d0000c7000c000107f0fc034c000c000c0404c40c34ccc4440cc0f31d07570004d403017500040d01013d000054030407c00000c00000000041f0c0cd00000c1004044c033f31c3cc3f1004100700143117001404fc531cc0000000000cf10c03cc0310c303c500001003c03400c30011030043d007c04007f000000c1300030000171000404ccc33314c70000435045010300007700df74f03003f0ffcc00c40070000000cc40d0004000303000074000c1301130f305c1541400c300040514114100100000dc04c3440c31c0033d04c00c3014c011317004000041d0c304f3000c000c140f0044c4000cc31014cc4c3c3700000040550010f104c4000c03000130c070443003c300c40d1400143130140000500440c0c0fdd114030c4043101304150404303100170030d00300033cc400c4c11c00000c10c0004cc000441403071030c1fc10001f113105d050c00300cc3d0030fc01004c0c707c004d31f000cc5340f0c43c0540007c3c00f00000d00f04000400c13d103430504cc430073c00300030135c4000300c0c4004000313005c000300cc100c403500c04400f03010033041d4c00000c03d3c7c047003cf003001c0100301001dc43c1c1033007c00350440dccf0040f5f0000cc3003c1040f3000c0010004c00410740c0d071c4147dd00c40c0043340c30c000d30403c04c00c131004047c0013000fc07c0d040c05700500003044c013300c0030d4c471c01c3c0cc0f4410c53300c0044004c10000030130c44cf00c140003041c0d00d00c0000040311c31c0040d0737f74c007001fcd330d0c3100000303c0c03030ccc4c0040007fc0041433d04300030131f003035540000f34000f710300c0000707037c00f0fdc00070400c000041040000c1c0f71ccc300300001404c000c01030cc040000303530fd113004034004303047c4303c0003001c1c3004004c0cd0f0000440d00c00c3d3cfc500d7f07d03040004001000cd000c371043030040743c41c0044004310000450300050ff1040010c747043c000000000d0051f400004f00440c003070d041c0003170d330007000034354714703f31010010140c3c0f300f00c00010014000d01c1140034c0001d070010d4003c00000030c041507c0300c00c00040014d010003c003004071c311135004c704003001cc03111143140c0f540404fc00ccf7c7110004c3041700104c040104001040c00f00c100c440f3c103c047700001310700003317000c01d40000014f010c770cf7c0f0307d7004c4013303033100c53003c704cc4f00c300000c0033c33000003d1f005030050cc71001f00d3004c0473044404300c1031c010;
rom_uints[612] = 8192'h44040010030050c000007f400114450540000001f040cc00441f0c011f3001000c3d0dc314300040500010f04c0dcd3051c0c05004015770f030041dd0c004710300000000030300000c4001000400103000d300f00004174010f300404000000d511300030d041000c000140cccf0000430100f0030fd1031000c3c300000fd0f300c301000003c0300100c10007c0c3000000005434c10c1500d7c001d10403c001350c000c300c440100c0c00c500100000000004301500700cc03340304c001000500c403011400000d01f34f000000c3700cc100001750010d33df13c103100c1c0c100404c54c03d10000400c03004040140f001011cf0451000100c3cd00c1cf1304c000030100003310100051001011107050413310033cf04f000c1c000000011cc0c0003c404134000c0700050110010010000000140c70c010010000000d1c7d3c0c44c043040c340000040c43015131000003c0cf30100000307344010f540c0c3cc50400000000105400000000df040c00430100010403440c700015530c4c004c4010040100000000c000c40f00104000c7000033c00cd4d3f1001001013103001004000001fff3c03cd003040f0003c3cc3c00030cc13001003300003000cc400f00400001030001041041000010004004c10000c1c000c00301305000000301054030d00110115300003051c100340100f0004cc4000700d110c314d00133401314010c03001000c411f3011f130043c007173400015400003401541c1001c010350f00000d0000c30f000041503c30f001001cc0130fdc3000d4c1030000100300000340c0510540054c0fc040001d1c04330d110041404410c4cfd130100044330004350040c0101030cc00544000c37c01033314c0441c3034c00501004005d44007041dc00fcc04450057500000040dc00c03c0cf410c71400000c050f0c7010f04030001c0c300044403c04110c01400014400040f03073c00000c03000303000141500440401050c4033c1c000c0331100013010700000c33c040070100000010c3040007130007f400c3100330003c0010cf431103040c0d34043c00f0013cd001c10700300330000070040000031003100033cc1cf003010343000c7c3340f00c004000010c33000433000170011000c100410d010333c43303001000c13410c031cc00c00003c10313cf100010c00c4004000c000000d4c401c005c0310070d10003cf4300033c0c0051334c00050c44c0c00c0004307000430001c013130000430304c0304d4014c0c01141000003fc104c041d400000501c01413300cc0000003010005c40cf4001040c40007000004d054c07cc04c40047c1c00100d3c04cc0014001c0fc010f001df00f43011003031d000000100000004310030000000011510010054c000c01500c00d034104000d01;
rom_uints[613] = 8192'h30c00001c0c30cc05c3c04001f000301040c1d513c34d0000d0c00cc540d0013030c3c3f10cc403511700f001307050c3c0300111f301dd14c070504100d0030140ccff00ff500c300000410300114c03100001715c1000334030035cf0013050d03c303f000400fcc13000fc13031c010c00c70ccc04100034f0c33000c00033034330001700f0003040ff300000d1c310c300000001403d003107df00000fc041c0001000d33c0cd0001f000000f30153ff0c000000170cc300771740114003003c7301c0fc00f0cc0070c0d400c0400003c440fff0f3001330f3c013003100030030001004c004cc104501c00000000c1c00cf4000c10030010c15c100c03f003c00c3544003000c107130c10010515000d503d3c30d51303340041dd3000000400050300d1103001000430c013cc040300c03000100c001300cf300f1030301cf005010300104014111000000414d407cc4431c07334dc10103d31011310040f00053333010c30cc030f01ccf0f0030000d00030d01001f0cccc4001c000c1074035cc3c31000c1303d3ccc1dc304003f0000000fc0000f0100300d10000033400f3fcc3c0c00303100010d03031dc430dd3f4c1cd0c3140cc31070d7000d3415101d30001001c33f001300f000f043704cc003f03fc01000330300010440000d0400030001cf501007330001001101500f374033010c433010cf00f00cc0c0301330041fc0c0f01150030100d0c0c4c30d3c307300010000440004fc3c4040c001514f000410000c1043c0c340d1435c00003300c00c333301cd00c3c1c3100430000304c000d101cc00070000c400303000c0400000430d1d4c3413c13040f00cf51cc0070c0033414000003011134140cc11d37d0013c10c1030730000c01300c1001050c0c300430300334314c00100103c4f03000ff3003500301c030100000030030d43430fc03c033c4700cf3040305f1d1110c1414ccc000130cc3345f00300c3c043000030004303001030d0c430c4044f11cc00111034c100f00070047400013c000300f1040050c3f00cffff30ff000c03000fc03133000130301d0033c010d3030003c100c000335f130c00f3100000003cd10043050c03f034000c0043000000c0100033d11110000013c400704100c000103c00c43001014041c000014330303cd510330034ccc0f003d0c15d001d100c0004cc00033401c3c3c70331004403d10d303000dc11cf130c0cc3c010f0d00c000300c330c3f00f000fd00034300301c01130c30700400f0d0400011030c3000d00c041c010c0140c03d300d300c30130000f41c033115dc1150c00cc3c1c40cc0043000003041107374cd3330f7074f7010041301000000004000300cf00fc14cf3f003c31c353003030d400f00311c3001030c307f40100430431001d4413cc3040000400;
rom_uints[614] = 8192'hc03f10013300c3000c00304c14cf33c704340c0341104c113033300014f1043000f00013c330341555540501040111c107f5cc10100c00d501000300100310c04000d3c300f07103010000004c0003d040113040701f03d410300015fc103143c10330cff0f0d0140350df031001d00153f0100c13dc403d00dc35dc10440f3053d0fd300033003c00c404ddc103c3c3c3d3000000c0344c33004c00f070430c0100030043003c30f3103c100cc004dc1030df4000c0ff4413c00005131f011000f0300107c00010330c0c00c3fc111414310fc104007003403510c000c10343c3410040401043000004c0c0143c00410050734500f0000535c00100040300000f0033350f00d01004443050f0300430d5c400170000000070433017040f750033014400777033340030c3c035c440d00037f00430c04300040004001101000d03004c0d107730401304704130004444c04407100c10013c03c34c1c053514001c3d700d3000301713030103530001740004103010474f7104331c0f00c0c50c303000407340d000c01f744f130fd0fc3000300000d0d5c4041f041ccd1c433300f100c3107000000013400030f700000c04c0c0c400cf30c03110f004017cdc00d330010f00010304414004070003034ccc030400c047d3007100c3000000150c000304110ccf11d0073317f0f0001011d40400f0045f0340001c30304030ff30c4d0f0701c7c10001305310fcc4100307c333000500c1377c0500100030cf1003010d434fcc107003c000131013d0045f001000047f040f00c1400110301130034114c04133c03f047441f31c3d033000300000dd4c441c000c1003c03c334df35400103d70f31010070c03130c30040c0700c4c0c0031f1c11c0000130f710f00000040c0301043734c03730001c710c0333504403d50003cd0c01f00c004500004c4077ff3733054c1413303001500fc00f71c54501530400530c303330031730003310003c003000100100c00f3100074c13044000d000f3140350000070c007414d3470c0c10407034003cf01453d00035403c000040c0100d30440103731003000c3104411100030110001000d100000503d0cc03050774010c0074c3d31003c0310c340044001cc0400cc7307141f53000f0c040d07fc0f410003c04300c01d013700c01c030c70f3000d030050030d500001313074005030313d3c040cc0303044000000dd11300cf004033333030700c0f75131000001c00d4401000cfd3504110403030d00001cf0030133ccc0000000c0100c504d33504c5300f73010301d4c340ff3310001370470cccd0d53001c7000011303c00000130003400c4417304d37307050c3447c0311010c3000011000000d31000010000cc534000001313743400133cd30401f30dc0001c100040000334c0434000300300c0c0;
rom_uints[615] = 8192'h314d40c0c515077100f000cc3c0301cfc1c4114c7310c333c03c3f1007d0000fd0fc0c030f7744504433c30300104343c0330013f0700477c003f3000f0f000074053010000f04011000c0533c007134771cc030300c0c4f70f3f01f55033fc003cfcf00c0c0c33004001001c010f0700ff34c0040000cd0003f003041c500c3c340d0000337330f0c010010c00003d10474000000300c0101f1c0f0001c0701c133f70504130c14000000044c10c0300031573000101c03035000300f0c1c0110300311c00044000f1003c0cf333530330c300100c4f33c03030000513030030f030000cc4f1140315000f00c4300ccc5013303400d400100013033cc000000d031c000c0ccc330f04f0504d33330c0507f00000c43cc40040cf13301c1c50000000400f7300001c004070dccc003034c70d0043030000013c03c103c100c5c0df001c173c3c3407cc030000070047343f0c47304c104f433035f41c7f030104003c341000144001cf004453001030301c00031cc4c100773c310104c00c0c04c04000003c30000114000000f0c10d00d3000c4000304375500344f0c34c4d50407730333c300113007c30001d0040f11ccd5401c5c00f1ccd15f00003c03104070005f403000fcd0d3300c43001c07340030000f100c77001403045500133145457533001040f0407ccf0dd30f01c04c003cc3013040310337330f0d00c0d11000cfc1001441003cf000313407000110031743ff0c4033cd333150133407d0c44004100110054300017f0d311301c0051d450c00001d4d7441c4f04100f00c3c03c014c00c33300001c04301cc400000305043c00c40003004033c10001450031001c0cc43030154f1fdc0000000003cd04c330d000d30f3c1530c1400c0c50010010700104013c0d37c3f3d30f5031f433c00313301c303c33c030c45f03340104033d01373c33373000cc1101c5011100c0350477cc0030030000043100d471151700500000dcd40d0c0001340f000cc3344f0c04f450c1cc004f0700c4003000c000034304f00170c0031300103c000d417f0030030cdf04330cc1340003d111131f311c33c0000cf14340010004010001035f1130c0000370c01503400001030400403cc1043c500d0700d33c1400c131370c100000000001f401010000c3404c0430051cc3013c1c003000044100100110071cf01c300010033313ccc4305004373d1300c501000c0c100f00070050041300c0503000c1000c4dc3d34000f3c03030014311410135140300103dc50405c14130d001140370303fc10c0010c30510c0c070f000d1f41104030f3001300f53c001f03001c4300c40373f0010000f0034fcc33400300c100000000f4c04443004030104f00c147fc030c01005c01f000301fff10c003000101ff000f04000c030c770030fc40c33c1f1c00;
rom_uints[616] = 8192'h33c73500300401c13d0407410400543cc30144000c00014100d00304c415733000f3300cccd1000d3c00110001000c3f07f1000051c0043d0113c0000c01c00130c034f3000101400000c110f30313f1011303000fdc7f0d00c00c0c50103d030d33c31107300c303101f31010f07400031c3000cc1033430cc07f4d30401c00001dc4304c0c0000004c0000cc0c00430033000000300005cc340c3d00103000040c0403c41f3314c71c04c511704004c00df50400137c4401331c0c301dc054300c01040400071300f430041010010c00003410043d34f0000c10000c110c101c100401110cc4440007c1501103d00c0704f00f311003310cc000cd0f0000f0141c0001cc4c034dcc0044030c0373c0cd133c1000300700043300030007c4c13c0c10004030075103101110540dc00cc40304d43f7ccd0010c00d14000c070fc7c0c014cc1c0003dd00d01004c0300f10004400d43151c10c00c1d010003007c0040010433c0c0000f0ccf007004113100c01000153114d00d001040000030ddf03333dc70c003c300000400d001dd70000010f1000003150f4010004003017ff0cf0c04104000704f01031070114001730004c14100033044731000cd03004d1470411d003310340400410cc1010c4c4300ccd1d0cc7fcc340010c150f00144000c1c000447000cc1f1d0500001705100c131000d1c0c1dc3d0d0000030310c500503f0714c00140700741033d00101cc400003d0111c0c03c303411033104011cc110d0440c0301334100000030c10317010003c004070c0040003d004070d004004130c00300300f1104140d0004c403c04c37c47c41dc1c00031f0004140c0000000d3f00007030300010c500413f404330070c7c3005100c00c7000c30f307510300010004147f340cf1330cfc100d7f31cc3d0011440c400004c40101004f140c00003000cd0fcdd30000c0dc74d003c0550c00103c0011000434010033035004040000100c0400c0104cd00c14fc0f0c07030043ccc00d0000fc000c0300300f50f10cc300d00031040d150c070d3c5500343c0d1d504d03140c0700000c4000f70400d003c000f4010c44007000c000f03013c000c10c01c00c47c30050403104c003c740040000040c4c400300cf44003100310f07317301040d3cc31c00040f0c400d03501301151041000034004013cd304c0f143c40000001000c0010550c1c0070c140110c0331c707c70711000030dd0000700000000c0000c0f1ccc1370003043101f4400300400f013c3534d4774400c00c3330c00d000407103c70c0303d1030000007c4010403030f4c0f0c000cc1145300004c1c0cf40003000cccfc340130d00c40314d4114cc01c70100030ccc4d0c17c0df0cc01070143d7c03001031040c300c1c033100533c030c10100d5c3f3c0030c1130040;
rom_uints[617] = 8192'hc4430000cd00050034440c3dc0cc000d070c0300c404310100f1010c000c344c00000f40cff030c0c0cc000cc010103c140d340f4cc0ff1040041c0300401310cf1004341100c0f00000303103000350d01070c5cc0f0c444030305c0001d111c015c111dc041c4400400404500c51f0001d0001c0010054007c00001304331c00000400cc0c004340011047d400340004330030000f1133f00dcc4c4000000d001400000401174c04f7cc040c3c1c00030c5000003017000c1400301044c3004010000004000030d01f00410c010030001c4f70000d0d00d00d0c5750cc003f1103304c374700070000cd0f1dc5003c00c0173014d000fc40301000104000400c300d0303304df0f0ff0cd030c300331cf0001c0c040030f0c043310703c0c0700300001000410c017030341c40001053040c1f000ccc000c00cc1d5410000114ccc0400cd0f403173d3030c43410c0ccdc340fc7f050cd40cc433100cd1c04000f01043404f013741c0410c003513004ccc3c14c0000cd10d3030470440141f7c41740cd00dc13544004014d3d40050c0010c430000751400cc04f403cccc74c35000c011040000047c0340000000cd0400057d010c030f140430300003300313c03c0340400430c4d3c00000003304404f10c5744330000cc0000c00f1ccccf0c000f0c0c000f5001000f043d000d07130c01433d0771f100710c107c1d041c1c40331c300c00c430d000100d000311003cc440dfc113307c030470011004c000fc0543705050003040c05000000000c7300000d50404000010f000045c0f17003000c043043430f303001c33300003c740304010c30c00300005000c57c30d3d05003000014400000df03d00744d0000c030c5003cc0cc00f30044404447001004c0330000114440130d111130003314c010000c000000104101430fdcc4d00404c304c7453cd1147dc7101100300f0d0404c00440000043fcc010534470000004040c00c0145cc40cc0037430041004d0f00031c0c41004fc3043c413007000000c1ff0c00000030400400d050dc04030510c0c035c00c0013044ccc310030414043cc41c030c10ccc001301034550033303030c000c000c400c3301004103300d00000430013c00301050001001013003304443000340c300d40107000cc0140003107c00c3c011501d0d000000007040c000c300c001c10000004f0cc4fd0c0f00033c0001c00307050000304c7d00c044004c70c1370000004400300d413313050003004c3701704040040004300cf1c45c3040400000c10333d01f014001c1030100ccc07054003334130550031c03dd00010fcc101000030043d1030001d140103d30c00000c00070c0c000110000c0011005f0130c500c000001c003f034107000134c3040004410401070c31010c003c4000044030c4c0030c00;
rom_uints[618] = 8192'h3000000440040033c00003c100004033c040007000447013f4c11c0fcccc0310003cf141c0d0c1033033145140c740c5510c0310c04100300000004cc000c0c100c0cc40001040000000304cc00d40c04c30034f30cf010000040fc1000000403d0d00c1300cd0000540700d0c000770c0c0c3c7c3340c1030c04001f10300f0d01000001000300011000003c11000d140c0c00000cf410f40c0000f0001000cd140d0414530cc0cc001017dc30c01d50307730000414c0c54c000040011300cc7f0c01100c100003010030040003104303d03c0c04fd300f773003330c4c00341001000503130c00c400f100c510dc70010000514c0000000031000330041c000c0c005c113005c0f30005330c3000d310c4300007000dc5010430041400001c000000330f30c0000014003300300011030cdf003c10300f3cdc1434041c111000c013300c300007f03310ff00110015f7010d00000044d3c0010301cc1440c1fcc000000307cc0104334714000440000000000000300010031154fc140411701550f01c0030003c0f030034001011310c330c000003004417030d00300c11cf0100000513c01c0c003f0400cc303000c10117000751030f0d00301c01f1010430c00004003513013411000300030040000300400000510cc01070310cd00c0d300001000404033303c00005c5c0015f03c0f00d3c040f140c100dc4c7c0741000053110110003010000701f0d01c030d01500c010c41f0c0411400c00341100c11004004c000f003cf030000c10000c1004030f540f17430030313300000cc4140100300c000310100c100010000400c3dc013cc44f01130400f01c03140014010001314105300000300cc03c003d03153140c30c043000305003144d000c000cc47f0c00c401c0d10f000f000c00c4034cf00c1000c1300001001d000c04501503333050043c304004130c30134f1304000004000f10030f1c4403000f017f0c07c31c0000033f0f3c31000d04340010041014f304500010cc0c1330dc33140000cc0d40000c10d4300300c000003c0c010c30101003300001001110040c10341743714000c0f0050110003c111c300cd00c0041110c15141d3700303410370f000c04f40c15047000000730101400c43003000f00045704445500043430cc00c0104050040130057c0010004f000c3c003c043c01c1c0140004f403d03130001d147c000005cc0004050d00c330103033030dc10300001010047434c1043c040014cf001d105401000710c00d4c13003c131f0dc700c0003001c4f1fc3c1000c31100101154cc00010014c031130003c3c0300c0c030301040005003107003f3c3c01141fd50cc0141103313d0540d410000cc01000000f0f130000030cc41414303000050d0000000000c5c5040100c00c1000170403001c1000000c01;
rom_uints[619] = 8192'h554cd003c0717003fc7010c00001d430700c00000140140c3035ccc174dc03400430104305053010d3700000151111d0700c30c00341001cc30cd50043003000371301311c710033d100f4047c005c00c7000130c3510013411400101cc1333003f010f7f033001c1000dcc000c0fcc0103707f00c0d3cf003c0c04c1030137310cd401300300c40f0c0105504c0fccc00ff040c00031010f03fc307df0133040f053000c00004d10d10001007c00c0034401d0100000173cc001001540f0c10343c73130f1350013433c0f30f3000400340d13000dc00c10300d5f44c5f0304f303001010510000c43c30f3500c153c3f0000d000cc003c043043c07340003c0330031033c0303007171300cc30300cdd17174501d33030cc004c3c0f3f00c134134000f033300330100c031710431c47c4c410143c0c00073c144535140003dc000c0410f30300500404041d700314d3370011353013303000f73033cc4f31000430404330340341c03f04450301c103dd0d03703037000004f3313000f10014c3f00433c0d3143330f3c71d0003cc0000d1104c103400c0c004400530c1f010710000003441dc40000c0010014c104c0331d0f03303333030501303c4cd00c00c400013330000cc3304c0000741c00070000c00115114c0001000f0100035d00c004d101c1c3130cccf13cf47d033010013f1ccd3003c03cc003303107d0f041f0340c073130cf403031c44030c303c10cc00301013100710407c10303d4101401431100030400c030f035001003c034303000c100110431000f0d0004417000f0f0000001370000400401f3d4dc030000d10001c000c0403133445c4000031f3300030003100010c37004cc001dc00017500f0310013303f11000035cc0330d033c43f03040c713d010f0c0103c01717c11000c0401703c13c001103c410000d47313f04051000170744d4300c0dc7003c0303150070f30400100000ffdcdc001001000034c0cf0001c13f3103f003f440130410014c0054100031150f0f0d003313c300034000c103333733033705001fcd00030010dc335c001131c10043c10c43c0430c450000f0f0dc0000001c0cc00d310003001310000c101100307303000f13017044100ff03311000f0cc00150c440fcc03411373034dc10c1d30100000c1354d001c01073f1c443430d1003100dc3d3333337455d00010cc40110014300007000011053c5130f0c3c030500004334010f3403c000173010400073f0f4d01f00340515300013010037030410303304f300cc45003cc301c0d031004077cc31330033c00c0444cc1000300030c0c37c404d01073343000d1dc33030010333304330d10007143c03d0047043001000401301110431f00c000c003f0c4c30cc0400303c303c30140043310c000d001031041100cc0cc33f00000031;
rom_uints[620] = 8192'h143000001330101c107031003c0d7f304403040c1011c040030cc0013dff0100010f3c77007001010dcc0001c101c51433130000104010fc0c0000113c0010000000c70c0300030700000303c400000303304d03030011003433041c000003d3010f030f03030403001c0700cc0033003cc001300c1d033d0010100300700003c400730050000001000d0000c10000c14041000c00100703c03303101c3c00300d00000003c3037f00d1000c0f04000000c333700000344d1c300001c301100130c103300000300033000003000f1d0501034340041033c004c0310100110000034c00111c00031030f000c4111400033730300100330000c0001413030000003133070400340cfc30d1300003cc00700533010cd4d0000c031400c0044f7110c0040000c0df310133450f00f50011140004000c311001000000000033000004d0031000013117001500033310040d30073013014ff013df3c11534c0041000700330000000001030013031433000d0130d30040c03131030d013c03c040c000300f0030f30dc10107030333100071730100c0101c11054000301c130f0d3000013111035333300403030007004c1000304400d00005030030303d3c1000c301030000000303100c500043013100004074000003331d3d0c040100010303000d31015011400c00d40cc0c0000003030030d130500c3703000c0f04c300300c550f111415113300cdcc300000f3450c0000010c0033137103103441314d01130103110cc0c00701100034030031000000304347c001433000000400043500041003000001000000070011d00131130303030300007c0d00000f000143331310040331330000c500c3c4500400c1031110c3c03d13001031c05000d4c00c400300c0317314130d00401f3000d0110000300000d7c000dc000c0013430303110010f0c00101100300c1000300033033040400cf05d030d0d03d0050f05000313004010301f30000f10031003043c0000003000f4c4003cdc503001cf0010301003000003001c1000000001300004c0c301c301015c000030000057055403fc0c003470100041304cc5c030c034130000f70100c00001305334300c00000100003c003011031d003404ff000347000400040c103314034030103413f1000410c500001004040cc300010d00400400303400031000301040504300c10c50041c0c000010d0000000000c0030100010501330440000300f130d10001040030053104000014c70c30003c034143014535003000c013000013000100f404c5c1d0300333340030054110c03f0c000001000000c30141014144401c1c0433000000003c03001104030c45cf13c1003c000c5303733300000000c1001110000103c0000003003c0f1003003f003c55301c113c0303f300010007c014c0d40000130f033110;
rom_uints[621] = 8192'h110030c1cdc004010001f7c0c40c101c300004340c0d504004f100c5010c00003000304403c00007cf133f340030001c004010057030441ccf0f00ff1030070000c440044cc0011c00030000000f333433d04054c140dcc0500c4700003730003035c0f730c07700154c40c0011d403c03000f4001001c050000344c117000cc404d7c00c4c0014000040c743100043007003300000010430040001c0c01c030c130c4030c4cc0c34430041040c0004c34c330000100410130070f0370001c030c03c0c03004300041f000043077f0c04c3c4c3400c4130300030301d434070004000070c000040000000030301c033000c3300743c0000003000045003107000c0d5030c0c304140000dcc0473000d7cd01000c0570f03401100d4cd0033430000d3003c7011000cd100037c703c30003d170c0c34c00000c300003431c000004c10034000c50004004001d4110300c77c0c4c03004ccccc40f7070003ccc040400303f003c0c0040003cc5040040001010515c400c000331c03031000003044553033373f00000d00030035000017400c04000f005043401300700030c1c0f7cc000c104c00100030030001c33dc10dc13c00fc1043c73c0cf0f100c1405c3000c00c40000704000c0c40c00003004c037c0003c33330304c40030d30f000400c517f30034cd04c7100043c100110100000f000c430304c05440030c107c10c7c00c010c0000003c10104c00c40d4400f3cc40300d13c3000c3ccc00c03000301000701c300303c0d4d00f13003054cd301000c3df00000c530400103c3c3f101cc4c00040101000c3130100434031000f0c000737c03c04d0040c3010c1440c30003c000130301004c004c04040704007c0cc0403100cc1504430cc10000743c01f1f1000000c0d700403c0000007d3c0c0000001f3100041040c030f7c04c004c0cc300100011d4403773033030000f0000003054010c00d3113434d0f0300c0f000000d0cccc00030000c3c0000c03c331173c3cc40100000030c313c1f700400c3c000c7d04c00010101000430f4000317cc33000ccd000040f3544005130133004c4c00c000010c773430c7cf3001000470417c3c04100c0c0c40130003f0400400d011c3000700110c403100311030c30370040f4501cd10c003070303430c0703c0d0304c0c30043030c0000304f4f00d000c14c7cc30104040000011314d0000c000d4703c0c51300c3017300000c70c0ccf33f14000010fc000010330440030c3c0c3400130f30d3cc34004003440c003c0311c13300c3031003000f4c0fc7004c170400030040400000000140041d010c00dc000c003000d750000010c333001f0000cd003300c3004f404300010003400c04131c00dc5340404c10313140100434041334303c0003300c040040050d3ccc35c0731304000070;
rom_uints[622] = 8192'h3030000c0034117f03000d1f000707c45005111000f3000000f0000c414cc30dc3c01030071004f3031110131010333110044111050c41400030003000cc00f0c4140500c351003c000014030030cc410d030c1ccf1454301fd300000001000000114134035300c07c0400f00f300300040400034f0f1c00cc11413d0143700f00c100501c10c3440000533001c04444c7001c00c0f44d0dcd00013c350c0f00c00c400300705f00000c300003700430003304000c0003570301040730710c30fc0d00cd001040c3351c14003d00fc0010c33405fd00f004170000c1ccc000015d0031130330500d0000dd03313c1c0000c0c3433d001110040003400c0000c0003d0044cfd74113004010c01cc73c04c134041031c1435153013cc0cf0151c3154000d31100d104c700c11407f110040701330004400c00003430f40300410d41000d4c304305c000117f000100003c4103104001704d00d750003404f113d003030003dc000000410104000fd3d37c0001003f003103351511013500140c3f14c154130030043031340fc3c0c04c0300300cc003440400010c0300040307130017014d01100d0003000011530400c13fc400404000000300330c13300c0004400d434c5410cc043c01141000003034040401301011030073030070d3c3144301500304d3400c700431040f500030cc100137400cc4c30c3cd31300f704ff40044003000c10351cf3f100ff171c03010700033c0cf004c50300f0c30100344c44c047003300730c0000014c003d00c10c04c0c10000f003074100310411df00003370d400334100441004fc11d040050cc4c3cc30033f40f107010c33c7007c1400003f1040030030010033c000df14403d00c41c47f00cd3d3043107000c00fc40143c00070cc017cf00f3071c140c0333113c50033c03107000ff045300010f34001c40031300c0103c110cd700410c3c104013cf03f4f4340000c40000c000c43c1000310101340300000d4cd4301177c03ff0340d047d01373310300010000104cc103104c414300004303100000cc40c0d300501304c3c0c030030fc1030f03110d3140c00400004f35031f03c000c03c3000c01000c033d10d31404003c10300144300d3001010d030000100344434014c10140005137f1c30350000c417003c0000517c004040cd00c7f030004430000c00303005401000301000330050f3010000c43400000c340413c0040034f3407ffc71330030105303f0100f00413013c713f004c103430c05c00dc130c000c7f3f0c00f4c71707c30f000c034001010013414c00314040ccc3013001cc031ccd00430031130000000130410310705700403473c04040411f1c003c0040100030d050170c43cd0004300100510c0040c410100131c0f400333050103cc0010000001c3cc0c0035050000000;
rom_uints[623] = 8192'h4d110400105000c5015003d003cd03143440d0f00cc3d10740d0dc003c30c000000307f11013000040c30c003c4000c00c0100c1141040cd130510f0fc030d570140400000030351030005c7c0004c10f303c000f04fc00cc00c07f003c304004101003317403c1043d71f00103cc771000010c3000050f000f3133301f0003c734340c000c000430000000f300104014411c00000d4c014140304170713c04004054540014c4c50150101d100c303c4430343000003fcf3d0400004ccc4fc00f74f070c400c0400c0df00c0c4c0cd001044500103100f1c11010cc433c01700300300073030000400c300c4c0017c004310dcc1c34003c10fc140d10c0100d0d7404433d00040c34137314300c000c0cdd004040cc41000c400731430c1cdc51c71300000110071345f3117340300100c00114000d0c1c0030c5c0f13c043305d0cd003700c00000c0cc05105010004040c00510f0c0400c1340103d0cf3300110cc0f303c0000f00c000410140c30403030001000017003440ff01034000301c04cfccd1f001d0c0c0c000030000733000140013c04000044c100100111040c7d3fcc007c0c0404001011041000003d000040c3f0003044030004000334130c070050c110cc05034d3400003000400340c0000033f0100400c13303c00dc0c000c113f03cfc17013330d0733f3004071000c03c430c1c103051310101013111000c7004c40400003070d000000014c401cc004f33003d105cf1fdf030013103cd300003c0300d00040c300400007003d73400cd00341011454400c10010301003d0300c30304004131000010040001000000030fc50300344104cc00030c000f0540c00f0d330c100c410c0000c1c7d07f0cc0143403400c005410c13fc001c001300c00330003000314004c003005f0df00030cd740f3004137000c00000f3c4c311000c3cf0104034c43001000030003dcd0301710400403001d1410440000cc330140000000c4040001000f301001cc01c341cdc0031100c00103d3c1033000c001134000104030c0c03c440314301453400107d00c043003303c0001c0010c0c00405300733000000110f003ccc3000c0cc0300403030131000c0044c100c3011001c00c110034000000d0c101c040040d403101c000d50d131050f400c0051c400c4110030004430d440300dcf44004f10044037ccc3d03c31100d00044010000c000044100c000100d00340040031050010cc33c4014c03040ff01100cc0101400003f00c10001f0c00003ccc350100f0d4331c0540010c44cc0c0c110ff0313d0111dff000000403c0001030ccd300001c00300400c0100c000c330003c330000ff40c001004440d3c10c3c3cf00c0070c10c00c0c00c310050c3d0400011030c333cc3033050000300ff40ff0000c403000430c00c4133dc003c00;
rom_uints[624] = 8192'hc0f401104050c04700f0c0007404c03c0cd04c0143f0c1c10c03010344c34401010cc00ff5cf10100330400c0f01300035f040ccc0c5340c0000004133d4330104100401c0c30c010000400337c04341d003037f4fc33c544000503c0130044f0c0007c0d1034471c00c340010f0f1100c0c00340cff004050010d34cc004370c3c3007000c33000004d4005f30040400713c34000f4300c0c340cc1f00031f03704004c401c133f3003300c40fc10d4c4140543001000c35001140c3f03000007c3c4370100f70404043cc50314403d0cc7c11000c1740730c400c400101003d0ccc0f30c73f0004034c00f340517000010703cc5c010c0340004f0450c0010c0010cf00400fc50301300003c70300c0454000707033401004000fdf045010000704d00077cd11000cd10c1d4c43fc43403c1c4fc0141005040070431cc700c01530404000d1c0077000343c0c001000c3340c0d00c0c304ff7c3cf000cc30103040003010d1373f13dc0c04010c414034440514047100c40000f4000145c370ccc4100531c0000dc000100f30050cccc30f04c0100d0c41043407330d33c1410c00000d007000040f03cc040c00fc01100005fd0140000340040000c00c400cf10c0074c000c7fccc3040014c0d7c0c0f3405341c747c40000c1000c451701d0cc53f3c330cf00d44c4340ccd04703001747070103f03cd3cf0003d4f3131dd030d000005700c0043130ff44dcc343f3040d440470010040030530d303c15404d0000741f10110003003c0c0000c007dc50410f0003f00d00030131c00c040f70c030c00033304003c04c4c040040c4403070c30f40c04031c0407d4c01000c40000cc443f14c301000000c3c04000730743cc01430103000103c04d4000cf03331c3030c00cd1c4033003f1004c0300043f040430144c003dc000c030df00f0400430cd1013ccc3c0c333c711304d00c3fc3000430107fc04040d054440030103053000000014f001030f0010d33500000000047000dc0104c04340447c43f000035035cc03c430f000010110004037533fc000c01010cd14c5c0304ff000c0004100c30400c30300100100001004c1103330c104dc0004444000d00c4000013c0010fcc0000431c1440703515040430cd3c0c10101703703c0000c34d730451c1cc0035040c0cf1c000001c0d1c10030c17f041c0173d473c00c0004000c40000000030300c0f030030c4300f4c0c0c0d071c103404c100100c400c000001cf100110010400403100cf007f5c11000cc0403340df300c1f0410c43100001c41013f04c0100d7cdc0004403450c050000401cfc001100c41004004440c0044053c0c4d014f50c0353550c3d10300fc44000c104cc40d003cd510c1c330c0100dc0103410110300050030000001400300100f3040747330000001f00030000;
rom_uints[625] = 8192'hc400000001000c0c000c00000d0400c40d03c4030043f403c00d30003030000500353700333c00000c100333550003440c330343103f0fd4001401004f030c0f001cc44000070d453000330110004004001c0004131074d41050000c3330003104f5015301130010073734030310030700003000000f000030d005074ccc3cc4df30d040347c0030c00400d0303010c70c31000100c0014d30c00301034c070104030c010d0c100d30310d010704073111f0c300000c31033013004000100303300303300c00003c0d7c0c500700000000130000030010470031303c7f070c051c010003714000010034030010c4110c0030310c0300000000c4c03f0301000434171cc35400014111303400030104430711403500030133f1d0100311371d4c0055fc00fdf10c10310000070f0cd00310000000343000003f3c4003cd0101310004334304cd30011043010c31113f1101051c1d0070107dc00035003d0404000c00ccf300304c0c41013c04310730000d51400113d00303310000301001310c0d05c3fc3c300001c0cfc100330010dd430003d433030c033001130033050001c03700003304300c0001c3070470100c04001cccc4000cfc3000cf0d030301443d1110030100000053013010d0000c0c0d00040c0cc30114013300304011331400040407330730000404001c01301f40d0030c0c01000135040003300c30041530000333001d3c00311001031001045c005c7040c00130001101f07cf41f33301d0300c10c7330030041f710000c00c1101707c00c0f111c34c333401f00d0144c014f03f4130000034010c143d003fd1004300500004033001334c5c000c330113d0df003003c04000401110431c03303000104cc344400c30301000107c301c03c0005010401030cfc33f4140dfc334d7ff0ff3737041004000f0010000304107134c0f347cc00000f10dd3d30310100310dc100c50300000ccc31013c0004430103003000030c33010c0000330fc100dd3c0c0100101f030033411114cc100d0010000c01d00d1030330010d00d0c410043331034c10100001000c0010c1315140400c03c011c100c0c300300311c04000d010c00cc001003000d0040343400170001010330010c0000400130470000400c400c1d0101003501c7010f33cc000c3001041100300004003c04004000cff4054110d44040000403004001133030000d031340004070300d0c7d000c0030c45c30cc4143051014000303101c0d5133c01c310014010133c0400c33cd707707f30700304d000c3030000d0300010c00040100c703c50d1101c0010340000c77430cc0001400000000000031fcf100041430f004f407000010c0f15003400073011c0440443c073cd335c0000c033030000c0dc33c033c0003303c0df300f1001000010c1f5f400c0c343f000400;
rom_uints[626] = 8192'hc03cc100f303430c30ff10cc005030c03f00133353c0750d03103003000d00300043d31c1057050c004130504cd0c337c311001c01401c0031000010f000f0cc00110410401004c703000c330c004030d7f03fd7c3dcc307131001fc003c304c100350040f001c0ccf3104003d33303f03c40304407d00fc030300100003c40c0c00d0c4c445004010c000400c0c47404330000000c07c50c43c01043c00001431c10317004037f740700c07113d00701d0d05c0004143c30400100353430010030000000c00c44010300003510130c4cccdc0fc00f3fc0130711033cc0d001f0d003031003300001c030371c0c350d300c3403ccc3c01001004000c100c0004f101ff03c07c00340053304401100700015130c01130ff00030cdc71f400350403f3d00073d37000000300c15c13f033130304000041040000f000100fff50c01f0f001c100c3f0313000cf03013cd701000044140dd0c7034411d014000075001117103c010f4c3000000d0c7cc3cc30004710003d334330710cc307740f30073d4430cf30541c0300003000c03c4df5d003c040f0003103f01303c0cc140440050c4c00cd33cfc00cf00030c00f00d30334cc734f40c3300c013c305144c300700300103103c30f0cf003404c0700cc35d0401033cf10100ccc310c311f04d000c1350310fc3d100d3f4430000003350c05cfc34d003c0cdc131311f00f10ccf05fd0300c000005030f0501c3c4000c01070000fc014fff041c4300000cc0170cd153030fcc34c30c3cd40000043c7133f300040c3c30310c10f71f0000dc70fc730cc10c30400c0140000c0470433100003000331403c00c3070c04010743311f0000cfc00410c0103c03cc01c03d340013043c14c30f41cc4500001304000c0f1007330030fc70003c030f441000c07c34031031fcdc3031c004c04031434d4c10033c0351700071535f4331034000c3003700040cd004001df730000001f000010000000030cc340030c0c071340c5000340403401c00100d33034347001f00cff07d03c000003730300034403430f004c1c03300c00cc1fccd5f104130d7c0c00cdcf10170000c4d34004001133c305c0004c04100000000c00c4c4404c1d00304c450f30c4ccf40303c3100004005cd13d7377004c00300cc3c0004044110c000c01cc0030c30303304c0c1000035f033043cf334300731544c3104f04440043100c0004d533d00005300030310300d43103007d077400000fc03d11137c300003c404300550030cc0f3c0f01c0033010c035cf0413300405003c030700c3c7fc00034f410700cc5000c00c703031ccc033004400000070000047411010000171000003130001410c040100f0030014013000100ccc700157d030c00404110000501101f30f00003033c004034100000c104010040ff104030d3c0104;
rom_uints[627] = 8192'hd0170300170c4303c0450c37c3030033c0300c0c0011c70700f4110010f4c30733010d03f0cd007d500334404307403300c00c03c70df30411000c0004c01044c350f333040107330c00003004100c1407010c403734370017c4c3070004350c0411dc000001c0070307d43f0303404c1f000c730c31074c00c03434044f00cd3f4443030c0f000d0300040ccc440c5fc071000000000c34314c0404077c1f30c07c0405f311000100140007d434c0000071c3030000403c330000330c05cc00f4c000c50000c0010cd54040c04415000034c3013014043d34c000c5cd13c000370000c300300f04005c10c40c3d00051c0cc00c000700c300c111000000000004d0734c3c03c10703c10fc0d4cd3f1cf3cf400331410000401c00313c0701d00cf0cd00c030400cf00dd331c00014d1413100cff031cc40c303ddc3511411331100100d00130c0dd3c3c0d30000000330c303cf00d047f50ffcc71c1c0c03401f0c31317c001134cf540101c3c3001c33031300c73f33c3fd0f003c0003c00740c30f0153c03301c440005300340f70c00000330100cd0c3c0304074431f003703d3d0c570303010000cd10c003d5c013d04053033d040001403f000010040c00c131cc103000000044000c0d000040300100c04335d443c0cf040003330cc10c043ffddd3007d4f70313c044300004c000f4c500f30331c3700300c3c30dd41404d40307d3004004331c500c00040c010000400c035c430300d511d000040103cccf0d0073300307cc033c4c0171c74c4d5c001004474d4dc33130040051030c0f0400c0040330000d34c0000f3f03040fcd4701f404000d0401513f044300031c0c0400000c0340300033c40017443103040f01cff34c00513c010350c0073c41dc30010004440040c14047340003c0cd0c31f037cf0301004700cf30f0cdcc03cf0d05054cc03347f10dc0301d31f3041c00003f03c00000c340c00000003d33530301004c00050300400003d3330314000c001d0d400300f0f3000c140404004731cdfd0010003cc003001000151004113404700000000353037c0430140300530d05c10c41c4003c1d0f00004047000f0c001d00400713c30d000c01011330004033d11c0003070c0c703031004100003cc034373300470f0401c0d300cd400d310f4050fd004400137003074dccf1354c034f001f00c111c0f1c00034030013cc30c730dd00100c0d000111003d03cfcd3d4350030c0300c400040c0c0c74f3c70500003c0373110c4c054403c3434033c0d103000c130c01103c30003f100100100315f3c00d3400f7f7000403d70f411c3304cc4c5311000d330cc00c4cc00100030507f4003c010004040333003501000c0cf503000cc04c00070337003344040f04000113101100010000300000340cc00c14070000c430031c40;
rom_uints[628] = 8192'hc0040000334d00cf30143c7011000c007d130051c3744c1100c003c000c0f10443005474c0d331000300c044c140300cc4dc003c0c100fd174c0430030f300040100130c31000000300000c304001007070440ff10c0041004cd3c0500000000c0500c330003fd10c4440c0c040f500c5040004cf434304c004330fcc04dfdfc0407400034f00050030000000c00103c100003000010104cf051000451140c1005030333003c0300101003f700f0400004c0d10c0010073d0307c430f0041003007c000000000cc03c40000f0040cd0500440d0003f005c10c44f0143ffd001440000cdc000103050c000c45f0f4303c0000c344c7c000000030d4c3fc400001004f00c074cc34401030f0003c05003c0d0c0c000dd0403013043c000d0fc0c1000003001cc43c40310f150c04c405c4140010c304000000c50cc00307710fc410c0000c004df400103c04031cc10d0043040005dffc0d301f00035030304013001f0040c0030f0300530ff10403040c0c00400f3cfc4305307f030f43100000cc0c1cc7d03c001105c0044001000050030051000000050c0003c3f40c303000cc070c3015d3030c0305c0d00dcc0c0f0000031c3f0014440f4cd00c014c00c0c00310cd0fc0005030010300d00040f00c0c000f30c000d4000c04c4cc0330003000ff00c1f0001d07004ccc053f0104dc0000344f000401c3df0000c3304335330d150c004400043050c0c05031373f4f07031cf3004c14010f010704001700d00dcc03c14030c7000001040100c0000100c04040d44014c705040d000c333300cd4334000030001f7d04c00c000000000000500000c0f00333c70040101034143c00007d4370cc003004f000000041004c303044300010cc4300c40f54004300c00c0030030305350035f031034d000017000300c07f00007c40000000c000c404c0c0004700004314c31000710c40cc10100300d0003dc004100c10000c3534005dc3000004544001000d003040cc3000000c10050c100ccfc30c01f31303070000c00405000403c005310011000c1c0330c104000000454c1543c00c7504c7340c0004f300f3cc0c034d11f0f104554c3c0000000000c0c1300c3000100c05f00001cd043103145c44301343100c3d40000310750007cc0303300cf1c400f0313000c0100030000c000c00c44574003400cd0300043100040c00054513004130410000f000cc00010c430c04d0311300ccf43000cc3405000003343101000cc7c1100300070ccf000050110401cc300404430f31c3040040c700c3f030001dc0c4010104035f0000c0003cc10001f04cc15c310100c3007cd000001003c00001f1fc070c00c3c00c0d4101c00030100300003004c0f7010c0110034f0404c40c0005c17c4c041c01430400013300100000030744d0c0004030c0c3c1c101;
rom_uints[629] = 8192'h1301000043370d13313004003c03013f3514c37034131c0c001d3cd30c150f000400d45f00140cfdc41531400113f3f170114333017c3d0030dc0101c700c0000000cc31007100504100cc40ccc030001004430334cc0700011c4c3337c0d333003d13010000d53100fc00000c0430700d3333f03ccf00030007300010100f00cf1c11f00041307100000040dc000cd0100c3c000000015f30001c00d444041df0110100d000cc353d00401c140504fc00074c0300003cf0c0c00005050d4303cc100000000d00c40c34000101100c3f04d1d03401330f0cc3040740c31d003cf1300031f0c103000013c005c0431d0410001030c0100c300403700c0100014cc011100703c43c70c3cc0773cc0000105401013141f0f030030f003503fcd14303f300000137c015c0d43d051400754030c11f1003000000d333011d01000003010f00c30400473100d4000c0f000001d14c0f01340c03300000004f000301c00fd40c73f40f35f414305400fc1753301c140540c4cc100000040c3c000107d0f0037dc000c000000400001041c70c1c1000000c03035f0003100000d30001130c4d00100fd0700004710c000713d40103144001001003140c040cc030501c0443001001cc043400c0073000030004003c013030050037c000000003f034130730341374000003cd0ccff433031500c10c00054307010d3c040f000440004c1fc0700405d3c0f00300c031700d0000000c00030cc000100c30015034433035300074504c040141730033c3014000c413d7d0030000d40d0010407f40030004f3f0cc3400053010301dd740d004377d430117030401cc040040d70003700011001dc03c0001c0100030c03010c4c04c33370033344000f31d35044100c0310c000c0f0340c0011340700300c3dc05c0d0d07343003073d40040c4010c13000144c10d3d4f3d430000040140c003000c07331f400003303dd1c001174300f1dc0300401c3c0000c000004fc0000c71101cc0cd034010cf00010f30051c1111144300000dfc054c00000404000c34041703fd00500c30011010cf00030355071c00400f130070041140c0040334001530113303003740401410013c11003c00001445c00c00c073d4300003c00001c330000010543330c0d00000174040300df03034cc0000010cc0441cc04ddcc4000014003c3304105100c501301001344010311010cf400747000013000000f000100000040133cc01777c33c000000033000370cf5100c0c0010011c300d03c03c0c0d31c10c00cf30300004cf0f0000100c0cc073c0344047005c0303040c30fc00f00f03c100000310300c40000710100434000333f0030fc00c10405343034c4000c0c300500fc4104300c034c0c10003500045033030c0030cc1000405cc3000005000cc47d01344131d4007144001000;
rom_uints[630] = 8192'h400000031070001300407c333007ccd0033c40c30c4c41400430703301d40ccc0c0f044cd3c401000113000000000cc140cc003010c0400c0c4c1004300000007003c3d00c3010300003cf114004f004df0003045110c0010444cc700400f040c0f000100070c0444c0fc040014044000c070303341404c00d001c314c3443007000501cc1c1000c03500d5004001031443004100003304fd3000300405f0000c3c3703c44c5f00000300057dc1dc040001d00c001c0c040c0007005c100c0741c0c0000000330d0000000000cd0cc73440000fc0c734f0000f3c3c004000000400000171d0300000003035c5c003ccc40c00340000400c0040030d0f0300ccc50d0000003cd30000000c0050300003dc050c004c400100cf54000030f57300000003000f35c0040c300000c3c01331034000c003001c10013dcfc0000ff00030740d001c440d00003c0c400c00001000c004000d071405d13c1d40f03d030cd00030c30030c10011c4004704001c010c0010000011c0000cc700c0031330d07d01301fcc0d3003030d30c034f004530d00c0010c00c0103c04041101300000440133c304c1c117c004303c00c3c44df0c0d410ccd0c70010000500040c0030cc0004c000004d0c00444000000000100c00f100100c450400010c430704300c0c04cd003c141034cdf04300030c10c404003ccd1f04130041100500f000c0070c34c0000000000031003f4cc1d300000f04c05c3d011004035c13000000c0c040cdcc0c0314000100034c013300011013f4030010300405000003c1f30004c05fd4070f71044c00f403070007440d01010ccc40044c0c033d04f0411c7030c3c0c0040013700c7110000000cc0c0400c500000070043c040c300401c40070000000300103c00c00114d001030c0413ff0107c00404133c4701cc0d00100f0357303f040033d50d00070c500000cccc4f40000030c340500c0103000001000030733d400000000040100000000c10c00c30401c00cf7cc34d3010c0c043310041300000045303303043c4c0533003047300034c00400100107c3c431c404310300071400c033ccc14c00407cc41f000714004500f10040000404070700cccf0000041003f0c00f040014c0cc300d3100000c53000003c004cf300cf000400ccc00030017300700000000c303ccc100d0074000000c0c001003c1000c1cc300f0f00c004d3100075d0c0010001000c00033f30c03c00c4043500000c01c00570403c0c00004000300d11c00cf104030301004d001c34cc30000c3ff00c40000000000000f0001304d3000040100000c0400034c341400cd0c301c0c000c3d4c0007340300c000f43c0340410740500000d4100431f1040c0044010404cf00c4030000010043044cd40050000c03301c00c100001001103100c01c0f05fd100000;
rom_uints[631] = 8192'h700c000000c0000000f0007004003c30c0c04c043f103c7c000000001c1000c0000c70403ffc0004f41c3030043045041003000143d044f4c0c0c400001c00000c340c0c0071047c310030007400d400131f0f040f04300011003143444000040001c403400030004030c400404045cc100c0c404c0300440330003f0cf0030c407400003004000c003c14d010340c3115c000300004f340c440443c0040014004f4001057c0d4c00c030003ff70034c0013dcc00030c440c404004cc410040004407c100040f00d0fd000000fc00c33007040c000304c1f000400441000003c04f0004c04f010400010007003c01cc054c0100700000000340400000040000034004004c0304400c00c00d00100030f13fc004c5cd700f01431003c44c4c010300c0c004c5c00044c0000004000cc4ccc040c100c34040430003c0400d10000440f3000303051100000cc0c000c00304c0cc400dc3400140c40041014c3c00c30c00057343410004c10c10c144300000040040000303c04307000d71014c00433111cf004000004c0dc000c0c400c4131004003004430003cc00c0010001cd440dc00c0500f0c000000c30c0c40400c00f041040cc30040034000c00001c4d1403c70000c0430c47c00d0340c003c041cc3c0dc04400c10001c100010303c3c0c003034004410000003c05000100400001cff10004c00001c30300430c400ccf004403100c400100003d030c7fc30d0033410f4d00000044c101504c0104000040cc0c13470140000001c503c0044030400f0001c000d0000cc10005c0030f00400000003000054d4044c000c0c000401c00c30c004300000c00cc0101c1140dc001c3414c0000774007cc0300000703410c0330407003c00f04c10030d140400000d00000040504434340c3c04470000df04103774030000c40000f04000cc1c105cdc004cd4400474114004c0c0705053c0c430001c04c4003cd100c330330000400c00000000004f0000d0145d04100004f1d0040040f0dc3cdf04f0540f000000c37c0000c00c03d001c0140004d0044c4c447c10100c1c0004003f4000c0d0040c3ccc00044c0414c040c414004003040c00c0000400c0c01c0051f00c0c0004c0075130c0c400c07c0000cf000000547003074000d103d03034d4010400343c0000007444303000c03000014f4c0000700030300400d40005cc34f70040000c0d0000700104000c0c0000c000c0000000c040c0000070044014d100c33c5044cc00101110d430cc00000cf430044c04ccd4c4000430000034103c40c3c4cc1c04c3fc101000d04c0447c40014000f0030c00000cc001010000cc01c1c00345c4000c430357cc10500c43c0010cc0414401c43c0544f11130000c4104c05000040c0400000040c1c0000001314003c003040101c1043c4c04fc0000000;
rom_uints[632] = 8192'h40000704144c50010510300730010c133cc100000404c007003314f141cc10404100430010411c070050000cf70c500470f740d3ff70c0dcf43034407f10440401700f500403c30040005c03400040001470c0110d47100c4c1f134703c4c01c5030f3d11001cc1001370d405040013d3c03004c0054504c313f4d0c743cc00c3d07701410cd00c0041f404fc00044f373d104d3000030f41041fcf334440c50c4135510000c01c100fc04f003c30c0340f4c50000330374000c00005c30000045c10001f0133300c334c014d3d40d470340000c7001710041c43300403304c405c0000403130000005030c740044cf00005003000f0000040430000100000c0c05c04c000c315c0713400003c0d10340043303054c40503c54300f37c4c30dd0d74cc003d04000c0401c000c301310040050d3001f3f000c030333040c04c440401044c440c00c140c1d103344300c040c4c474140dc0c040c4cc00300f0cc03000c05000fc0570500001c0c401d750004010103f504dccc00d314c300011f3045403c440f0f4c0fc103400c0010410c700f4c400040103c5c4014cc0141003001cc13100045ff0001030400c1035300c3040031c34040103417cf47414040d1143400130c00c3003c500003c0003d7c7301c0000307010000400000101c4cf01f00c1f0010d04333c70010c04000c44000ff3000c0c0c70403130013c71c0c10c0f000c41005c45037fcdc4003d03f000cc40c1400030001043431f0011434c04c000c00001010c340474c340005103c770c0c3431704000030cc731004000300300c03040c00100f030f3c0c513f40f01d3c7d0c4d0c00c00100000000c01100c40c04c100c100504c400f7c000c433fd154404d000fcc10f34c4505000040c3c30500c000030500314045cc3401c4003c440f0f40031c010300c0040d3cc43000034011c400300c04070d3c01fdc01c43403cc3010130043f410d410c0c004343701400001000001fcff1c5c30514c447013033143701c00f3300c00300003003304c0c1000400c50700530000f03107c1d700040c01f44c44030f130370d434030cd4001c7c3104107104c0c334c71000cc00dc00f0404f0030f4540d5c050701c000fc3500403000c0c0401ccc4ccfc030401f0c130cd0154cc40014d403c0d0c0007d05d40c0c00fcc0100411f0c4c0fc003c0303305000100434f3d10041544410c10113f03c00f43301031011041370710071500031004044f030f03c001fc4f0001c0450c1300740c01c1f0104345030d004005c0730c470cf30304c3001c04070c0d33400c450c0c33050003d030c7c0010100150fc003140f5c0003cd1cc044413d4000c4c0d0c10000c00d3403400001005033471c001003407c3000004c400003d30f00000347c1c0c0f01015053000d1c100cc4ccfc010c00;
rom_uints[633] = 8192'hd0503c0001c041c0cd3f00003354055330010000c0015c000075370040cc300c1000733f10740000d3d03c30c04404dc014000fd0c00043fc00010000310330030153004000c00d01300004117000df34c310c14040301c014df037001410d3000f04401133040d340001107c0d151443000114500f010c400033011014731000f71c4301c00130c30dc0001000070040000000000130c45005f00c30310f1330cc37c00004cc0f1070c1041053c307400111c030030c313f0c00c0310c0000040f00c003f007751371d1044c000c343400010cc070f1c1d03c3710c30d11730fc000000fd303dc0c340c0ccdf401c030007134340c100300400030343c0000054d010000d3df31cc00c1400000003003f13505000304031300000cf0057cc031000fd00337f10c040100c330c031c0d133f44dc0c303000fc4013033034053014413000dd7d3503c00c70f373d001034c130f000331c001f00c303530000170130374f0003010f451c130d037003010c1d010c44330047c0c000105d0c003311430f43333054010010c37404c403305fd30030cc0c0c41003c00000051c0c00135fc030100541cd04c3400105011c0c011003c031c4043703110400c3f35f4501c04010703000034451350cd0103100c3000300c04d5353140c000001cc05dcc10d143d11404c00303c03d301c1304003d0c04c340f001c01310030400c00155c0c4d01140d04cd0c100001000ccd00c1c00074c00007134f1f07c14c0d011073010000cc30d3000000f000000c00001704d003005510000c04cc3d0140c130c3f00c0130c00c0010f00000c00c0430d0004001100d3d3100d00f4400000030c350043311010500c30440c31c44700fc3310730337c057300dc0c3001357001015f35414101110d0047c7501300c303fc1c10c4300400310f34050010033c43cf3c1f37f001c34f34c004c07300537ccdf0c43431d0c3dc03c30501d313f0507140dc401000030440010035cc11300300750fcc145fc0f104100c00dc1333c00000c7001c000003c031c0d3c000313d54340f404f0403d003f0c00cd74070c03001c1c013cc13110c00c0000c00c14c1c31c040310331000040f3010cc03f35cdc1030000311310c0fc10011004040043000c400330410010740114d01c4d330c3f10f01000f4004331fc004700c1c04fdff071cc1000c0310040017ccd33110070ff30107d00c07431311337003f3014cc31130403000ddff40044c40004d0c1000fc04f0141dc000433d0031c33c0400730030f33330005043f0043c3007007c110007011000070c00130053c0113007431030400c0c301f530000f40c100c040d13300c0d3c0c031c00030c371310000011010c3070fcc440074f7040500cc30000170cf317701000f01f43030004000000300c0cd435344301504000003;
rom_uints[634] = 8192'h30cc0000c303031314c00347040c0c000c004c1011f0c340037fc100c00f000003c7004103c100000000044114500100c040403cd7d500050c3030c03c00f300c0401501050c400f00001011030fc41010000000134f0401000340000cf0070111d4f0ccc30040c0c3c3c103110c3010c033017011003330c01134474c5310f30f00ff0d0001c0004013000ff04043333001014000000100133c0350fc1131c1010403010741f00c0405030030cf07f400c3fd00000c000f000c000d0d07000301cf0000331003000071c3130050ddf53003050004c303c0c0c500cdffc3c0000153000333040003003c0017f000005c0000f10050f3101040031cc1c3000040c330331010175ddf301000054d150101310f34041100c040134000fcccf3d010400c4300c100c35301f304c0010dc3fd01d100f0010104000337c1f0017134500000311344c00000003340c1030034003fc7c0c53055030410c031031135005341f74001fc43c001010c00400433111d030d4dc353000304010004c1000030330c4dc31cc0540143c3300003c100d00f0c00f3000700470103f113330033c1004c4d0c003c000130300c070400c33c0cc00f00340040110003000003034003f0104000040c0041131003c304c000c30003c00010d1cc0fcd401431013c03c10411301034051007fcc04dc3040d4c00311504731100000c13331011004300000353010400413f00c01130f03cf0104300f304c041000c0030170100300004013f070030400743000004c0404c330c4c40c71c3cc000f403003c310dc3c00030c700c03f03d150dc30300013313fc05103cc3001140cf110c00d33c110c00130f13010f35174dd40033003000037031410d500105103430000d400c0c0fc01034000337c10000307004070c100f40c43d104f034014df3304c0000400053d4300d4c44c0c703034d13c3fcc1040cc00070033cff010100c073c010c30ff00d0030010334c0010003f1c0113303f053dcc0301135010f30040c000003070010000000001301d3c1c04100000d5013d000cc30c4013c03400d100700f5000040c30340f13031cc00d00f7c0040d1c010400000c1000003d043c343c004c31000c0c10400001303c001000433c0010cc03100c0403dc111130300301300017c0001c010571c03c1400101100013c350cc430100010403131000c407c5400001c300301400d007c3c31307400001037c013304c1f030c14330454f1100000003c0407c4000111c3000c3c007103004410d5c10330c00c3f011f40d00f0d541c1574000c040d4401400c4400f0f0c300f0430fc001104403f1700d000430d00400f1c000054f0401c41f31100401c04105700c001103000cccc40c10000ff001001030530400403430043100c400001007f5cc03050000c0001c434c000c1130c111010;
rom_uints[635] = 8192'h131c00030c104050053c4d40f00dd0035cc30cc1070fc00000000c010031000010010100c430403c305101405000030f0040cd4f00000c34100400c730c33000044c11d30c1d0110400101c3340c303c50703003cc700404c00d407f3c33f3010750030cc413040c0dccc044cc334c44c7043d100030c053033c105431400300c00c5c0040c004005d00c4000540dc4cf03001c000c40c30c333011030c340340704000c000c700434000010003030300003c0300d00c0301077003434c33c3030003000104150011000c01fc103040314c0034c000c0f3034c040f343400111010000c114000c0cc0d01c7000503c4c3004c07dcf0000010047101f10300000100c031dcd450c10c3f3c4c405000300744410003430d00fc0f007cc4f743d5000f00003d0cc11cc0001531c0300c307c1c00330000f30c1704000050074c130fc000013405c0000f341d0f0701034f041dc3734c110043f03c07134100340040f3410c05c00c470030c040400053dd00030100c703c1d113c0d034000c0fc11cd17f1d030d040ccd30000040c00fc0c43cc310d3000700433003cc473003304343c0c4150d40c31c100f4031103330c50007431c0003000c10400003044fc7d14004f0cd0c107314050400fd03dc3703000c414131d04d00c70040d00344000031fc047c3004733d17374f07c1c400300007d3c0040c050040000301440001c30fc005041c07311c03004531011001000037070000400f107c014d4303477d075f040c001000c003700044400010100405043034fd33433f04000cf40005c003c040f00303cc0f3304dcf0c3df0470fcf04f114033d070000103ccc070734f70401014740c000c40c4010300003c100ff00c770c000103510107c0030104030070d1c70410d014dc177333f7d30000c33ff30d0700cc10000c0400071307430053cc0341dc4f0fff41070f4fc10303c00100ff01d00f040303c3013c00c0c404c3c0034000f03ccfc3f300cd010f0cc051c303034c30c1c70c4000d04000c00000dd00cc00337001130cc501c00c7003d040c400c4030100d170c47017cf414104f4040d04007f400cd0430031110077cd00400011d033000cd7f004000c30fd053030c7130c3d5004c3c140cc00c00c040cc40c1104d10c003404104cc0314dc50740c100300403c53130100cd140c3400004ccc0143010f373c5033131d00c001005fd11000d0400cc4c034d400040c10134400007dc0fcf00000000004f7c041d141000d1cc71070c440340451030f305fcc0340400003030403704033403100c0300c030dd0070d00c04d003300010c01701140d010411c00040c03c3d0017311110f31cc400100c011015000470c7c07000730000000cf0c73037000fc000c300d00110000004c043310400c03300f30f5f0cc0034003c0000c130010;
rom_uints[636] = 8192'h370c43000104001cc444004043000331c003073401c00540000f00c10fdc100c00c031c44f1500000000000400000000c4d0c0004f00307010c00040dd4030400300010c000100344000000cc100000300003d0c0100300000c41c4070c10000c0f403004005d14033c703c000f05430304f0300f0cd01f10fcc4d01007540313104c07031dc00c0000140f40d0000f140500001000000400c3d004040f03030000c00000030003d0c700f0033310000031f030000c3c4cc0400000cf00330f0c0010300000000c710c300030000c00cc0d1003400004430003c0010ff33cf30c0300040704000000030000f0fc701cc00041700741000040004000c10000004c00340040431130d00c7000c00dd3100005f004001100107430000c00f30f03031c30300511d00c0004d000310000740131c0d700c00030000004300050f00c000cc040000443000370100f4400011014c5000d500fc535c10c0c00304f30c34c0cc10131500d300705dc0374c34003404c0040150000410100130300004300000001c17010cf010c3c000300310003000004041400400010d300000101000c100c01f00504c0c4c10044010c000cd307c0011c101140d5004c07100c00030040cf3f00343403430001003000f00030f43c00d1007d15d03000700c3040d04c001040ccf000000304340014140d3000034300114003037f3cc0c44005c011040fd0c03c4f5000cd310400c007434c0300035500017000c4450d004003c0c4c10000cf4130031001140300f301000000330f54700301d31c0004514d0000000013033100500300400f0f04f000c310031003110040010c4004cc01cdc0c0f00c00d0000073500c00c5500503434104043033413300400f070f3340000030443c3c0f003c0000300400cc005c043cc03000c5c3c100010413000050000040000c3cf400c400430cc0c0c30cfcccc15d4000dfdfcc00001c0000013034441104400010c4003050000144d030c00003110410c00dc0cc00003444c00c00040c5000df0000010fc000304404d3000c4034f1c10c010dc5c140400403000000401c00000007003d1cc0001d00404c1401000035001000dcc07f7400040000c000c01433d0400003c40f500003010000100034c01c00cc144c4001000000301d0001113d0031c04c03000000331340001c300f100031430004300000c1c0100d00f070dcfc400c303040100c300000c0010f00cc40400c50c000400c3140ccd037304303c000c0000cc3700c00003000000d4000d00540010030c03c4c043103cc00010110303051030c00c010003100440015400003ccc030010c30c301c0010400c1cf00cd01500c15100c000c331c00700033100000c1001113df0003431c0c4004000333c40130030303100040003011004c300100f40d0500d0dc130c110010cc0;
rom_uints[637] = 8192'h300004c0ccf04101cc047cc00d00c0013030ccc000743dd1304d33c31c0700000d40c730dd41100057000031001047057c400c3cc33c00c004cc7c00070c00c0f343100c0d4d3fcc4000f04c03c0fc003004ff407cf4c003315c0c041440c03c004d4040cd400000c010c10c01004413304c0f411c0c0070000070300104c40000004447030030340010004000001cc0001300c0000070037c03700003c0c310c05050f0c33c033001c040f353030d100004dd00005d0cc4c3cd30003300cc00504d110035001040400010540c54c04070000d000c0f400000dc000000001cc34040c00ffdf4c0c000c00037c0cdc0c143033000c00410c00030000d05c0c0c0441000001cf04df3ccc0c04d41c00000cdf300ccc353000170c04430c4440ccccc0073003d0040f3ddc40001000cf0004c004ccccc34c3c0c005f010f0f04014f704104004343103c140005cd100c04010000d105c000043c000074c0c00f0000043404044f1dc34c43c3c1c00c000d100c0c031310110c3473cdf004011003011c04cc077f00030fc400033140cd07400300100c0000300104000f040043300035107cc1040400000033011431c003440c0c0144c0c00c30c40700f03040f000c7041c330010000cf773c00fc00dc0010430c004170cc430f0d3c030c07c30c0d303dc000f7000c0cc043cc17c0d4c311c04000c07300f01343110000300cc03fc0103c07d0c000400cc04450c0c3ff0c0cc313c1c0d703cc1c00c7f303d40c40c13c0034c4f0100070d330f40c40c0044404003cc0340014003f34cf007c0cf00700c0000407100030c0cc3133dd040000c400044043000400000005d010c14cf3c0c0c0d30037400c0000300700c3340d000300f40c0740301030c01010c01000c03010c0c0c40044f400c3c004c0c3c00303c07031c300cc400c0cc00cc0c30410cc011c1000104000f105fcc1c13c7030fc10000cc0000040000c10c1004000c03003003340c0d0100000d0103c004000d040c4c4430d4000dfc4300104f000cc4304f000300000cc00000040404cd0d057001c3040007010004700003035430714d3300074430c0cdc50040050474c0c0300c00000030310c33340001000c70001f3ccf04000011c01400c0000000300330c40f0003070c000000c14003370c4103053471340003134f0040114d0ccdcc030f7c0c7d000100031f07003c00dc000d7f000c000c50c00f0003cc0400d4031cc001f00005001000440054f3c0771303000410c4d103cf4040040dcd4c0c35000c0370cccccf470f3d0047400c000c03c003f1f0c400030cf01f040000cc01034001c0000004100dcc00c0170005c010c01c0f00001c0300100000100cc000410311404000d3d30300c0cc0c300cc04010010cc00c10c000034d000d4c400c4d1d0c0170140c34f31033300;
rom_uints[638] = 8192'h400313c30051d433144010141101c003044c0c404430300c4ccd503c00000c0fd3d714000040d450c0c1cc1cdc3fc43c3c03443004f07cc40cc01030000041d4d011ff400010c00fd01330000c03f0c35cc00cdc11034c00ccc0fc500c01f00407c1000dc443000fc4000304c030103400d0004001c000000340450c0c0cd500f003030043700030c03c00131dc3344000000000434043300000345304014c104c0030c04100003c4f34030400301107330000033c100c0c1cdcc00d000304f40c0000051344d75000d330410000100330000c34100c1d30dc7d0000055010d00400f130100c13000030cc0c50000c0c0f0030300000d1300043cc00030310c7140c010c003003f0d00f0010c03d3770c010000710c00c00c3340f404100ccccd00070c0001030473000cf0d0c375c70033c30010003010004c45d001030000f0cdd30d03150c17013c4c301504047dcf5041c000c7c00101c10100405c04c03510dcc1041501000f00313cfcccc340d30003f000c30001cc3340d00f01c1d441c0f00703047fcf00300f00cc07000001100417d004530704cd04c4441c303104007070000741300c340001c730001355d340003f300000c10000cd045045300403300c0000104d0d13704000c00cc040033c0c417400003c0c0c04c4c100100447c0fc0f10034140301c0000300c00340040400100001013c00034c4033017400300cd0003014701dc0000003d103077010c0d010441f0110400440007140000100c100001130000004d00f40d0303000400043050040ccfcc1000c10303d3140c0f00fc11c0d10c0c03445033c030c41104031f100040333003730030c0c30000dd0d0cc104007df030303c03000c417300d03305c40357030f4d00c03114c0011c0100100000c0c3330003713c03cc0330040c1103c00c00f1100303f000c00003cc343000000cd53503c040c0f003c45004c1310001000300450700c0001340000043030c40030000000000c0c100430004044134c033d0f005dc4300003041c0110005010403100034030401c301f3004130c03000013c0440000030cc0cc075f00003cc000010000f01310703f0cc10301004040d0d00f000400440c00073013004040503c00404c040c3c01dcf0d00d1130000314c41c7003003410000000d04040704d003d041c30c440f4000dc300c0011c10fc00013433411301300440df0001000c00004130303c014cc04001140cc1c10c00000003c010004f003330000c0c00400d313d0dfcd300cc000c0c040d000c01cc004c70f031c011d41104f40cc0000001d1003c3010cc454d3d00f0107c03000c700044f700c0d101cc5000f7170030037000010004c030cc434000000c70000004f4403707f030c1040d1010c30c0d3310f0d000fcc000000c10403f5c33000304c340c0c00;
rom_uints[639] = 8192'h10303000031300004030033cdf0033030c0000505000cd410034000070307400c0ccc5031030000c1c510c100cc01313133030100070031c0c141f0c14013101431f3303100000d0000043000100d0400130040040311c5410c0030c000031c01c13c3d03300010303414f0001107000003070014c710100003000417047301070c1c3d01070003f00001c10000000000401300c0001303044303033c030c0300010700000c0033030003c0401400035310077030030c0130100000f5070100070f0000fcc00337100700030413013cd0cc0c3c100c30030310c01300110303c000f7300cc000000c0d3001cd0101000744330404370c01000100133540000cf30ff0c00730d0c33d00100340c030013c05300310c00330d3330130113d70340004cc0000005000333004c00340051101c3c3004c1004000c03103c331d00033dc1103c014dc170100c0344cf110d047300000300430d40cdc0401715cc3303c0004f7c0503f00400c0300003400001300104fc03070040300d030c30c040fd00c70503013343c0000310000300030f74000c1130000510003f30c0030300300031003003000c03000d00003103100c0c0731cd7f0404074000040f01010f0313301400cfc4010004c003cc0130033fc043050070c30f05003c003003dc001434130d4c0131004cfc0d0cc00000510700c1400110043c14000c0000014c00010c30c3113f0c0000000103c10f031d0103cd3c0044001c4303070c0030040050330f03301c030005400f3d05cc50074001cc31000000300d0c000007070001f0000107001004d0004131c4104001f1000c1c0c001003000c110000003c40013400100303c50033410000c014cd000103c5334103305c4c000f3010f00130d33000000c000300000000003d400d300d003cc050f000c30003100730100c140c300000c00000340443141fc030cf1ffc3400304c1cf40df0c100c0100d4000030001000d10130000000cd430001000f310000c0000004001cc3d10430c013303440000000004c00f3001000105010000031313053c00000000000c0d130c0000300040014041d0fc0cd30f04cd34004000c10303c3c30504d3043ccd730f00cc00300110000105130030d0000000330500000000031003c70341034000f300334d0431100f40c100fc000c0303030df01c10103030113507010c1000c00c101000d07c0000cdc0000303011403340003044d000f11c30000fcdc1440001111000034050f373300001071000031141303000c1d40043c03fd01001101c03df500000030100000030c0743003c10140000007001011035c000100000d00000cc074440010010f00d0741c303403dc40000101000cd050040114f0403050c0003030c001010004300c31733045000001d0740030030f000c74103c1c00010004001000;
rom_uints[640] = 8192'h435050040d15c0070444c0d4733010f0f14f10040744c405001cc13000040d00000303c507010c3c00370034c50000f41c004c3000f50043f53d00044c0700001c401c0c0fc3001c0000fd10f5303f4c035000c3333d30403c1f0ccc030c000440d11303440cfd0c4f1f30005c00c03440c0701000553cc1400d30c405110f301d000cc03c0c3404043c30105cf4400140f340c000f0d00003cdc4cc0104f41c03010003000c40f0003d0353f400004000f443110000000d0734744dcc30434410f000001300f5c0000000347fc13f301c5331c3403d030140cdc733d0f700c31010003cc43cf000405010f1cc01c1f05c0033fc00550034c0f00007300d000c0511140c00f0c0001f3d103cc10ff0f00c50c0000c701c040c3d00401f400c03f10c0400cc00130ccd040340033c3050ff040c44c4010430000c0411040f3dc0434c0104331053313c01005c0050f00031f70300500103303f0cc7f105f0040001031141fffcc44c0140007c0471f0500435f5140c40400f0400450500100c1f13144cc3fcc30c0014504000c0507010033030f7c0003c000437000f0301fc0001030040ff000cc300334004540c41345105004c143d405df0007c100403c503530d00000c443470003f034044044cf34c04c40300c170371000303057f00030100403f00c0cc00404344c3107000c004c301f0414150030030311001001505403f030c110404400300c0c04010400c040f30440c770000430f030303101400333040f000003f0300c1307100000cc00041f00c000405c4003340c30050010104000c0c30c4c005030cc3071003003000043c1fcd03c3c00c4400450d4044d0f73c000f0cd004cc35707ccf0f4414df1c05c3fcc30c01d310700c0004134c33c403c47000040f003054101f30f4c05f3f0c4f300c0ff10010030000f10343f003000433c440f003c4003107f0307cc1475103003df030010344c3407703f040cf003f13f14003514035c0000440050c3c3004100000cf01051530031c3300c0000003f033c140473040c03c000441c0740043003c003000000140c4510cc4d00c0fc0d50f7ccf7c01110070000fc07000311301430c1004d000c1c0511c4045dfcc7f040fc00c053cd15040403100c003100f33000050500140c0000c400f0c30cc0c40403000015fc04101c30134f01310113c013443d1000403000040cf3d031c00c33301f003f30f110f0f00000000013d714001dc54c7c3c1c0430030f1050030f730010300c0003100d0c33c0fff073c0f743301cf003333000c1f0000c0c1337f33cc330cf004c7c3c0403fc41003cd3c40000170cfc030000c404c4c700d303dc347c1004c04304003c1304103014c0001030000000044cc3c014071c34303c0003005031100d01100030003004c55030010c73c0f011c4003700033c;
rom_uints[641] = 8192'h3dd10f03014c00c00c0000134300030300000c0004d1c10300d1f40cd1c4304c00003c40cc0cc300073c00403f00340101c0730f04431400040000c000ccf003d0031c030cd04cc000007c003400c00734110c0700c30c3330cf50f77031030c10440001c300003001104c03d040070110c043f7000c03470131703c30530cc41f473000000430c00337003fdc000f0f0000000f0001440305d30001340c03dc00304400000c4c00f01033310d71401d0045cc00000c3033513070004d04cc43c4c340d40000d304100015c00d0114300030351c30c3dc31dd3c0dc1dd0c303f313314000f3c0c0000110035c05c0c3c0314f004030003004dd01c0f004c00000c071440403c304440c104c333300303cc07431c0c455c3c440000340041c001010c000000f4100c030c0300fd0dd00000c400cc3f31030000c34c13030c000300030110c4340f000100010415cd0007001003045c3f0cc40701cd3f1000c04f13f0f407770cd1010c0700033400051c000003400114100004704cc1d100000300d0004404100434cc14003df0153f0c3000cc0300000c0c53f04f00440d403337c3030413c400130cc03f030d41f4f011471430d030070001f430053001f7140c100400000000c303d411c300003ff3010400000034130c000c0104143c1d001330013f007031c3300d0500030d03d033c03100000f01000034330cf00c003f0704f0430000001134301c70373c0310c00005070cc3c003c030d3441c00730070cf3d110d5f030400c00c0d0300373c07734c03000351f3004c07701040070c01000400040cc010013c0d031100d3000101000f04040f53c00f3014c0307f10034000401f00117c0000030033000137304005070ff04f0303110fc1305c037043c510c0000c310c04430cc0300c30003130003500744c0f407f01033f3f300d0d13001d00030401c340c0cf01c3c03c00c4703c0f03c303033c0040cf0010004f003030c4000c34c10c0053001c113c10030433cccf3c37501d3100340000404c003c04033003f0401f0c0d15f00037d137033717031c00c000df3000000c00c140404cc0003437040010003030101737100010330c1f00001c13c00700300c3ccd0000340c0cc40c105c00040400000c000dc50c031f3401043d3030040c30f03c5305000c0dc400301044c3333f1301040003031c034c33d4100001107403cd003033010c004ff0c000400d00040cc403f03300015301f47040dd4dc1013100000c0505104ff0f110010d000400300d30c0030417c0c04c0c0d04c00c1000431000d05d40c451000100041c030c0f004f13377c04040d030c0000031510011004f1373c3d00f00004003300043c1c4c34f10c00c1000d03cd3033c303100dc11c0044110c1c13d74f0304c3404d1301001000101033174044000001000000;
rom_uints[642] = 8192'h40001400040540c40010cc1375007cc17130001c044011000003000400300400037cd40d0cd30c00010c0c04000341173d0355c173504f7f43045c04370341103c010140c0d00c010000040c140c31071c4c0101331107c30f33054404cc70c40d003f0f04010403013340000104d0f010f3000003c500c40040000c4c003170140d01030c0300400cc70000c000d0040300000000000003c11df040141c0f0d443100c00045300c130430000dc0004300f3dc010000300f0004100470000303000d0c0300000c00074400c30411030d0011cc4f0cc1110d0d440d174104001ccfc4000014441003c0c10357dc4d0040c011001500010070430041003400000c0c301004444400c30015d10300033001430f3050414401140304000c1c03310f044000000113045001cc0f0c0fc00d0c4001c40303443c015044030f11fc33130d30010004ff0c0c50f74f00000f3c00141fd3400c0f300c0f000534040000400007cfc0c00430410c0c037cc305113d013704004004010303c31c00000f41003ccf0340010031c104300c010d0c43d1030010d0030004cc511000040f414330030d43003c00c070004dcf03003c0000040c0c331004000c3400133003010d370d340001015f004c0c0c0f0f3c0c1cc0431c0fcc410c504d4d3f11000c030130d30104540c04017d0413071c1c0700000403404d4c3c0d701f0100000001410c01cf33031d30000c05c00037cc04c3000d30ccc000010d0f114701300c3c4d3000033f35171300070c0c13040c0fc40031c001000033c0c0001dc01c41303400050304100011130c00c1030300cf050c0c0c0415c04100010000000d0cc34fc03d7000044131000400031070c33c03d0044c0140c034c0c3031340c00c4d17400031c0003033030c110d01130f00070c330ccd0c040fc10300000030300003444735c30c0d0d43003d700f310d01000f3d0d0333030003c10f41030f1071c30c0c00d00cc000f00c1f003004000c40150cd031c0cfc1430ccc3c0f3001c101340d00d303c3400041000c170307c03004c14100403c10400003c00010c1001000440103014d73c00c0503047cd00705c0dc41c0311140040000cd000010c50f03401103350100003004104400f0313040040d03cc0c3040043d110f41031d13030cc00c0040c4051013c001f53f0f01000050300000c0000770fdc30001cc3f0c1440130f00cf00373c000c00cc003003410100c104050001f007000c170c0c340cd10f0f40000531330cf005051303c0c30d00c00f45000f034004000c3700310500cc154c030d0000010c3304100010004740330f0011cc0000430030010f00073cfdcd03405c1c0500430c33030003dcc07f010cc440df0d1d0df30c040f0000000d0c4303005c0c34c1030d07734030300014010050300001000c03100133;
rom_uints[643] = 8192'h143140000347047c3c07000370000441c40004404400c3f004cc0333c5dd0040c0403335051700431300400570d4c30c000004f050c5f1511037c040133c4c04c047cd104fd010f7030033f3030141513d53401454cd4043c1cf005f00331300c4d4cc04c434c0313c0cfc440103f3c1040134c400c750030730f300f0c701041cd7d530000d00cc00114000d3000407c303c00000c001c040000031f0c0fcc03010c33001030cc10001c010d0033000c051cc4000c17c0cfc3134d00d414c011300001c3004df0101c4fc0d001d015f00c11100c54c4440000100000f1d01c7f000d003034c30000301005fdd34cc40104005543010c050010400413044000307c00000d00300413c0c000750073040dc0c3071cc3f34344f0070c55701c43c0010300034c00030030000104505444c300300c0f405c00030454000f04035100311c0037cd403003dfc00cc1cc40000c033100005cc031f4dc0ccc33140cdc00000f4c10330c30ccc003f37ccc0cc01004c000401c000c04374f3400030011c41f04134005c001003d3c0c0ff300fcc0000304700c374c034c00d1d10c4c0000731cc0c0c40543d07340003113cd317550c1c5c3c0714c0c01f4cf3331ccf47305cd5c01cf7005000d7c01c40030d4c0011075c00c073350d4c11f5c03f0104003343044ccc1ccc3c73304000f01004d051510403000c14c00c0c0c1cc10c45d0030000000c105d04043c0cc13c0c0cc3305c0030150100003c00fc0304350c1010dc4c0030007c01cc0fd10700c00010c740004043103d5f3104400000503cc00c0c7004c103c0107700003d3c0c00f1000f43135c30305c043413d0030135c1c103f07300f040004303fc000c403f5101040ff0407000000d3341c0040cc3001700070003007030c0003c300003c0c35000050001004004c430003d003301f3430d4100c0dc311000c00cd30d0077051c4350301301c0c33113403c4103003400504cc000040430c000330cc00140c1014d0f01100c574c011100dc0c4143c0000c00133400c001000cdf0cc10dcc0d0c31c004c3011030337c03f040fcf430000304040c01d3500030c1400034030f00311d4f01c013c03dc030004007013010010c1000ccc1301f014f0000010443501cc034d510ccc003cd4cc330cd4d343c0fc00300040c30343500cf5ffc003037304f04c40300133500703411410fc0440cf00c000003cf5cc00c0000c4001300c000100c51070c3000003070500cc041c00dc0407d010c01f5c0c0f4c3030c1ff30003f313017170405c0c0110f0f043000071004cc0c000c40c0c0c00730040001710000f014d0c5c004010fc300d500d34070ff4cfd407c044511101040103cd1430cf0310ccc50c03050c344c5cc04d10030cf0050440cc1f400ccd041407430d3c005c5c001040c04003c000;
rom_uints[644] = 8192'h30f5c003013d7304771f00003500c45d331000d05c3010070007c530c40734300170000c4c0dc03c0c04400c03300d1c0340017d3430003300c401c3f7140f301030570d00004043c0003111fc000cc0100030cc0000000303401d33003000c033f0c175d4007f3700f470c0140013030071ff4400cc10f100c301307000f3f3430140403d040003300c001c3c3004c40000000c000000c1d0000403d4401050000100000140c0d0001300100550003010f1000c0013134404000d30331700f0504000710030053330ccd0401430c0fc0043f5c0000040d04041440031d3c540404d0003537301f003c00030cdd1c00001000473cc0000303f000f1c00040033310540f000770301001c41307ccc01010350405051f14034d07cc05004d1f3303dc40000003045500140004005004c1c3c5c00070000c4004c3370057000c033c1fcc0000cc0054350000000f00c7c50015c0f30c570017d100101d400c04c7c17fc00c43d0c000c7000ff0f01c01d0c0000400107400430c3010cc054c00000500404303cf0301470c0003041003004d030040c0110c0050133f10000c13005000dc00ccc0300f400c3100f003400040430417071c31c03350370310034003c553c000000310fc430f03cf040100005140d415333cc04c13030370d400f04f0403c003c03d0107f0d1c0304c004430030c00c701040c0cc04d043304c0000f1030c044fc404c0c000004333447f3cfc030c0dc400c004310010013d30301d004ccc0000534cc0100c70c4400000c0300171c00001400d03000c3c31cc00407c0040114cc50c4010334000413730500013307c4c3c30000c3f31030010003c150c30403c3300040c400c4041010450000000010c1030101c00005c01304305cc103d7700c1f043134000fc00c3343400404c5dc030000043d0c00403c400004ccc4cc11ccf1033f405c055370513304740fd103d3010c100fc03f4100030f300010c003001000100340c0000c14cd33cc0c0010c0500103104c01434f050075104001cc1f000000c00c1003c03df04c1c300003c411d0ff00003007c0540440c013101c101330070fc00c0c700f03701c30f000000c4c4d040403003c0504d04433700c0107000c0030000410c0300f30004710353c300001011310ff0004000c403fc0100c0714543451731313c4400f040000053d3cc43c3f1044450300c0110010040010c34400500c00530c00031c14344400010000c00c400c134d4c40c300040d4c00003c340c0031045f03304141000c1f0ff0033344001c14f330000053700c001010cc3c7003303000f3000303c443c31001c3034c433000010c00c30c0400f313007f10340170c034f303c404005000010314004c3f0134400040f30c7000c0307033335dc70000435c0c00f0004004003734050303cc01040c03c;
rom_uints[645] = 8192'hfc40000400103f0030001000c04ccc0c17c0004c040f040000c5100103cc30300cc3773d377000ccf0f00000000041f0000040501404ccc700410004d0300140ccc4c1001c10c15000034f03730300410c140f000400303004c00cd41331045c3c0010130040f4c4f43000400d0340cc3c000410304c4c14010737740010d004f4000f400540040040140000340040544d00c0400c40c4c073030c00400dc0c000003337140015c400c400004740005c0117fc400104fcff70c0d000343000000000d417c4011cc1f00000503004cf4ccc440d4f041f00c05c304c0cc0104c304400030404f500c400000310f1403d034c140d5033d000000f4c0c310050010000c5d0000c03450cc0033300dd3ff4001400cc0100c30044533340003757f0c7c040000f3f301f4c00c0000340003cf0c03417547f44100010c03410c4d04c0fd004040c301d0c04370cd4c0c330d000cd0700cc0440c4dc770073443cc0d0c113004400440cf3d0c0033dc00c370c0404c40711007400701053330000300310f1330c3c00004f31ffc0031c3450c1d550004000000c304c04040400100500c3040f0410340c00d00c37733c3453f000100007dff071004010dcf0c00300f00c3c3cf3c3000040f0c050030cff01c01cc04cc005300cd1fc030c00341f0100df734c1c00f3000030cc0300401d30c0c40003dc0c53c0fd700c0300031741c130d3cd0311dcf040c40300cccfc3c414c4c75410df30c050ff01f0c313000d4fc3c0f7f1dcd03d0c700305100c0ccc0330135d00c044c3003c30770001c00403340110c00c01034c001705c5151c11c040434fc0000431003cd0004fcc03040140f7040001c1f103040d0f34073030034f750cf03030c444430c00c0004134140043105c01c703f400304340300c1000f300c0300c0100353007043c04c037c000303f04700d3c3041003410f41ff0d7c4c400030000c03030c1004f504c000fc5001010c0000d300c030040000131030000404cc04c00345050f55500000040c4d0000fc000f0c0f00457307c000300c4c0040013c447c000000c0cc31d00400c03045c0df4000013c34370d300c040104c07000501000010330037c0443f000c011003c300d0001100000050cc0d040c0401044031c001000440f003c7fc400f5c1cf41cfc344300034307101f0cf030440031133c40041133c410007f04c1fc40044030c03c04f3000000cf130410c3cc04c7003c0fccc3c4701001001013f73c1f00001004f0370c04340d4105cdf45034003f5033cc311c400307c0c10001101030c01d00cc001c005f0c40cc0313c0cd1fd0303303fc010fc000d01c33300c10cf4c4c3071d0000d075f30f0000c0054c000000f0c01034c051c3301cc130d4001d0f001c1c4fc404cc0000c340700c4037d0000f401c40030d0003f400;
rom_uints[646] = 8192'h3040400c1003330c1100c00f000000c1710030010033000000003c000c0f4c43001c733c13100000141100cc110000007c5130c0000104c43d003000701030303000141110033007cc00c0f13000d140100030c3430301113440c10003f700fc0003cf0303104104300f0500330c3000100d11f3143703010070c0f0c000d1303000c3100041000100101000c0041015003103030040f100030310403f0150104c10101001d41cc30011c300c0c04c3f0c4cd0c0000433300543000d10f0100000330310000000c03171000343001d0c3000000403433c000430cc430ccd400300c4000cd000d00011c000c01c0040733c33440c33c330014134000d5033003703f333303000c000001c1001d0000433117c0011d0053304000100040c1c31cc4340000044040000f00001330f0030301005301c00050000000c310c000f1cc07030c0003043f30000d1c000f1f3110400104010101c00011c03003703c133c0700c30c010030d001170c04110333100010100340030040031c033004011c03cd011530103fc3040700c03000130003450c4c3050010401000543003c001d00030f30d33c0331003013000d01fc130c01030c1ccc17370f000004d3000f04d0000c333c030403c0300000004cc000311f300130d00001100c01d11403011f051d0330007113fc01031dc43003c713470115d0ccd50cc0c3500c00000fc3340400fdd0c0310110000003300cc11f0d001f43001011d1c04000001c50c3c003400dc0413004cc70044011000030100030100033c100003d014003cc00430100053340300000c00d000101730307004103340000130c00010100d000c10dc1d030f041100040014003f03c1000031d11030300010c000c030300000c0115c00007340dcc0000000304300404f4170700411000cc10dd0113740300c700001303033301050105033510030140103317001114f017300100043001070400300400d00cf0300dc1c0003cd001010c000000004000c3004040f050010100d010c04c041000000f00030000100140000005030010000003100301400301014c0000c7c407030170c30004033c000077500c10c003014300040004400041c37000003000100f33030c00003000000313d030100004000cd0300500c3010c0301001100401410000311003103100c00000111c7000000003d0433307010cd14004000c5d030d0010000100301110d30130f0000300c003c1001043d1400c30000c33300c003f40170d40000f10140040f3054040001133d04c5011c000000c0101000d30000003007100501005014403011c00c050001d0cc53300c1cd0030310014c0015c03d03001c1114c0400004d10000ccc00130c1730c033c0033c3303100004400005071300000001c0d00430013430010003100040003011cd030014000d0c0000;
rom_uints[647] = 8192'hf0030000c1c430317fc304004331f303c313c003c3c000030000c1313070c033000000f7003001400c4c007033000040d370100000c313331340000001000100f10001310441000104000743300003c03c0010d0f0c030414000033000d3c01330c000133004304010ccdf00c04003354000000000d040340043c3d0010400307001d40043033f0000310041c000343150d000300000405fdf3733371410014110c03d0011404311410d0001ccc0030503c000c300045001c3c30400030040c0c0030000170031433310000c03c04100c3000dc003c170c400c3c000f0310003c1c00013307cd030f04031030c100d47d0110c30000300000000003010c00300f0c000030073541001f337010430330071dd0dc30013c30303000701c1000c3d0131000030f3ccc00301f0c03d0303310300000135ff0040c1000401c300000003f144007cf1c003f070ff10c530107cc000001010c013103010cdd0c370034300c0c44040f4010000001340c3c5d10c0041ccf010f010000303c3c00340c0d1d030070340dc31100333304c003031114d00044c0300c103c371000104101c00c43440000300c04c30070000c0c10130d0d411110300c1d053f04101c30130343fc130cc0000304c0030f300c330003f40013f0dc317070303305004c30150730003103330104053c340c40300030000510300d000c3c3fcc04d70c300001c13c00333c75cc010107111000c00c000031014104133301c0f4340df1404ffc3d0300c4d4c43f304c300303140f300d000f0d3000035d001000c0007000000c7d000114000330100c00001cc4000c300d3c00303430003300000d140c34d301400f3d3c0c430300301c34c3710c310c0070cd000cc037cd7043c03300cd143c0d340c0d14030c0004040c4c3701440013300f10f404cf0d10310d000000d0f033f337c03c003034000c0c3100c00c37f3cc01113c000cff043cc0330c303030100d1000400000000c0f0033001000700c0310110000d3100011450f04141c0101051000000c303001000133c30000100dc03000440c341400030c030cc704000030303d40103c34cd43003000d0030c00004c01001f0f00400c0043110f4dc034c0fc04000d300101003c54110c0c07000034003dc53f000005c01433710004c3003c003500c0fd3101300c3c1000cd000f3d00304030d040c00f041005cc0003300c0c0f3f017004f513000104fd3c10010c3c0000c010c400c41003dd0430400510330c0040003105d00004140f0c333f011c03001c0013000f30c1011fc710d0300300c00031300c100104000000044003d00f4f500d04c7000330000044000000070030300c3c0010030f40331000040c01001404c00f00300011101c3c3340f0000000f4310c300005407c0c003000c0000f003740c0135c133c3f300c030;
rom_uints[648] = 8192'hdc01000010c3703cc70033f1004d34140c30310c10d004400170000100340034045047144c51000c1400000dd103c700f030130c00000c7030041c01f0030d4140d41544301000d000031053c000001c11c30cc030f0d7cc30c405000f0003003ff17c044000f7400c3c543c44c173f4c3040c70110440cc0303000cc4000c01704c000013c00414c500071d00004dc107c0000007013c133134044c7014150000040c11141f00103301404c310c304030704c00010cc0010c700310c130033c3140401000c550c01c0ccc7c003d0541400c5403730d707c040c001c3c30400cc0c4073d440000100034057473c0c4f0f1fcc704700000400010044c0400c40030100003d000c0400c3ff00711030cc1cd30ccf74c00700c34000c055c30cd070700300c3f40013000c1005000003053f0007517104103013034c114010035070cc0000c0c03d0c00d3cfc0c4104030c43310c1000dcc004d13300703440051cf0343d0417300434000314dd0c00101010c13000400c01000cc030cc710010c314507403c4101c3c03300004400cc411000c40140000c44511400003c0f10004f444cc04dc370004040c30c30c5cd07f30c410d04001007040c730000fc000110034000f300c0c0ccf3c000cfc01004c7c501430340c471430f0001c3001c1f033fc500cc000d133411cf030040c0c1004f0750000003414330150c04001cf30740fc0d11c300043044cf3c037f0cc0c31010cf1000d071040c4c0043c134c000305540345101400030d040370c4000c300c00f070030cfccc40313f4001333c01003003f00110fc3c00055d7077d04f0c04f00c3030140400103c3700cc1c3c04c40404c4f000c01000301031000174400010c0300000300034c030000043004c0c70141701d007040c7cc030471403d0c30033073c0cc00f00000c004c700c03c0044004c7000d4004030c1c430103410d74300010300103013cc040f03000103c04403000000c40407c4c34000051c405050110010013430c35d4c0fd34401000330d7001f3003411c001010d003cdc7314500000c00c3040fc0517403001500c0030143003c0f03c00c570300010c03034f45000000401000c3c00cc5330550300000c43ccf03c030c0c07f400000dd5cf3703110053cd0003d1c10cd3c0f00004110300f410001c0000140334044043c00110300c00fcc10c17d030341c3c01013c1700010103c100c3f000f00f0c0003c4100c0000d70c00013c303000f04414000003c0c0d7313d04f00534100c7f0f3004000301504c0004143000c47d003504037300400d037333d10c0140c44015fc500700000c0300000050300130c0003433074d5c030403c4133003051c1d107003c014d40000f00003fc3d314c0540005d701400303007c03715000c344c300000c7040300c000c7000030c;
rom_uints[649] = 8192'h3c040001c10004471f0030cd0011031d303001c000c1000003140000714307c0000001dc4c01c5070014d005d003c03c0303003000f330f0430014c071031004000013310f50000000000513cc0007cc30cc105003f3c113f0c414100f33000011043c300000430f040cc103405ff000c070c0c1d41f03d00040c3cc11300305cf4c4f30fc47011101300c14400151004300041000c30cf074003104135d0c00c104000501401c00040f3131404130000c0c0000000000130003000f0304c03f3c4c0001c14c3cc10c304c307007c0000f1cf14003340f1c730d330030070000cc00000003000530c30005300330f140040301130310c40c00000003430001003443c040c4c0703c000f30c013c3cc470c44140f4373303c00cccf0c0cc1c5c00ff1f003430001100001c1107f370f0fc340fdf0100410c1041f01c0f00301ccc41330c330f00007104030041033030c703101014dc04c104f0d040d0303011400030303110457c30071c000000c40500010410040f4cccfd130d137000f403151d0007f0110d3540030000c53030f1103000100000400000cf3cf30d00030011033c00030004ff00000c03030041f30301c510103cf100375101000114300030410031330001303dc3cf0c030c510037ff0114040503d304400300c007544c1030004070c100010000070f03343c00014047041040305013040300c7c41010070000c00f33cc031101700030131d3704d0cd31034000fc1304f400c1c0300140010070470c30000000df401c01010100ff3430313c303c07f40c103300040331c0c40fcf3004300010730d3000c400301033000000101c0c4c3304051cc1300c0300407d0c1000001c0fc41f00300c7410d4c0044030f0400401030000d0033d70c07d0710410000c0f07043001f0300310034c300040d00130c04714cd305710d00410c15cc030000c04dc0c000dc00c40300510450d1000004c30c335f030c00507c000000c03300003d301104f040c0c005d03070f0cc04075100003430c4000301400d07000ccc300104100113003003c40c33c0040c103c0cc110cf0000030000001f03314000011000370ff0cc133000030051c03000040cfcd41c4017d300004000c1c3001c0c10031100001011f7300710000007f000003400000c10070001334003c0f00f000cc01030001c00134d00c000134c00000000000f10450f150400100040cf4c00343c00f030c4f0173001010001113010033037ccf40dfcc4d30c304140004000400cfcc01313030033101133cf4340330101404030f001334c53033300d0010c313d0000c0005ddc1cfc00044400404c00030417c74051f3d70030dff3000110130001300c0010c014000d000c503c1050005033df0c00043100034103005c03013003043734103130c40573033000004dd0010041;
rom_uints[650] = 8192'hc0004100f370cc0035c1cc0c5f01300570330000040011100c0c05000c0c1400c3fc133c0f430053c01f013300ccc4404f11003f003344010000103010134010400cf00fc0c030c30000f570140047c3043143c570cc03d0c00f3301cc3c3f3107477000130f04010071c7000045d1300000cc0dcd005c010014c3074340310c140033c004c010cc00400334033031011440030000103140c5100303000f074400004d30503034340430713047300ff4000c13f10000004104300010110c0c30054c000773003301034000c0d4000f000c0303c000c4cc100cd4300500311000f4330004f0d100000cc400150000c333011d0cc00c00000030130cccd000000c1004000cf0c0c1c00031c3c0745100300443000300010001010c00040001730103303000d3cfcd03031c00030f030cf30c000d0003c0410c0f010000c7f03c004f0107000031c0100013304c31c003150013000c33074040cf0330050c00413c001cc100cc0c03010c00000004c04437000400f007c0c00000fc13300311c1053344030f010c51403c41030041c040770400004003000000ff1371104010000001d0c004f3000010004003fcf3f00403000774353c000cc0c005d30c573740013003030c0100005f300073003f000134071000030f015f030044c740000f00033c00c415c010f370f340741300005040301340030304d050143100000c330100300430f30440453000540fc34c3c4040000443010f0c34001c0003500010075000cc43450cff00d1001340c0cc00400071fff31c0c0f50cc33303c1300300073400544005c01000034373c030c0001c0100031307c50d300301ff03c40130fc10017cc0cc4c1c0d00f0053005003300d1ccc470cc040c70031c0440c00f3c4401041371c4c330711c171fc07c50033c0173f140c07c1300700410000400c0c101c0300df3330cc010ccf3f33340c010303100c0000040c4040001fc5df100d1c3310150c0000131c1c00003c0003d5c3000073004500013c054044400cf0340d43000c400003000300370fc5c070004003c0c3154331d3001030037c5350dc0c0310c100303f40033041447410300303cccc4c013100010103cc043c177000c01c400040c00303000df4d4fdf004d44101040cc0cf470000043403040403f4f310300d11d04ccf00c0f4cf300404300010030cd1c400000d00070c030040d04400704100000300130331345000c0000003ccf303c1f4370041c100f3c0000010400114034000cc1004003c000344fd03c030001050310307c30fc043700101011000c0000003fcc430300311030c00100043744100004c3c303c0000074104d000f5033f4cccd3370003507003070301df10070300dd050034000100c10030010404001c4f0c0f1c0305130000ccf3d33d34441c0c00d3511300000000403151;
rom_uints[651] = 8192'h4030c000c00c0344c0d30f0d4300000c370c433c4ccc0404cfc4c00043fd050400000000400000700c500c00310050c03fc14003f410c431000c3440c0004c05400003c4c0f3101340000f1f040c50c0003cdc414d0000404404000100ccc400ffd3c7d0c4100034503cfd003300c41d0030043000d414c00030f30dc10540105400531c0d0000c000100000c300c4001343004000c00cc547043000c0d0d000100dc04014410ccc04cc001404cc0cc30c0ddc0c0034004c30070001fd1c00c0cc44c0100c0cc7c3000003c00c3010c0000004003c1040c3000400cd300c045c004c000040400031003000f1100f5040cf473034300f04044010003d4043000033c4430c403d0000014d0ccccc1c0c00c0700000400f00c0c004000400c0c030400c3c0004dc034030c51c343f404d307f0104d4d0310100004070c0040c3dccf00cc0c04f1cc3404c000130c44440fc1440104010003007740cf0d4f0307c10c0ccd01010031c40ccd50311c014c00dc040c00070300404000c5cc300000c001c0314340cc004530cc5c40000001fcf3100304c0cc040c00c15c110cc10c04010c4c4c00c4430f40070101c000d1c050cc3400f3c0cc10040cc500c0dc303dc3c43c400004000100ccc4c007f3c0730c0104c40fcc0070430303400d00c340000c0700d300c0c400c4c3c140cd7007c40404ccdc3443310d00044c030c00570fc1cf003345010030c405cc030330c4ccc30cc5c4743040047c43f00c010d5504ccc130c30c0000c0cc11d00c00000000cdfc3030700c4130f10c001000c030cc0100000003c00000f0f4034041443f50c400f700c0f3040ff01000c0340100013c01304530c404030400401cd00500140f041fdc04d0010dc000300d300040c00cf001cc0cc00c04404f31c0000110ccdcc1d431cc0d3400c0000030000c0c0c04310343000000d300d004cfc003c7400c014c000513340c00034330470140010030404cc00130330cfc0c4407cc4004034cc0303047000345c341401cc30400300004c000c400400ccc0c303ccf4cccccc00dc00073000c40ccf50404403cc0500c440543444dc0c0000c00403000000c04030100044c010445430c10000dc110d0c13cc0d031c70cf00cc1c40000004703ccc4cc030c05f0c0c4000df1000000d0c000000000030ff00c0c4300007c00010f047110300f3cc440000013000554010c03100003000f0000030c0c710cc001c0c03374c71df000000000c3300d00040c0c3004c10533003cccfc004013033c050d0c1cdc00404710000300440434c1c300003d405c400c04c005000140030010c10400c000f130f004000040050004f3c0c3cc400001cc44c004d400cc370d040000740c0f0c04cc07cc000010c30040000430777c00417c000c00000431c030030cc51104100cc10010ccc00;
rom_uints[652] = 8192'h10700000101000000001030cc0303c0d103050003c00171003c0030043c73c00040cc0c00c00001c3030001033374003c404103c0300003cc0000030c040041010001100100110000000010cd3047cc010300cfc0c040341c7313dd40330c0d31f00f0130c3004301100100f4cd05f00401300003c310cfc10100f0033d14343131101001100040f0000001d1030313310c0100000c473133c5303030040300100043c0f003c71f00c33f04000f30350000451000030410d0f30143035030001c10000100303d0400c01300000010310000010000000130d10037000504740cc10c00000c010300001710403107050c0cf1031c0c0010130c00010033010301c17cd1f00000cc0543170000075470c3303050333030f403f10c0013030071c01d0100300001c003f000010100440301010010053530c0c00c0f037137c1434000000001d40001c013007007137101100005310700d1001030033fc10007000c100040c01f0dc04004440c31314070d45403007030330001cdf03d30377033d5131071000f37333010f430c03014cd0000300000330001313c017c01000103004dd5d35004010410000010700503d030044344d3c400c131331001030cc3f30440d3c1f4031404001c30c00000300003c11d00034c0c1345500100c1010c033ff3030103d340c7c04040300170f4c005033003040f00305301c0d1100c3000014000037d004000054405d003011c0303410d001311f0004041301d0100c5c500130003500c31cc04c031310030f100c0c343c003003310c0000000c131700c034000115d340030c01c5ff035040100100444000000c00030cc3400c510103717c1400101c53f000c044001330000d040000043d311c4350c314003d400cc1c00d1c307c001000305000c10410014c0cf0fc113000003707f000f05cc0740ccf3c3030403000f0314300001ccd3001c40c000415c03c007050ccc107cc500500d43c1033300000400c041c077350450c0c03d130c00030330d103107000c3d04000500c070043c13c03030101300073c0c443110301030040003404030f1cc3c100400c31041f3300d77000c0c10031c110c00030400003c00005010040c0400003000003c3f0030303ccc00c0000100403c33c03c00fc3f0075f33000c04513413cdc0cc1500d340d30000133341000000404c0f3004c0000cc3000004d101730300411040c000331f07000410c10310c3d0033c000010401f00c000000040001003f01170300c4003500043d0033f0c0031d1c40c3f0033013000c3034170303310c5c000071040c040300013300305f003000c01110c040000c0c0041057c13003c543340345311ff30c103cd0430041000c0040c0000d43301000000f000d403303000000301d00c030d01dc0c003074c04031440c0000300000c334004030;
rom_uints[653] = 8192'hc50000c0c034100cc30030030000f300dc400000c030d4000053f1030030c01003000154403000000010004043030ff5c003000c10040c53000003c01000c40010001dc3c3c0300104000133d103c100030334003dccc00010700003000301000301035031001d010033334030054035107013730110303000d00007130410011d340000000000c000f000400c0000f0cc17030c0000007040030000100d000000f04d000040c130001c3000c40010300300437000130530cf5130dc000000c000004000400003f3003300401414403100c140f041000004010000000001003000030340001d00030c00000f0c3000cc3cd340300005004010000113c100100f000340030030c1000000c03037000000c17040cc11400300330c050030c3334011c3c3000071000000c000304100010000300f0cc51cc3000cc0f0003400000011000373004400040c003f4d00d4013001440300434f301000401033034001133001030c1c017313cd5073740000004000c003144011c000003300001c00370070f340011c0011010043cc00f000f0104000d0c00000c140c00f4f1177030c307047c3030310003340100300014730000003007004c0410300005c4c0300313303000101dc1c00310040330070300073500030100000c0030000104337c0030c30c00011c4150003100330c040dc00f333c000001003000cf3000000cd000000000070d010f0100300000033003cccd000000340c301f0433030c0c0f4400c00400070c301c3031100c044c0440350d330030031010001c070130cc300000105d00301000000004303030d100cfc4013d00030003000100003c430300c000700001130f3cc00c3d0d04040400c000040d11340d3001c0c4030c0f00333030000003130101d0c00331133d1c405000010c3400d0c1003c030414000c0d01c0f000dc104004003000035400003334130034173000003f0000140107c04014300071003300d00000000400300000000c0100100d34033001c0c3303304101c0d0d30c0030403cf0005011c31d3000000003c000370f4303c00033000f33011c410115404040443331341f50000f00cc0040c51011000c070073004000040031450040c30040c0034000c030000003c3f000014370c0c0cc000000c30300000333030c4333103330d00c40031101707003034007c3c0d0050340f0f30c00114103304040034c0004001c00c00300ff00d0f003000c30c0c1000071d000c30013400300d040404d007003051301430330014003c100050003c00000c0c3c0c07300c05000300003110c000100000000000030001c400044001c001030000001410f0000c0011c70100303303001000340000000d0c00000c1010000c30030c010000f10c010404100c0d303c000407c40dfc000003311c0f340401d01400f53000010;
rom_uints[654] = 8192'h1050000f105c00004130c0300c3000f040cd50707447100000f0070030c437000013307f3130000ccc3100303000f04040c440107033c10310430440c000d030000f3504701c4410f000f03114c00c33341f000445c034c0c4007ff343c034cc334010410354003cc444435007103c3cc330f054c44700030300c04000c0f0000400033c00f4004c0030000000044cd330f000000004040cc3300100340cc0c003c10000d4c43c04c4300c00d44030f000f400f000300003343400d0c0044000003005c04c00c040717c0c30f41c00034c00c0000cc00cc0f00330340c3c0101000103f04030c000007000ccd35000310007743f003f00103c00100c057000011010300d14770000c000c3440f003044100300c0f0f30f04700c0354031f0d44c0004000413100170053000341c11cc0c0c00000037040003c001303c00c3f000300c00034700cc0030000f0305f0cfc31d13437001010c73001c4070000cc0c0300000cc00f01c0f0c3310c1014f3403011103035f450303074141003f00c700034fc74d41f44f0500c4000f000c03c74007f040000d000f00134c00f1c40044c3004f03fc00cf00000000007551f70500003c0313433fc000cddf010d0047cc1c10030337003c0003c4c001000c000001734c070c00005404000417c3c3771d00010c1f00300c000000c303c700000100007c370300100c40030304400d340030000d0f47304037100c0000c3400f07004cc3c0c1c14030cfc0d0df34c300040100003703000000003f010fc0cf0c013c354004cc01f10c4d33070c00000c000c7c13031f0340030500004703130007300103c003000000fd00cc30c701c04cc00c0303c3440101c00cdf53400cf3cf05031c0003053c04c0030c414400400044314010000307f100034f5d3400035c0ccc3314cf410d4003c34300010c0300014030000043040f0c0f010003334101000f330303403003000c03003fc00f000004033c000cc03300c003c003dc00000001031401f0010400004c40cc0c4f0010004000c4c30001030001c003030300c00c0f410c0c000304034c30034000c5010101c14cc03030f304441300043dd3040f4c0c440c03f300c3400103c40104c000000c340100c005c0000c10004fc400400c000710400c0000074f00000cc40f00c00c01c00104c40440cf4cc04043000301000400050f4d300000330f40440f1004c31103077043005000000305041077350000c0c4cdcc0400000f103c41030003003301d40c130100300341005c0c4c0010000134000700400d003040034040004003407340000403cd0300043004350005c50400c00ccc000010074c400330040fc301401043071500413004c0d00001c000403003000dcc00034303f34c407fc70700cc15370c0c0301070303d000c04f001c5004000f03030c00000;
rom_uints[655] = 8192'h30303000040c33034300fd00c0300310040cd314110130ffc0001c01131000c04c07c5001001cc540004300400cc4c0104c03307c3dc300c15303c0400000f0017f04004000434005040430433101403440010f30f0434c0d7330400d310c33003d010004703c0cc14c103001f03f00000030c00444f00043000c07000700055031014510004003030004304f47c450100000000110c4c5c50f0011d4c0404140010000443d400c7c000001001c0007034000000030f013c4100d0f400005034033c4000c0040c0f10c0000000400043000400000fc1104c340cc4c04cc01cc0001c3110cc00300c0c4c0cc733050340f1f0007000000400c0053c4f004053004000cc04300074dc0c043300000ff0d00cc0d0d41330040300c0cf40033000073000f030001c00fd1c30f0f017c000c00f4c737000c00030040133f0030c140305000143340cf371f00307c0cccc0311100df0cd003101d410330fc0c0c700004c0010013f3c0050f0300c71d4c30000047c031030001c570c0000000770c443343454c40000c0000c30300430f40000400030003c00035d044030310000cf030541574c000403c00007001053c014704d0440c01433440330100d00501055035371003303d310030f00c3c03055c11110c000430ccdc330f4004041f033c0440031fc4004f350310c0cc0300f1c37f0033140ccc000403504000000c1341400c04c044c04004035f004100f0004075401043500f000000137c07713c431f004d400ccdf041014c30c0f300c4000000004c000031ff1d7c00051d304430030030d4440c01110043f0305470000010d30c034000110000400300c010054cc050c31004300000040041c1741c00000cd0030d0cc3004033c04c53100c4004c1443cf100440001000043c101304305503004c703340000c03040c000003c0131cf04cc000134100c00140fc0713d43cfd74c51400003000d0300c104cc10030c3303100000000404c000010000070440c00043d0c30051050303000000130033400003000c400c41054c0030f1c140d3fc34740dc130400304300c33c001300113030c01c73c1401040c03031050c0044100c000c05c04700000003401c00d05cc000005440f0000c03100c0004c00c0313000f074000003c1031cf357cc0c10c0d4401150f5440d0d00003d400030c4c005304133303330c3c0400c4301104c00051dc0330003000173431000030c7040310000130330ccc434004f533007ccf1514cc0300c300140cc30700000011400000004104130031f011015431003010000c0034034c3000000001003d505103f4300c00004c00000cd0003000010c0057034c01130c0400004c001434c0044175c0c00010004c03d000301153005c400310000704c30700337004c0057004407000401040cc30c0435c4100400000;
rom_uints[656] = 8192'h34000000000d00300100000c7430041c401400300c030c5030001100001c4c40000c7c5d0c0d000030300001103c30040f510c00000000c731400c040cc0f0000c04144f000c300c00003c047d003400c00f0c30ccf50030cc0000cc30304000004101f14140010330c04c00c0311cf30000031c0c100040304373000100033050300c00031431040c0c00000010000f400400000000143c3010104f730c0d0c00040c300c3400d04333003000d4003304310330000034f001400000c700300103010c000010010000007100140c370f000c5101400003040140f04c01f400c01100001003041000700300c70c0c01400040113303370c00000000003000000c0c000c010c1310300137c310f037330c0404071414070340310000140f0c00c4000c1000110c00000f0c0004310cc0333000001103040c0030c0c3514f04000355f40c0c07011000470c00003f0300000d0c0c1c0400007c01010c0d5005000031517300470003000c011004413003370000434dc0c0000000110d4140443430f700500041d0040000034c0c300000031530401c00007000030d0c3003001100304f73001c0000400040000300cdfc00010000f50340015000003004001031f4c0000d30000100f1c03cdc00c4033031043c0f05300c000300330010cc050c0110000c040300f00405c431c4003100c104c454310c17000cc00040d00d040001340c1000500c5503003037c00c0f03303c000c001c003030cf140035c0010330c0d0c400001300430003f0300000400c303c370130414010040041c1c7005c0107000c0c040013000003314030cc074030030fc300700710330430033c050000030c00000000403004004f0400100000c30004030000003004013300401f00030037c1003000f007004c400307143dd41c0c1001c4040fc0000d1d00003c0041440040431c0001010404404730310c304c044c1010000130c170041040043100c300c00001000040010000000001000300004130103304c10cf30100303000003f00000430000000301c040c00400400c330c30c300000303cc00000750c0034013000030340100cc01010300340103c401101c00c010131070040073c04000410c3000c041c334003003ccc054004033c00c4d0304c0000073d014f000f00004440c0413004340000005d00f000cc0c404f10c70300030070040010300054100400003030cc0c40100710000c40700c0000103c1033c70c3040003c0733c3c0f30000403000334340c0003730000000f1007d0d400003447100040033100cc07004f0d0400050040c040040010300410003c03dff000d3300c00500041c104c00040f4000044cc1330c700d030000104001003000000000c010001000403cc0310000003350001300500c3001350d3534003030000c30030311114041003000;
rom_uints[657] = 8192'hf0f0000411050347300033f0c00f4117c030300c0051010d0c4c1c00f000003000d4cc040303373c31c03004c000103150071c40370c00f0040031c1dd00c100f001f310304003d70000100cc100d003004cc051f1fc030f03fd0430400004000300303300070d0fdcc0110c304c5101c0c70f4c031c0550000d0040c0000000cc40c7100501000000f0c0130001434100071033000df001003100c04dc70303c0014f0003d70400c3c033000cc10131034c0c0100404c00c00310d01c41c0f14040300cc0003c3d04c444001f05c00f30cf100c30413300f0f0001f0d300143001c300013cc0000c5c440f1034cd00f704fc503333000c00cc0000701c100f07d00700c000d03c3014d0c53040c0000fcc70c01540040004304d300c341f00300d3c10017c07175c301c3c3330c001f00003030cf00c100cc30f1001cc01000010043c4304541000d0004340cd1c14013c4c40304050010c170301100c40c0300fc40700f34cf0f030504d0c30c13140c107c1000c040030050cf00400c130c0013c1c034c4cc04cd5130304f4333c41c00f0f13001130d00110d3f51011100314c0010c300100030033d033041010130101474000c13001454cf70c1dc074f10330003f40400c10140140003300f34055d01d0005c30c304c3030c5104fcc440003dcfcf100040c00034cc40cd003007ffc0d5070d40cc0c040c00c3001001304030010d0c703fd00dc0003001310c0f4400453c00c1c0f0c1d0000d015c1400f0f310cfc303c000c00dcfcc430f3030ccf0030cc4030007fc03f14cc004f041001400003f004004fc3dc034c403000033c50d3003300100700304033400d301110430cd0000dc4130030730001401cf5c141040cc3f04c00003c40004d1301073c03c313c0040000330013370cd000c0304ccc00000cc00340c03f10df0000dc0330040031101c1001cd4000433030c44413040c3f000030030440d0133c01f307dc330003d430f00013000101c140000d533043c0d00700300cc0300010dc0000004f014c00400fc0177f700334335003c53f740000031440fc04dcf3c30100d410310c01001c00400000ccdc00440400040c30d5c3400c10c1d1000053305df0004f0100003013400400310c04300d034300030d0045000000d04001f00cf04c54cc0c334000040440d4c3371000fc070303c0100310307f01041c00700400000fc000c00d033001011c3014401c707400310030544c04340c30c1d0040040f04103000cff010c1013d000030001c33000cf037cdc3c3031005043c0071031c0d00c03005dc04013010fffc000100dc0c0cfd0040c3000c0000d1001cc300033fc7c5c0030c30000300c0c3000300c300c0300f00130040050300144044c30c00400434cc3c003004000cdcfc0070300441030cc0c00074330c07030d00;
rom_uints[658] = 8192'h104040c7f700d30d0434013d030c031400c00c0c510f01000f37343c43154400041444cc00300d00dc0100f0f3311c0407dd4fc0d4cccd37c0101035cc00304c0111337440000300c0053f05400010c000400003034730115c0101300f3f04cc1000fc00005400000031300c00004d0310044c4f030474400cf3d030c50000414d17411f03d000d0110c0cc004cc430314c00010000d01c3c130010070443c000c000010055d00c3450ffc0d0f000430010c1130000c1c40034004511c10c0c0f34c0404004400030fc0013350ddcd4000513400000d3d513001344c0dfd0c00410031044c040d100c400d1c000451c01030000000700d35100c00c000000c0c000007c10c00100140014c05cd4413fccf1ccc344010400dc450135c107d00000107d0001c400000400c004303400cc1c0747000400c000000300301040400010c03d4cc050c000043cc35447014101310300ccc0030000c1f103f40010004c0033f1f07540f040040170430c1004d400000003d00503d00075d7c004014140fdc5044c034c3000c0030310c03cc000cd0047c40000401c500400040cc0f041d0f00500c0f0c03c0304300c403c70c040000c1d0441103341405503c04c7443c13041c040c400400f03c00cc0c0c7404f0500c1137534c000cdc0c0003310000005fcfc0034cd0340340711000540101000300717c00f01c01dd0004d100407f000c05c310030f0041003ccd43f3350074301110570c400c7015c4d00c0d531033cff0003300435cc04d0404f0031105345c00430037400c100700c1050010f40117310c00535c00100cc410004010305d10310d041030cd0ccc3ccf00041001140000c5dc0010140510000c04c0317fdf0000370d10000dc04fd000710c0001173010100300000014053c07700504010d170301000334000434140d0c0c4c00100034000f0f1f0dcd0f101004003c00300030000c10310c0c0fc000701401000001c0300000c0343c3300300041075c00340c00fc300057cc43c0000f3c3c03100f30103c0c04d114003c0043000c130c00034d37000cc1004f3c0fd0040004c100f10c13c3030344005101470000cc5044700f400000f0cd3c0001001000f30d13041040d430043431000c10c0010047035374403044301ffc044700001cdc03fcc5010004001003034030cf510000734331305dcd30000f030310ff00c01cf0000c000cc40010010c00041007f0001403504403f13f0dc700010010040013400000c030ccfc07dd0000f41c301d00304307c440c300074000f00c10c041347c0c0441303300143f4134441c03c030010d0d01cc030cc004c3c000034f500000303710c0577c0c30c0c400cd113d0d040000cc4300130c043174fff400014410c07100301401340c10100304731300c00c73400f1f140001334300c01c004;
rom_uints[659] = 8192'hc4401040031334f000710f311d04473073110001dc40c10000074300c0f4cc0000103c44074000000fc5c00340050cc0434440030450dc047403440c05003001433c1110c0140010370003c13c400c10007143fd300403c3150044c3c344774f4c4034403010c004ccc074000033010c1331037000c031dc033401104171c00c0115010330100010003c00000150c0f0050f00010003c531ccc10103cc70c1100000c500c011014c041c043003007334000311000014c0c10000500c174404c3350400c0010144c3030d0030031d1c030400001c05c005100003003507c3035d0453440c4cc70c0000330cc5f0500c00c00c000340000030330404503000000004c4c110400001f0c0c0c75400400c4c04c5c0c0445703cc00070c40f3c04f0000004c003c4d14013430d00033404104000000c440000004c13c30c440100000433010c000c0430014d14413000f4cc0c47c10130f1c0303430001004c314014400004c47074400300010c1f43030030c43c570033f40dd04340340011d741c010f00f435003570073003001d30033011004fc3103000300401110c01003141000073041d00c3304304140c0f0570c1400031c10cd0050c0143cd3010c01cc0c15cccc04f1011000404553307300f0101700317030410150c004040340c103400004c33f030c040015cc313001c40501cc0c0c073501404000d00403f0400130040c003cd000440000c44007c03330d00110101c000c300f3007c04f47300d3dc0044770000000c40000d0004f000000303f000044070c50040410144410070c440000000fc3dc500030f744c40d0040c00d001000003c0004103ccc343151c704331044d41000f33c307d04050010000f140c0300000f40015c4000004000331030cc040010f11104070007f315cd10c045310303c004c00f50c010c0000303f33ccd13400314300014d370370134f50550440500dcc0d01d73070001430d001f003404000003c03300000c000d030100004400c50f074003000710c00cf03140003c10175c004c105cd030cc0075304c0303c53000070030c000000cf03c405300c0004130f0540001140001c4d040013513300344010001ddd00300000d7c003c000dcc1c40130401c10410cd400000c1443c3371000c0340103010d0007003dc1d04d070fc0c4000401041003c0330070000d00f00c4733f144000040401df000101030cc0c3c10314400c00330c5d03140004001c000fdf0030003317104000c1030100330cd00001c5030014d03001cd0c3140000000403f005004003100030c5730030c14c00740000c0c00010044d33530004000c5000000ccc014000c03c47101043d50fc3c307010c0c00c540450300033003303740cf0030100c50100000007010c3040f75004077c03010401053735341cc41001003300000000;
rom_uints[660] = 8192'h3344000017100000100730cc030044c0330000c0010035f3030040000f30441000f030cff040001400c400c0101400dc731300f3c54354154040c0d00fcd04040040f40300340cc00000f3ff400753ccf10c44010c471143400410031cfc0cc0055375310530001033cd7013050033000043030f01010400000307c4c310004304c43000000000413003c03070007407330c0c00000100c3dd07040307f4cc3430004c05c41017003cc045013ccc0f7403c030d00000540c114000001543133040c733c3c0503431043300347105cfcf0331007440f303340014000c701c00003c0300000010c70003000c1c0c00310fc00c4f0fc3140c0001044007111040c0001c07cfcc1535fc001003cc134f0703d30c115005404330d1430000f011ff1500c00c00444400d4000310733003000c33c0340f000410401317c0c0440d00c1700c0000cddc010010147101574d0043f03d030141c0f0400000300d0c00c30700700051fd000c7f000f40cc3141100000c704d1473c500010ff3c0c4044040430c03001c00011010c404014c40030c4150033c500000c0310041000000041070fc00d0fc0cd0c4700070c0c00c1030000103117337c3c1345003303c001440fc14440cd3040005000034c00c1c13cc04303010c430f733000d004003ccc0c130033c10ccc30d140c100434700cc4333d5d0003000140300f00100c101444c00040cf1030400400000c70f4003c0d3030400cc00f71073000000374354c30f401105051010041ccdcc43dc00003c01c403430c0103037440013000100f00f30005040c010f00310071c3330700300140730004c300141100000f0030f100573300710ccc13c103f14303370500700c003fd40c00004004071c74f0cc3033d0001c543c000300d00fc0145500c3533cf5cc0c0303c00ccf3040c0000c140330003c43000004dc710100030703750101f303373f03000d0000c00313dd30700004f00013004000c00370304003400330040001001c07330030d1010f13103053003700030f4c030034c1000f00044d44c043c03734c3030400c3f0c000000301030100130d3504c530c000c1df0701f3c337000504ccc1c01000030c70033c03043cff0014000f040d4013cc0001100c0401c0303030c3040001110d00000001c000dd00c1c1044304103040544300f00100740f3305511cd01cc00700440300001cf034cd01000000340f000c740c4330010371c3010300c0d34c00c040c0030010c0353c03000f4445001313070010c31033000d00c034400030c04c34000000750c0d0030c00cf14040f140333003f00003dc100000d0c000c00c001003310147103700cc4437c1c30ffc0f00f0030f00c045300000113c00004c00000d00301000c010434700034050070c007000004dc1c05100030130000000010c100153;
rom_uints[661] = 8192'hf0f41304c010000c3000100f3001000fc0f7004504113000000c40303405c003dc7c1fd0310c1000dff403103005d03dc4740c05f530440c0000103f57051c5c04010171000000300000ccc413f3303030d710c47c4534c40c3011500c1c4c0cc07c000c4010c000f000000c430d100dc131f051c04c1cd00004111c7f145000f400070034000300010c343cc0d0011530303c30004cf070001c0c0d500c5d0404c0013104c03101340c7c010110c0004417f1000c030c104000d005d3047f3010c0117f0c007010040fc4303434051c300f4030c04cf50004001000f0104400c400003c70c1c04000401003d004000013d3f10c13700000c0340c0430304cc01010030740f0c07cd51cc000000000c445310405044d10044510d0c04d134c704100700cf500500104414470300c040400000c4c1400100150ccc0040d70010f4c10c0d14c00f00540c00c041d3000d4057001c50d370f0d30c030000d3c4003100110c05c043005007030314300400104f0033f04f0dd404cd330c105054c04f441f0c0df4033304dd000c510147f50300d1000000c31440c70c150143cc00cd5c00c403031034000d0f433f0540c000f13171f0f711c10441cf0c403c01c3300fc003040f0cf0c1050304cf00f4c44c311043030d3f4000030c00c44003030c3d030c0f413000740f0cc040fc30c7430043c3001c0c00170010c003c137030440430c0004300431c00f7cc430010003c1c440ccc34007c00cc7fd0d00c430034f1305c054730300dcd4c1c00030c03000300c3407dc5c074c0f130000cd0400c430c40c001f0dc70000473c5750cd040c5040010403047005c011014000c5030c01401d10c00f0000100403dc400d0c3033100700000000405000100003fc300c000c04cc0c1440cdc040c0c0001c340000cc335000c000cdc100c307cc44734f1c0300f07cd74354110307fd43f30001f41311401510104043c0c44301400c00c0430000cc0005cc1cc1000d0430c00414cc04044f35d54c530f007dc00000000430c400000c0c030400400303050040104dc310c30c31c35730c00001c14305c10f4c100c310c0c0040001004f7403000401000f1040010c0004d304044c0c000703d070300150c4000404d54004000344503030000035530500c50430041d404f054c070040c10fcc0410cc500005404c100c3003500c30c00004c1703103c5d00440300c300010c31f110c0074400030c0cc0f30034d0000330070d4dfcd05f030c00f0005f30c00140404c0010dc010c1c000000d303c000001011c45c3033300310c073000ccc01011c041000530430c401710300c0350070400c13c00134fccc50c1040c3007fcc330c0cc13c0140000c0401405cd0017c00c04010030c440cfc0cc3c0c130d00000d0c000103cc0504405304cc710c1f431c0003;
rom_uints[662] = 8192'h30105000c00f0400cc0c00434d130030d4003030d3013cf107001004f470333030cc35005cd334401c3404033334110003cc00c44010c05dc00041103101030104515c150cd100fc4000500744004c0c1044f0303110cc41dcc15f100005c000100017303500c33000c01d000cc4f10f400c11f01013f14400010c0c00001300305dc000c0c030530005cd004400d7c70c10000300304300f001030100f73000501004f0f01c0cc0041c04f000c033d40c455dd300000c3300104070101d0c11c40000010030c014f03430f0ff0c01550000f530f001703c0030000100f70130f0c3003cc0c00470000c007400f1300030300141f530000003000000073c0400770c0000110c0034001f031d4f0740c001fc4047031c350c3c04700034d030f7c4c0000040f400fc0c340c01340070000403107000004000000003c0f31d000c0c07045013f3c10040f4f5df17f0c000003735c0071dcd0c4c00cc3d0c5d011040f5f0000dc1f401030c0000f004001f0000d00f300300c14c303f0c30001011133401c4015c50404030c1cc1000c0df30000007000043400f31d1d404740003313100010c3000d4c00003044cf404101c003c0c074d110014004d1404103343000070001c0c003c07f0c0307c00000cf43c14c00cc40441c0301d04c1f31cf000400c40d0004403c313f340c1f000405c00f0cc001c1044f455110ff03f4c01f40c0c4c1c10dc10700d314001f0d0d3c0cc3003f0301c300100031d3444cc0c0f101c5030cf4011000030304044400130fc0c0051101300500010700410f4141c03011000005cf413f300111400d0c00c40030c041ccd00500500f40c00c00030c000010410f1fc0030343330f01030c0d04010f053cf700d0cc44cf10c01070d170043100030d103cf0f34f1040c10c1413c3031c000c7003ccd01d055c01f0000055d04cc1033000c00cc433057f400f0010c140733c0cccc51fc0d500401f0054000c0000000c500000400fc04300404cc10c14500cccc70f4040033d310fc00005170fc3c144c30410300300c0030c335f54004c53055c00d003c017010f344300033c03c007700300131f40071c50c0000f44100f43050300071000c000000001c77cd0013330311c33030100000c00547c00141f013f01cc00000040130fc00505140403f0cfc0c00c43103303701f4073fff010dc1fc01001070013330030c3000f100c3c4530030500003c11330c40c50cc1f005d00000000c00401400c0100000040000310305c1000c011f4f030f0011403f0105d3c00c0f010041700041351f0dc30140030400031003d0001033030000f0c00001c000c53c0f04057f40340dff4dd0040300c3c3c00c0c130cf010401040303d7400300cc04110c300000c7100015007301700050f030c7300003f3000d0cdf301000c0000000;
rom_uints[663] = 8192'hcf000d40330030000c0c0ccd0c044010033400c410100015c031c0001010cd50c4010303c4070d000c0000fc0c3034c4cc0304030137050330f4000000c10f001404040400300034000c3c44300f00000f04413331dc070013f00c30fc0147030003041c00303c0045130100140c17000d3001013004c4040104c03507d3430c0c030341330000c40010014ccf0000000303f40005010d100c311400300f00350030170c000404000030050041340000013c05043c0000df010400000d40070004c000d0330c0003c407030000070400d0003fc00c040004350003070301000037000000c0017400c135043c0dcf1fcf0700000c3000cf0104007110c500003c000f010311300c000003003500000cc3331305413dc4c000770c04443500000f0c0c04000c4300303c13000f030c45d003000c00010330c3000dc504041034c000cc0000041c00100c0c000044000001043cd037c4c44104030004034010031f3c410044073c004434d000f0710400c3c00c0cf34c75000c0070c01f01040c0cc5010c0430000003c435d40400140000010d040437000004013001c50f30000044cd11000c100004c70100004100f0c53d000d1c0031000000040003000500434c00001700030047000107cc33c3403c0c1d43003430c007333000000c04030c017034001c530000410015700041d430340f0c3104300004c0010004040cc505000c113000100033000c130401400f0d0c000f040c0c0c05ccdc0f34f030174c00f04000c4044010000c03cf00000c00d701c00c1c0c07340cd443c03413040003000003c4033300435c300c3cd303103007040c3d0f030c403000c331143040070100030f14004c00051730303c041c40c003430031000003010c30c37d03440400101dddc000c014313f7f300c00300c00351003040077031700cd0c34100f050c04301300ff000ccf00370300ff05000504f7f0303100cf00031f00f0000000cc400c000404044031030501c07110130c03000100c5300710c4cc000c0304c3040c0030000c10500000100c4f1fc7030000c330f104c44107000004300c03033c0f0300043000400300033100001c0f0504303004040710033030140c1c00170cc000047c070004000304030f1c0c0031007c300c0c0004030301041300030c33100f04030417040301440700040301001f0004cc00d0400717000c044344330030000314000030c1000c0c370fc00c00130f4c0004300700030300f741000430003100c033c010c070470c047d003cc00c0fdc0f03c0400434cc0400001c3f0101040107fc010c3300004c0305000030034010300000100d4c001005fc0c3c0c070403003c000507374704044000000340c01d0d00030d001c07010030110c350004311f0701303df310010c0d000c74000cd003147c00000c;
rom_uints[664] = 8192'hd40400400044cc031000344000d0307cf00c41d0004030c0000d0d004400500000500c1000cd000040cc00040ccc4c0040c3044f0000dd104c313043dc40030304400400437c0471f0000cf00000401107040030140040c1040c007300034c0400000700cc40c1c100357103440f0004f475c0f00000030c00dc304c10ff043050f134fc3c11000000034000f0000110014c0000000c35107004cd003004303074003000001c3330c014cc1700c03c030003001000c31c443c001040cd411000ccc00c01d431000c1044cc74010c0003c3300d0030403043037c40c000c000fc00010430000f70000400c03c307030fc11310c470f00005c0c1c103f0000000c07000000500c4c17041030300c000c7300010f307c70c43c0001c4f10104c0df1c0540003d3001d44334040433005000000010c4041f03000f03f0c10443003054c0cf0373f13030070d041c03004730c00430703005007f0fc00304c14007310304311dcdfc3f007007c40300304f0050c00c0c1c15141000004734d00c30073100d53f03730040f4f033317040003310003030000000f00400d74cf3430c00ccc03f04f30300dc00cc00f003c030f004007c00344144005dc130004ff030d30000d140010004141000c0c00400c07cc0773003d3c0370443430f104d0c7fd10003000f00001f04400010c00000d004d103014f4001c00f4070000c0000440503430d7c40c14070d113073014000f000c4c40cc030040d0004d0d1133003740330cdf00ccc4cc000330300c03300000c034c00010f3c0c0501343c1d3003110d000404f0400c3304c00c0ccc7f1c00c04c03c000c40100c301303340dc30400c03dc4004c0d14c04ff3000c00004010ff0041003000400700013c400c010013403300c000000307cccc534c40f0c00ccdcf4030430c001530001500511cf133d03074c113400c31303041c1c0c301cd1d4fd0c044fd30010c00cc7cc400c75040c000000300c0003f01c0030003c00f0404407c0c471d0044040000c0001010c0000040c0030010000c043f40000d10344015f0c0010c00303433c40c0cc4c4cc431430110c01f104003cd0044c300100400c034010c10400000000c40100c0f00d0054001c0c0701c04040007007003c017c11011c0c043d504c004c33003f007300103000400ccf3000133c340c000343000fd0c00cc04040f30d100010303c1044041043004dd00300700d400c4043344040c03074500011300000401c000403c100c7001104cc3cc4d3ccc30c4000c33004304c0300d4c3417f300c0403cd70004c11c0503c0404c3c050704c0010100f33c0004f430c30000030f0000014103070400f34110000c00cc00000f300000d00000030f003c4c400044304004c3013003000301000000000401c0300f100004c000103330f0c40f3cf70d000;
rom_uints[665] = 8192'h111c0000300cc401005335033c004f3c1f33003341d4130000001f03103403000001c410400f01000d30100c0330013033430f1c3053035173f01c0c07010fc3011100043c04c30c000001c1c400110100c0153cc0040c41000c0c03004004003103c50ccc01c00400001f030d40d74050730075011100c400003100005410114010c70010700c0000cd0014c4033000030c00030000413f3004733003770c03100003010051003d005100c04c07400301c0f03c00333100c103c14134c440073dff0000030000034137004430050d100010c311010757f1cd4c030cfd3103501f4003004c1010130000000401050131d53f0d30103000d00400010c33000100030c43030f4170030f31303340300010507743400c0110001c04033c0434017c13c050003d310100701400d030000100310c000310000c4047134000401000001dd030c00d13130140300031d001004014510400013f000f4031df003141000c0504430113033007000fc3d10f0030401040430c0700cf000010c3cf04f405c05130313fd144010000341c007000030330000031100004000cdf00d4f10d00000435300f070004cc100d4c00100f0740f003311571c001334d340030000300000f710430304000000cd00c10400003003fd31d7337030311007fc0000303010007d0fc5d0cf51000d03d3300003007131d0d440d304403000cc00000d1003c5fc30c40c30437c00c30174011cf14c0030114f037000d101c5370333fc003443045000001771000401000c3501300350d10101131044f000400ddfc035000440c034073000c074004f00007d40437140c05c0031015101d0003d001003030d110003c4c03140cc00d10011040073c400034071d104c010050300d07c1cc1d0c1f04f103000cf000d347071c01d7010d0c1301403031c004430d1c040003110411454c31313c010000000cc0100dc0f0403337030c0031c07f034047141001000055071000c00013000f0003c300030301033f530007004714ff307313c131435007000c31474f301010345044013400c0403c010713d4303040300300400011033c0c3000010f3003053330100430051015f30cc4c3f10c31405c3030c3377d0c1f000001350017c14004d43300f0404401000000434110c1303c0f703f105c0030cf10000d00c003000000003300041000c4cc30005003d4407d340c4037030d34003c47310f033f0001300005000f1011404001004f1d41d110001c000304f500d0303000001334030400001300011d01c10f31cc401301031c0c0013000000037101c50c00103300010000f00cd0d0004c0d0010000010400010001001fc73300100300c14130cc000f713003300155403cf340400011c0010710c03cfcf03000c1c1374030c0fc0c45543000cf50175000034533041003c00003d3c000040;
rom_uints[666] = 8192'h71140700c074004501000011c0003400d470004c3005cfcc000400c0103410000110cf0303030003c110501c0100113134d00c0f7013c37d040c00c0310cf0001700df43445300430000c043050001700071d07004003cd3f00cc5f14c34d00000f740040d00003c03031c0000c00030103c10c0c0104100500c414cc3050c00d31c4cc000c00000c04000cc0000001f0f7000100030300d054100101000cfc0100f0370404000400000007cc0c3001f0000df0000007fcc1cfc1005fc300000001007344000cf03050030c00304004c00c0cc7000010010501c1011d0cc4001101000300c0000000000c371c304c0f54400c430005f044100410434000000c400010110013c3100300dd0c330004073ccf30431030004c045c130c330d300000cc074000004407030007c00001f170004c040d33c010400c0010f00c400c03410000d05004411c0cc0c35d74130000000053304370f0004400043cd104cd00cf44cc3000000d4c0c0c01c41040f10f010310040cc0040300005d04010104400f500303100034cc0d0151000cd00dcd01c00003340dc41cc4c1003c00101c004f303c51c3334004500304c04404fd0f000031071030013107704c0c003c5d0500475c40c000c507143040540c104003c015000c0300001c001c03340d0c00034c000330003dc40d30c400f0d001341d033407d10f110f040100100300f0f1040331000f000c007000003d05dcfdc1330130413000c30100041cf30f01c1403c440037341013c3d0010c0cc304103f14c340c0f0000000000c04c4471540035c000c3c4040000fc1000f100130303034dc0007d0005047c0075400cc44c030000543701f011000000314054330410040cf01c01c414000c00c070c700c3c4000011440c400000501c10000001c010c1310000d00001c003df1040d000cc000c00000043400040c0331c3103300cf100011c0441400cf0d3c030c000411031c4c007005d700000070010000c1c130c0d40d03473cc33307c405c3000c001300f40df00c0307cfcd004004c400445d333c7150303c00014000015d300c0f000c00040004c4130440c340104dcf4c0300000001100c0030c1350030000d301c0033000fc30c0005cc0340335400004c143c0044d0003cc04003000f40c00c034c10cc045741100004100000401000c3dc0c00c030001404030dc10304000dcc4f000054100330000004c030004c00045c000f4037c4030500c7104c00c4001fc3134f7407f0f1010c031f330c4131c01c530030c7cd307f000010c0c00c4300000c0134014004c00041c001010041c003001404f41403104c000340403000000cc010141dd3040d010030000f30004c01c000c4c000004d40cd3d01c000c0007d0c44c0040114100d010404c010010011030cc30000040c30cd43300c01004c03f40;
rom_uints[667] = 8192'h3c1000054cd00007d00f0303301047c000d0c0040f0130f40c4c03001dc0dc40004030040500c0000000c0c000000c0040c430fc705c3c05140000004cc0c0000c3cccf4f000303fc3003170cc00530044011c0c3031303d403030c0307c5003041f404007c3cc003c3cccc70f00000ccc010500400ff0c01003f7f030040050c0f43c00001014d3003c00cc4c00c70f0c0000000004cf007cd40c44c0410000103c057001f0007303007344f1f0d44000d0d04c000000ccc70410c1314010340cdcc00c000f41114310004000c01c040413f50334c513c10c3f401130c00030c40700c30000f40c030100d5ccc01004004014313401000040105c04100000000c3033c701030345c000000001010400001c004000005d00030c0cddcc10107430dc3300104c00030d74c00001100cf04c03001cc0c40000c303310003f00cc03100005cc004700c000c403d4370310c104c3410430cc01f500cf030401500700c310c4f30c01130011500d57300cc010c000440400c70301c130050110050c0555033403301101cc0010030c100c003f30cfc400000000404000130031cc4003cc743004070000000c0cc0f0137d10300c14fccc301003345c0004001300050044c10c0c0003000340c5c011140c0c44c0100d010c00145000033005fc3031010c040f0c00c10c0f333d11fc0d000101cd1cf1c54c000103cf0f0003040001334c0c0c0041c5404c0cd50c03403300c30330000c0404130031c5c41001cfc11300c1000c43004f1c040fc010100c034c0f0000044000c101070c0f401010c3010dc10f300f04f1011100c3510c031001c0c03347010f0000130037c0f001cf0000f0003d0c710fc3330735d0c0000f70cc0500300303c30c10ffc001370000cc1701040110040d3003033cdfc00c0040d05c5c31000010c0c00d30030c4f31310c04c50130c0340305400304000cd040000300000000c000440d0731c000000334c1000000003c000400010400c10370c00441010f000304310d700004300040c00700504040c403034030f4f110c015cf134c00cc3001033d0dc03cf01f100737030cccc5400010c000314c400430d34050dc00114000c003c100cc030400c153c005c3c0c001300000c000c3010000010054c01170070d04014c00410f0c010f30000044f30030030d70004c53fcc00140fc0004c30311d400c300c5d04c0c3c00cd0040c00f040004000000000c1400ccf04540f014001cc0000000c411103c4c00071000c1330c010d0d353400100f00fcc4c440010043403100cc403c040dc1014000000c3c01c4030c4fc40d00034c4c300000700003011000cd303500f031c07c0041c37c00c15d774c7031004047300101c3010c000004050000f00f4f004305f07f0f440cf70c15001d70c10001030c01cd0314700503011c0c300;
rom_uints[668] = 8192'h40104340c0f410101003c0005c004c540c003104c303c40000dd0c004c30c33000303c5c04c04000c44400000040c30d0040000303c100c7c31000c03c0400004c0043d4030000c000004440d00000071000003cd0dd0030303c50d300d010d510c4c0f0f0000cc3001054000040f3013400100c3300c0f0d070c13d0430d000cf13300014c00003004000300c0c17c13130000c0000c04c0c3f34400104440c1047dc1dcd5133fc3000c01110c404131c07040100403140c070c330d4d131304004100304000d3c1c10004040300003c050f34000000f14101440740c35005c301c000401f30010001000d700d00d400031d0fc10541c004040003013c0107c1370100040d0005030d000400440000c3034001040c3cc00cdd1303330c1000430101300f011147101c4c0040100d0071c0034f030c70000303000f31107143c741c30fc14074c00c03010c0cd0100cc4f50703fc4400f70c01c7c0c00c0004000703dd0303004f0130030401c3f4014004004044300c0000cd070f0c030c404d050f3403d3000c04413000003104c40c3c000000000f30000000000031c0c0171c31004c31ff3001c0330007f1003f0f73010c004d0040cd40000c04030dc1440003004dc50c00410dc0030041043344d7014c030344cfc0030100cc0cc1340ff000c5040f4100c5100c43c000000530404c0001334004c50f000f301c154f01103403053104003103c0c3430f030440704c50c0c0c70c00d400103007c4031c030f41033070010000c10c04c30310030f414c000d4c4001c5000005400333d40c03f100170c000d0c00000c33040403000f00d00c000c017000000500430cf00001010fdc000f4f3c010040530c4c0c0731c3c01d5ccc000f00300f050000054c10000003030d07d0ccc5430c03030101470010cd0301000f00c3430003cc4144000c4c040fc0d57d343011030d1340c00c0f000d4c010300d30f1f00f3c0c001c10c000003cf100140c0c003070c0001c01303cccf430c4004cc040d034307c000c0cc3041301144410005144040cdc5010140c10010030043f004d401000401030c0d3000015df00004030dd00003103c000700040c410c30ccf0c7410034400f000f43030c40c00110000c00300c070c0d00477c01045110000c31000100c011c001750f0003000c0cd0004103f005c00c1307500004cc00c0001c0f0c010300c74dc10c0c34cd44001cd007000d4c573c47303315041f300000c0003300004377130001f00f00034003040000000f03113301003003410c0cc43cc0c1001441040f050f3404c04c0cdc040d03000fc40f0001c10000000000000cc0f00001553d1d0714c30000074c43330c0c3f4017040030010c74f00c5c033051004c444f0101dc000337ccd3003c00c1033d400c3104050c44f0401c0300000c500;
rom_uints[669] = 8192'h3300000030440477044c0501f3f0700c7fc4000c000040cc0411f01c0c03c3404070c0f0c0030001100f03cc005043cc00f1101ff4434d1000000c3104d3403c3040c4c030400030c000000c400f00003c070000034c34d010140c00c0404cc704f4fcc3c030004cd300cc03c1c3d3410030cfd000034400313c0004c4030c7c04c43004700001430000071f00000f10d4c0030000c1f0d0cc4c0000c301c3f711c330030400fc47c000000c0ccc050004d3d00000cc031034000c001000000041f0c00cc004d05070000000cc034f0000c1d4400c0c03d30c340f0100ccc0404c040007030c0c0c30000fc041734000004c00504cc040000303404c3c00004c014c0010031c04c10300c007100c000f30c07f403334340500c00fd0cd1344f010cc3000cf5003430530004c001053000c30cfc4cc00c00000001ccd403cc0010c404f700cf0cc030c0c400f500740c03f705000cc0f0c71f0334710030cc40f407700015003cf0f31cc0100301300c0c0003d001f0003137fff5ccc00d0cc0410f0c001340004040c334003d0443533c00ccc0000c7010cc17033400030003004d100c00c30047c40cf300100c100c051c0341d3c004c040040d170101374c53070000c00000374374c3cfff03c1000300003dc000f0300000440c0c00c30cc0001cc0cd0041d700c043c1035fc04011c10d5300cc00041d4d4d0ccc311f54443033105c1700c0cc5c334110310003c0004c71fcc00411c00f4313413f5c0140504107300f100100100c01000c03c00c0000f00343333c300700005000cc14fc0c1345c0f4f00001f0c14100340403c104004035f0d040005401c40000550c0c000c01001c0f301300370307000301c11c031404c340000d4570c0c04101340d344f340000003cc450003044010c0f3c3cc7c00300030d04cccc00c4303c043173cd0cc0dc0cf01f100035000001cfcd0f00040cc0c0400c100014fcc0030135010030010043c0c03f00400ccc0cc0041043c50304cc4cd431fc7000c5c0c003000000c40000000053c000440c30003700457cf040400000130cc3c0f1300004310c003304007000003c010c4c0344711cc0000440000700104dc0f1c00400c00d00000c1001f00004300000144000040c0c044104000400340c100c0c4000fc00740d10c41403010ccc04003cd3040c3c10403373101004f3f10c4503f000f030003d0000004001350c407400000030050001100f4003010400cc43c01c317f00300d0000c1f041000044030400c0c15004c0c04000005ccc0740043c00c30c0003004013d00f00c040730cc0043c004c4c104000c001033c350014c04cf3030403ff3f0ddc0c000cc0ff3570404f000c400100f000cc337543cc170403cf0000004033c00f1013340400005c0f30c0043fc4040fcd000015c00c00040003;
rom_uints[670] = 8192'h1014f040c000030d10000000c000301003c0001f70c401100c304000c301100430000140403000007f4c001104000c11001c0ccc00003c4050c070c35c4cc000c10d0501000030300001070c0004003c40001370000c00d0050c0cf00440c0100cc40744700c1000400d0400400d000000000c700007301000133d00010133c5c000c010005000d004300c40c00447c0c00c0c40000010444000100cc05000c1000300400c11cc000000c000c0000000031100000000f3c05f304cd01030c00100303000000040cc0314307c411c5c07c0010000300000040d53003f0fd000cc30300fc0f0300004003003dc4c0cd000003c043000f0004c10101000140004334000703c00070001c00c000cd000400117d004000044037041001010140300cc41040001c4700401000034c0300c0c0f1334001010400c1300f014400ccc10003000530000d050ccc4074c3000c403c4dc00c0004000c370cf04c03c501301040333400040001cc000c0ccc044001001300c003013c4f0cc043030030cc0010f0000700c00c000001040043c000dc0301000c00000050c0c353003c000000c431d703000cf4003000004000000c0f00030000c3d400df011040000f040540c0040001040034c101000c0401010300350c000400010d4733c14104c00000003000c03730d0c104c30045340100014001dc403037500000304cc404040041400c0403001514000cc4004130c1131000000c03040000004c1040c1403c05010f01700c000150c1c00400003031c40004c40fc0004004030340c30041300400c100c0cc400000000400404c01c1430000000d04c0033000c3004030c4404440100c40540004101401c4d03010d034000ff0404005000000010300301004c0004000073f04003103c00c0d0503040000371033104f03400040000003c1000c0f0c04fd3d000040cf01030c0c340c00431433f0c3034f00c000c0d0004c040c00000300030c0c00004100000070c0000100041c0c00c41c0300c34005300c0133cc000c000f007c3c0cc1000cfc01414003740c000403c0c0000143cc0c03034f40c0c0030300d044110001000541401441cf40d003000101004fc00c0f000030c300003c0003000cc100c00140003304d0304000010001110d00007345130c0304000404330003301c0134c0c00007310c00000003fc040000710f377500004100040c000030c00c0040c0c0000d0500cc040c0c000c004f00d04cc0030030c0011c3dc0d00c0000130c0404003c00300100000f07004cc5cf00000004003f0000cc000300c404003c3540000030d000001100100c343100c4c40000c400400044040000dcc107dd1cc403034140433107c00004100000030400cc0000100113000005000000cf0c4351000c400000010100310043340001170c0030000300c03040;
rom_uints[671] = 8192'h303d0000004014107405030134000c00fcc0133307d3cc31c01c07330c13370030f00034f1433100104400403000d04c3c7f34304430007540f30000c403c001f104f1c0000130000000c010f330300030ccf0c303dc03003f30c4f114c40d0c0071400334300000334c7104c01033430330f4d00054f0c00014c71f3740100031010f000410007001c03030cd40303001c1003000c10034c0dd00c0cc1c511c00000103c40471040c040003c100403410003d10000c03c3000300f0f003700400dcf03030004c47c7cc00000c1433f401c1070000dccccd007c00f001d100f0f1030c010330dc00544000c130d00cc0101300c7501000303c30c00003130003d1100040c3c043000cd004405040000c7c13303f00d4d4705404330cf043f0000330340000004310030033010000f003f013107d473330cc0c3d734030c300f03400d7c01001fdc000000cf03430701010f040430000cf134301311004f00c3c1c57df40ccc11f033c000c4330041030000f0c450f0150340113c14010c00540c74dc3c00c000030fdd334c0f03400c170000d10c300040105700031041050c5c000004070000431c0c143033410c01054401f0050c3001044cc0000c030c7340cc30003404040300031303030000c1c003d000f0cc340c00030304440471074c01c1733d3d0c35c4050003dc0030c3d043f4340400101f0011101004004104010013000140d14c070fdfc0c41cf00c14c4347043c3cd031cdcf313cc0010d0304137000f3f3410c0300cdc0f1fc1330403314003030043cc71440403040f303c04d0c00401c01d000030c31c10000101cc041c0c037c0410f4054d71c00740700c0347c3c3103ccc434c0704d0041d00f04c303d0003403c0d4fc40cc340401d0344c70000050fcc0d504104f01000cf0fc5f00301c503300040303000000c0cc0040f400dcff04cdc5403f0500000004f0c35310031c3100cd400001c00013c3130034340000001100017000400000c01040005cc3035451cf1c3000130c00d000d403c13400033140330cc4cc100700c3c01030070040d05c030004c0fdc100c414307003004d030c0033fd730030fc0000c00c0500144c31f10cd11f700cffc400c010737c0004040343001011c140c30c0300f034000c0400000c317000301c000401c0544301c0003471cc0003014033010010c1000f77000004fc3dc0d10c4100004330c4ccc400cc3100c00347c01043043d3400fc77400400cff300c0003c10c100fc3c03dd1cd7410101f001c0141f4c40f30074374000ff300000c403030fd71000c0010001f5470d003103f03010f70053470c0c00004c101c0c3400004370734130f1000c44c7f330003d7410030c0c00c10011c00343400c0075dc010111100c0c13103df000340300300c00c00c503c0c10004000030c10fc;
rom_uints[672] = 8192'hd01c3000500101010073104470c030c0f3c011d00c005000004400dc71cf1044701001050c03003010000400fc0404cfdfd300370c1737cc30000070000043000c0004c330000001c0000401510000300ccf501d1c00033401040044c0004f1d300cc0003c0d104c043d07007c405c0c004dc0300c000004000000400001050c773f4c0c04300040040000170f040100c0430030000000445c41000000c07401f00cfc4103f7c040c5cc0000131f00370300074c00f0c01cc00500c00104d044000c0043cc0057043c300437cf00c3400c10470001504c40700c33cc000d0c30000c0003340004c040cc0c50434004340114c04000000000030000c07c000030405541c004f0700c034f10001c00c01703fcc040c0010c300103030c1c13f00d44c04300c00cc001ccd00341cd00430c500c400f03c00700370013c0130f3040030c0040000c030003000c3030d0030c313c700f004f0c130c0073000fc303040000300cf0f40d040300f4c043503cc000470000747c4c3c00f1771d01c0cd000c00c004c30c0c11030000004000433fcc003003c000c0000047c040040cc0c71104c0070c4c4cc530300c0014105cd3d0131004f3c37335cc5144000000c0c0cc40c0c33c0d00c1014f3300cc0c3711f04703c0034077000030000043040303c000103c03c10c7f037001400cf000733704ff0004c000f300004000d304c010144340040043000000cf000100f073047c03d305dd43100330cc0300143130d00041c000f330000f00cf40cc74101d0000c3cd00d0033f07cc300c4030000f4c0f0370701003010c00000c0740d3050010c3d5015d330f03034f01410040c5cd33c37037107c3401c00075c03f4100401cc00d0c30050f70cc10001c0c433433040003003073003005040043040d30c040cd1cc000001170c00c00001000c00d370103c300c0c00c0c7f40075d30f4c54000451ccdc33c40cc30d00d30c03474c0040000c00000010031000003c3030c3c4053f01350ccc45104df3010030540040044010f0c403403c0430c4d4d3c337000c7300001040073304f0007043c000d44000d10f010100cc0ccc370c030033433c0d070d0f44100034c03440c0134f0c000f110cfd304443104030f5100000c15dc03c333c00ccf03c343f053333100414c040f70004000000d0f050d33004003013000010010304c1400c00d1404400333c00c0301c3010cc0d00300c4330030c3d0030c0cc430030000f00307500ccf30c0c00013c0c0c13030c3504dc31011041c3333d3c0c03fcf1050cf0000f4011d30c0c00fc0f00130400040001300c00055c0410fd30001300000ccc30c00010c0c30c43c437330d3c001014000000f000c01000f110004c14300c04c04c301000034d13045540d51430000cc3330350d4c0c30000330700f00cf000c00;
rom_uints[673] = 8192'hd311110403130000007000100005c10300c01000000c14c00c340000103ff01004c00400c430013c00000cf1c00f440f3c3044c304c40d500004004001000000000374d100c01114000c440140017001c0001c40103c5c0000330c3c00400c5c444300c303c030004300000000404040000340c300fc03f0cd4040330011c0c1f007cc0000300010c00000c00400c030330000f00000040c4d7f400040000305d030310741f04074c00000305c00c50c30110040000d7c413000d0037c10f1c340c3004030044c01041035003075cc000304000003410d4000440cf300505cc034000f01040000c00c001d0c43ccc003f000c040004003103010c010c0100003d70350dd0c3000100370c00c0f00c4c000c10d00303040030cc313c01f70c04c4300c00c3100105000d005100f011003c04330004000cc0c000014033013d005c013140c33001c0f0c00d70040104001f0dd00300d30c40f00043300f03ccc010dcc4c3c010c0c0cc000331407004fd400000c0140c3000000d1c30010734034101410f335040c511c3030403c7d3143300003000003cc00413031431400f30c4000004f00c004c00c03d001c00c00d040403070031c0073cc0c300c003cf310c4401c310300000003141040c000c070417003c1707c01d0440000140df300f0c3c34fcc000c03f13000d01c013d00d00145133f301000115c7d004034403c140040407401c00040cc1cc00500100370c0044f00c000000000347000405171000004c04100140c0000c0530051c3f00000c7c000c00040303000c0c01003000343007110dc30cc03003004050c04c0304734414f101000c003d340000004003c3033040030403f001010133114700d4fd030d0c0000050103000c0001010004d00401000c000411013304c0010001f400c001c300000d0c01400300035110c0c03cd10c3000c00001113c3c740c33c00370d10000010c3000041dc4c0400300040007000000f1011401334c000304c431cc300700000f4034000300f4c000c0340014001c300c000004d1f110000013c00040c44c000000050030004700c3c1140004000d7c03ff030033031003000113003003000c0c7703c0f70cc00000c0c0110010c0130071000000000cf7043000000c470c140300c444400000040700fd074c0500010000c000cf4040030000c05100c0300100cc04304000341d104cc400df3000400003431000003c003740700000c00300000017c00030000444004504c010c40010c0331000c7c001331040150000f50c40003c00c0100000030370101d00430400f300300033071110540073010431c11300000c1000435c030c0c3400ff4c034c140101c03010300000c000440d00c000000004c110c003c1cc04c0c1c4100c001040c004c300400f00040031000000d10f0430033c00100003;
rom_uints[674] = 8192'h30010004d0003d03d00100000f00c70c33c5000c0c013c000cdd00031c050cc31c0341003001101000c00f00cf110c01033400c0c0001003000d000000034001c001400f01010f004c0040d040000c003c00033d0c0f0c0030c4003405d030301010350f0c30400033030000000d030c001c010000c1004d00000d000d0703030f3141300f75000d000c103041310c003004000000000014010500004130030000010000133c47d00c0d040c430400710c30340400000d000000000075c0f0c3440130c000000100000000103004cd700040001c000400040100004335c10c0000030437030cc30cc0000017f03c0c04003104000f44001c000001c10f10000401000030030300c0004c04041d3c0c33d0031013000101000c4c0d050c0cc00f330cc00031700c1040000c014c00004001c301c0001d0004001c04003f010cc30f4c0101000014000c0c17001d010000000fc400010104c7c30110030c000fc400040dc03c0fcc314f04c5c00c00431f0c0d0c00000d1130000030c00d0040c0040c0f0430050000330100004c00003107004c0000003300f430cd0f04d0050c003cc004034043010003f0c401c40d040100000d330000100330000403010c00d01d0c0c00c0000013000000c300030005040031404d1137000cf1000331c50c00c0c00300730330cc000043040c00000f1c400043c3100fc3050100410130033000000005030100433010341014c30f0c0c000d3310050000040c01040040000c0401004c0c3474100c0000300035130004030c0c004c3c300dc1c7030001cf0d0c500030003300300c4301013730040000000000cd100304cc0c010c0c3100031c030c0f0000fcc00c4000030150077c34cc300003300c000000000f1003c0041100cc0cc00c00cf110d40fc0c00040300070d0f30c40f0001000010d00170f00cc30cc113304055040dcf31300c03110000c000333c000c001400010000c0030c000c0000033030000000003034000c00f70f10400c0d110004103c3c300000000c0457330c0000f4c7001c0c010c1000c070003c0100c03000c73c0303030d0005007f010c750c04000c007f00003300430003000000d0070000040c000103010cc1cc0c00040c1d3000000100003310451c003c00300c00c3431cc04c030300030cc01c04000001041c0004130043c00300c010000404dc05000d0034100f31000003000003010cc000330100000c00010011430000010c000005014c0000c0340101001cc00d0700c13dc301004040010cc0073f000f0ccc00000703004c00000000030f334100100c0000000000040000000030c0330004000101f03c000c01330c000f0000100c300300000404030d000030414407053f0c10c1003401000c00010000000001004100440f004d00104c4c04c4040d340dc30107031c;
rom_uints[675] = 8192'hc1d00000d3c7014000f154001000d03014330300ff50f305c0c50fc01133c3c1f010c01750f00c010f00004700004131c4004c4070c0307140430000137031c0c100fc40040000030000704f3c00404f3304c0c3c3511141c0f0507030131c0500cc1403c004340000407c00001cc00443404413c0dc1000001504f170000003f04cf00c300103cd00400070c000300040f000000001f0fc01c00004700100c040403010ccf1000c03401030000f00cc044030ff0000010030c04031400041040c00c0041700d1335145000030c043010000cf00c700cc7000c4004c404c00dc33040033cdf10c001740003c00050043c5c0470740f3004400110d40c1c00010dc00c344fffc004000f0cc4045c30400713d05c3f000d0c3703000cc00ccd707f333070003d340c7c000f0000540c070440ff4011530310003c03401f03044c0cc03d0000315ddc04c3c13001c1454f0c0d0f1dcc34f55504300c3c0140414300d0344c07cd000140f0c0310d00c0d40cc0101f30030c30004d4ffd000403400d7d0031531c4d040d1d000307111430c300001cc0070c031003c3700035031010c444030010001c3c0d01303040ccc0d030c103343000cc404c34000013fc700501000000f030010c3701001410cc0001f3c00740571d007c50043100f035004c00003fff370404430fc0330000111010004ccd0033c101430703c00304040f30c300033310fcc0c40cd14703c040c0034017d5041c040c1c030154401c13c0dc0c30540c3c1000000004004140043cc04047c0014c0c3cc4f1c043f00004530d000500f44040c504014054d00cdf0c300c4c1cc53000c40740f40d7433500c03c74c3001040003310c4d3c000d0000c30015330c0c4cdd374303c00cc0c00d77c101c00d00c0300c131433c000c4070007cf035c173c33c00c0010004c003c40004ccd400f07103f0c40004d0f37000cf4d30cf40cc0303c40174f00001000303cc00400000c107000000c30cf000300000154fd1104040044404000c33f030cd000300c0c34014000c400d00d00470d0300033d0d10000074001130133041113700c04d044044300401045700100d4403405400141c0c0f00f014c3f100340f143c3000c10c0c0cdd110030f030400000071c34410007171c3740043417c4344301f1073c10cc100c000c0c030c4c0c0700414f1cc0c0003d00400c0dd701c10000c000330c034c0405343d000c3c000040340dcc00110003100c000401404444004471300cc004511003f0cdc0143f00fffc0007c0000f4104c000105000d00d04000040050f0cf1000010cc00300044400030010737400cd0000703040c4c0033447c731c17c000310d7043003003071300400c300cc715fc0305c470004cc300030dc0430cdcf3510007000010010401300cc513f0444d0000330310c04;
rom_uints[676] = 8192'hc000000044430150cc0f0c30400000150d330000c43054003071103fd10c3c0000040c30d03000c0005d0003c04f310c4f01d470140040007c0040000d14c01431000c03000000404c000040f000d11014cf400030c410300370c1c003054004c00c04131c030d0400030500141d0000001731110c140ccc003d01100d0c0301f13303010450000f330300c03c10c03c400c000400404c04130c50300c0c1d104001101040c41cd000c407100c430004300040400000000f15101003003371030010104003004d30004f0050141f10c000d00c00c03c0c04407500dcd0cd00f013730c000400cc054cc50cf0d400000c000004000000000100c003441100000f300c0010f0004c0403001000ccc00570010300041500010517311c30fc70c30c05dd4c00001400500033c010031000d07305535100100d0003000040430000c000300d40c5000030f00c0400000035040701340c1100437000f310c00144003070000000f00030c1011400c0100c45054040f55340c03300007310001000c400301411410000d40333c10050d04100000c004000300114113c4400c330300c410f40050000d010430ccf3031000c3f40370c0c3000c0c10c470c3000411c05f010040c3dc70430c0ccf300013010c0100f1405404cc14037300c15c000cc0030333c00010304040110130c0330110000f0000401001cc000040c0000004017330c0500710dc0d0000430c00010700150030c10305d0134040c1001030f3c0570030c0f055105000300c00c300ccccf4030300000045403c30c04101004013c30c034010cc0c04001443c0c14330c0414500070fc30c0c3c1ccc004300043301005010044fd0001c0300d0c044010003f1540053c000540400f5001140c31000404cfd3c0000c50c3035144007c4c1f30cfc4445101350030000310c0c00403c4c3c40000f00f11540333110000331310c04000030130c05d0c4c73001741033030303300000003000300003110440004000034500cf3013003d03c0301f0300070000c333f30044c003030000010005105c4400373003110330000100507c400043040c0f74040cf0f000ccd001d00703300000100030040003000000300043000cc04030c7470400ccc340f30000040001c403c3c030014c41010130c0115101013307c00f040010000030d40cfcf3c0c000cfc0c010c3dc0444c000d0044000100000f300f000d50c0000ff00010303030403c0014c1c000cc0300300d0d30cc4400330000370504410c0130000cc0400300101050fcc014c4000cffcd40c0541001147100d010030000113103005c00c5c10ff0001040004c100004041151003c003c40005310001f0c3f34c30000010c0000d00c01cc01140411101434005100c0000140003d003040cc10d051110f0c10d0000cc407d00cdc0034000c04;
rom_uints[677] = 8192'hf0034401d1c00011003d00014004f41011300c5033010000000c003d1031000033cf30cf0c3000050c3414c413070510030d000003ff00100100f01c003d4341144f33330ff1c1c3100404107000040d3c10f11315c44000004f0001c30041d5011cc1f30000001f3003010d010f3107050040403f3030100c1ff03c110000045333330331300030c3001ccc30331110330c30000000000c1043430c0f300430010c3c000100c0c0310001000005133105ff311000344130cf30c43503cc10004d0000301003f00300300c300c0c13040430000003c010004d030c3fc5d0131000000000111000000dd004100d10f0400000c1000140000c0000030001d00c73c4100c010400c10741d0330d1c30013514301510310c3d1110c00cf03ddc3510033030054310c1133000003330301333300cc110301310003050313333c003003c1f341001040041144000300c300534f0033341f0003f351c0307c131c11301004cf00f73000d0c3cc0000f343c7400000010c00433034175f33c1c000d3000f11333c101310100cc1300df10010f304000000000043000033c1003001134000f0403f330030f000300104013cc000110433d0007000cccf0030c004701001000103345301001000f333300000f00dc133004c0000f03300510c0000d1103000f0c13001130001335013000fc000000001000c0004fc000c4031000c000c0cdf0050103000c3001031114d505c30141333c3113c015000014304553010f330400000c141033030003743104c00f300101303010013033400f033011100c300d01005fc010000cc031011c00ff3f71f00033c0001c004304000010c3014c7dc00000030050cc443000c705370c3503101004000fd0500300000300110300001303d000d17011100c0fcc1004f3000100003440010314301010cc73007c00cd3cf570330003133001043f30d3303000130c3f00f0000100700010001c0001031cf0051c000000030030400300004100f1033d3f5001004c31dc0135503000150f0003003330010330ccf3400000410c40001c03c003340030c007010c3034300f0301c00330300d3c010303100300000cf001301f0000010000047003004c0d0f13300014c300011000d400003c11104000153c3403001cdc1dd030300f0304031010cc0000147f33cf001014f030133f037071100403015501cf330c0430f7051d0330704310050341100040300cc1ccf1f403030005030003c000703003cc330c0331fc0000130cf01c505303033f403c0c000004077003f0311030711000dc0d400000300c00000103000fc01033c00104001f300004cc000d00011000003001030044c3033c030300011f05000013010f0c30001c040003f01cc010400001c10010101000030c051030310303003010000000303010014c000300c004105;
rom_uints[678] = 8192'hc43f1000303f3347337031035700077700310c3010100c0400300c00043130034003f4c00f4c00d10003040000010c3073c010c0433c0c1000000000000010c135001f0000c4013c0100ccc05cc3030000d17c3f0013f3d4dc300404c003f0040033fcf03300cc030300cf030c30c3c043f4d0000f7300cd000000cc0004504050d03ddf30030433000400dd100003131300000000030400300033000003000031dcc1400003fc703050710430c004d30031cc030000ff4133c00031d0103410003030d100000c03433c000ccf10550404310301c400441000010000c4d10040c0000170434403040000c00014304305c3307340000100010c00c004403000004f003f051c3f4c00c001033375c3040c150c0147cf1030033400300c050f01300300010037440030c33003c131340d1000343404300000000005040000c40d3003131440ccf30303170340cc43131104f073540c001c00fd0330d3304034d00010110c013c4330000f030c1f430c01030f44113013404f0400401f0300d3c10c30440044f333000003134033d4004331c0003010001001c4d013c41301430003c07131140340103100134140c1c01c300f003f3504010f733300100004cc30100471c1cc0f33c00000004004033010345fdc0330c3354443010500130c0043550000cc00040c040d04430343d3f330001155014400000c004000003c0403ff7f31050f00c11f3070001105f0d3c001033431f000d35c0c174730104104000f013400401434c33104003cc10100013c03013cf00001013c10c31311d01000300713140d0104d03000000014d3411313033000000f40c40441111c0573c05410031f31000113c70f3f30307c0c400300c340cc000f43140c70c130f00400537000df4030d0330030000030010007f5c1d303d04705c00000130005cfc01304c40f01430750007f3000c514c113c3c300301f30003013031440034440f3c70301c1310c0500350043c070300100100f3033000c04f10054c3cc0300710400401004cc0044051343103f00c0113c70f0010440c00d01407000003003703c304431c37f1303100f3100c4013103d0d0001043010410c503000f77015335100cf0040003c10000001f40003770c007000d17000001f143007cc007104fc0334015c00035f000dc173c3100300cc00cc001c000050140c503c003d04440c5000313c430010010c00743300030000031104070004035c300033c0000d03400f01303001031c0dc0400004300c1d00f0c03310c1f5003300304303c00f500033510d04100300000004003f43303101c10300400f0001005c4c0003005000007000133303001c0047300c373c00430c003543400c3d704f0153040c0334000c03d10c0031500304700703100143c04710530c1f30050c00443030017010340c03003001001;
rom_uints[679] = 8192'h313d0000c4050040cc3f40cc3104fc0ff00451f003100133cc00f0103003ccc0c0c7dcc403d10404433f0f01d010073fcc370d5c30351737c10133c0cf0f0f0000050305104300f001001014fc300007f41c30303c3fc40c30c317df551f00f003cc050034c1fcf013103315001cff734030700f0310cc0c00cff10c400410f3f344d3000c0334030c0c000330010cdd003403c000c0030033f00cfc1f1d0304c103cff4c4070cc340700304401cd00f40055333000104131f1010700f4c0000033100c4d0c1f07c000003030f4f00c500cc040100c4f04333044043005f000fcc00000fcc0c1000c00c0fc33f7403cf31004337135c000c033540033d010010cd01c403c3f34404c133003455403fcc5f4f04100f43c0cc0740d17c0104c504cf40d30030fc0d01000133050003c31f4f3c0034f100c00310013d00001300c351c1130143c1c0004fcc33000171003c7030340003070103770303100033031043f00f071f0d570c1cf01705f011131001c03305c04341030fc5d3c74c0077dc7714cc3c3300703fd00cc030030304dc1d3c1cc00c03113015c44c1f004003c11034030733f700103300040001dcc73c015f1155100c04f373c00c00030330114f050c5000f010c1c0c4030053700c0734003c40cc1c30330400c005004140f51005010000534400043300cdc04f00f3444ccdf701330c01007433c03700c4d1c4043cdc1300050c010c0f34300c1f3d00131340ff007133c073311c1035c3dc0430001001dc050343f03f0cd7dfd000350d4100010301cf734115cc7c40cc304073c0dcc11c0c03500d0c7031fc4003034c0c0033005000037503c0007014d133530000cc030f0004f1cc330010131f7c10c30ffcc01dc003401f37cc33c00500050df40300031f01c00d4f0d0fc033cf473f0c355c410c0004ff033d000c300030c074d01033307003044f0400300100030f3c101403cc030000c4c074cc010400550001003101dc14c001001310f300c0f31300340fc40153ccc0334ddc40c0004f40c10000403c100040714340000f03c0133c040c000d01cc30c04c1c0c313011013304000001010f0130f30107dc000100c0301fc437071700c000f710c433334440c30c100cd1001c73004300400d4c5d3fc10cf010014c135c001000cdff33007300013330ccc0d1cf1000c0d0010410c041cc0d00340c0c340030dc10f5404303cc00004c13130ccd04cf0140110045041c04545330014101cc0d071c003030c7101000101cdf1000c53c031004df3cf07fdc04c000330f0ffc10cc01107400000c040cc04c10fc115300f000f001c43d00104f43000000c4c44fcc010400c5c303f1c37c3000c5c001cc0030441440000000d30f3003c04c00101107100334300f1cfc000103df35003f000300304c0c407350333f34cc3c1f1f00;
rom_uints[680] = 8192'h3071000004300c03c0400510040100df030000000c41040001c3400d0d1374000c041700030000c3c3311750f017ccc0730400151c014fd40070cc00d00cc41003030f04004014f000074c037000010c1103300cc103100ccf043534c103134fd04c404c0007040cc5c0f13103340cf001c30400c1733400130034c303f10c41571543c704f0041011000c0033cdc770407000000000711cc74000077c4401014d00403c50f301cf7ccc0d1d04100043011f533001c3c370130050f3f1cc01107df14c54003c0000cf400c50000c45c7000c15c34f040304c0351010cd4110011000411103cf050030400541430100c4700cc03f11000101c0007c14343003440000001010fc01100c3030043303303d0dc01cc70740400d17743c71744c4cd3dcf00000300000030d0111d001170cdf4c401140370c0331004f01130c0004c40110137cc44400000000300c0c430131cc0113030f00301dc40750d7030cc000c355013400dd0000401f0f0003141dfc000007c411300cd0150c13430007f01cc13c430f50cc0000414301ccd41d1107d001013100033311c053040c4003003ff41100044c10cd40704c030400134000430004f14cc0c0004000137001d7005d1037000000331c04c000400dc1cd3d5c0410cdd0d10d3d14c4f0030453cc0300544c00cc07400d3010f0c0400001f15311cd03043c0c3c0113c0c300043100f3410130f1014040c705cf001130d00001c3c0107fd341c0310003c0111000d07c13cf1500304f07100305005000404303447c03c0031340000037541c1004113f004104c30000300c43f1d0400c1034037f3007007043c40cc1d41001c01771010400033413010004c0300fd11c310410f5dc3310c11400101130cc004400dc031371003300000010073400f400300fc003d0cc00c4c00143470700004c03130f303473003cc3043cc3011c0c43100cc05d1000f00001003cc030d5c04330000331c430005000c10103400011311100004f0000c03c3f0444004100c3cc011331300cc0350000cc70041fc4007cd004c071cc04100040c0d1d545307040fc030051d4000c3c03045004471c0010d31cc4145c01004005004c3c0cccd41303300001f00313401fc047000504004434c105f300f5000310004d43100300037111c000cc0303133400c30701050cc500fc134c4000010cc304cc007004c43d0cd40c3301440001d007d010011004001c70004531130001cfd4cd043401000003130c041f0c13400ff07cc0001f0000470700030000004330000c0503343070000007400c030c004015000c70403c510733400f01c030c00400cf00c0000141f5cc00043c370303c34013010004031010100c141d4140030401c4c0010c3dc40104040c03c5030c0dd01045033000d04000010f00043101cdc0c3c4c00000003004c;
rom_uints[681] = 8192'h4144400c004000030057000043cc03474c004c00434050140c1c00c401c07404010dc73c0cc01c7c0cf003fc010004d54cc04cf43d0c0030004110300000050c0003434c41cf4f00400300454000050c04400f4c31c004440c0344014cd1cd00011300010070d470134c004440c0130c40d000103c4005400410000c0014300c5100000001c4c0000011044000004001700c00000404c030c100d7005000c040440c00400370400003300303cfccf00c04d500c003017f300d0401004400004000000000000cd30c35c000103000344704c004010011010034d0c440c1c400c0000000cf00330440004004c1cc41f031001134414100c000030100010004034000000000c304d30054cd0d0303c10c0dc30c000dfc30400000000c30003c0f0007000000c0100c0c030300000000f001300c050300cfc00014c001d10004030f3c000cc3c10c000030c313cc0f010c1c0d00400c031c70450c043c0c00540c300007d0004c4c0003010c30001000d0403c300c04014cc0100c3d0030000c10003c414110d1fc010404f000171c00000c1000001030c0410000d004040300011c130c00d04dc40000007cf0400f0300c0c0050c4c040143004004700c030c03001c0130c341700073c4430000301c03c314d01fc0440400030c00030c03030cc104000cf3010cc3310000010d73c0c0044030c4000f0034401010000030c00141c1004400c0010400374000405cc410f3d0000c501100c5401000033cc001370c0cfc0c410040c440040310c3000004f00d4f0100014c7c030030701700040c0133100003043f40534f0535310f0470040c70df00d00c0c0403d00c54d3c13340031053000f0000707000d005cc1404c4c000431040300c00000c0007400014751c0c030100400745045570d1004340cc7540c100044c0c003d30c0030cf00c00c0010d757f400ccd00441f300100c30130cc404f0c440003070001014035004c0010004100003405c000dc0000070111c04c0c100000f0440170c3c0000034c3000c00c1c30004310c40040010cc0010001f041300c044c44003430747300000f001404301040013c00ccf0410c040445d03f7c7030300030040000000c1000c03003c00c00c05010004cc0c103c01000030c0c0750005007cd3d050050f000003131440103043100c41401110033c44107c43c00013411110c10f0030001000cc304f000f700cc0c403000004410c4c710cc00400737c0534700c000405000140001405000c400d03103c4f03050d0c030300c5103300045043300000d004014300c00f400000c040000000f01fc550030cc31df0013030030fc003434f0100004301700cf10cc0d001c50440300c0010cfc0c0010504010f0c0145c044400c03f534405043034c0c04140000401034c0001403c00100010410c3430030010;
rom_uints[682] = 8192'h4f030000050440df1d0400330300000000000c070c073731003c0030cfc1000d30000c750330000030f03000010004c353101000cd51003300000010c4d0cf304f0c5504000004d703003444dc000040040000c00f0c000c0000710f00c5300000100000034001030034150000c37103c030c010000310410307335100013003010100000400104100031414cc0100001031310400c00030f37c0007340411000104030000440cc40000030010c010010004043000070707c51c0cc10404103c00430010400c01c07000043033040010401005100c303c33c0100040303f0c01007c3104010700000304003c0300001030c0fc0c004c0c00010000300000000030340f000041330430fc3314010003001344040110cd000f050c03f7c0100cc0000000000303003030041040cc003c04130f00cf4c0f000001000010444550101033c0000c43300014ccc0003c00113301c4003000113c13f3c0cd040033005c001cd403d1010310d004747c1030c54400001403000433000170041000140050001543f11033300c7c0400c00134dc01f000c300000431017c14130000300c110001010400c3d00c000c3f030c040000010400d0100070001000c7300c01c0f100cf0000c0c330030d051500700007003334000000310c0001d0003004c0cf00003d0c050c07010c1000cc3000d50c011103c0001d000340003001c014d4107001000c040d0c113f00f00c003c31010030141100cc0f00034c0314001c5c170004c0070003510003000c000000010c1c0347300c40030c004004000d30000001c010100d0ccc000010f0fc14ff11000407030c5133100c10003c0cf0cf0350370005030101000003000303140001043003000c310000c730034011c010101000340cc443000c0001c005000000700300005057c310000030000004007c00000044001f0370031c00d00c151014300004c03407000340dfcc00000c44000c30004000300f00000003c3033001c01434000c00510c53300040d003c30310d300401000000c3c00cf0000150000030330c03c001101c00111003c00007014130c000300043f401133d1fd00010000dd0c4044330000101004011400000734003c1c100c330c04d7031000300c00030000330004001c140f300500c030100c1700000c00f101135c001133037000050003003f005001313000041cd0cc010500000400000044001700043d300710d10017c00000c00330004040400001310004c4007304040333015f13150130f411370d30003cc0c31c3134001c0c0dc110fd0cccd00cc30d07001004d10c0001003c3010100c00313030000703001000044300c70030000d300003050000030103030cc0001015c3000310413030100000103410100414000000004c000100000000c5033d110cc000000c0007310c1003000000;
rom_uints[683] = 8192'h43001c00007000c40044d00c50010701730000305140170c0077c3c140dc030000f4d10004f7001c13f1c00c30c0151374340000004710d10f700110f3001010c01c1105004000031100d0045040110f330f40303341001040f0101cc0c433c00335c0c4f00300d01c43100c0c30f03010400430347530c400f0014033fc534007d100030c30c00400000155d410010300f400000013ccdc370f04330c75d0144f41f030c0d104c500531010041000103010150f0000cd73f03000c1c4404cd0f33d00400017414df57300c5f00304101040dc3000033f1cc7cc11300c0f00c403300000c301d750f0cd3007407000000f30c04044dc0040043040c07033033c00c3cfd003007403c413c003dc31300c11101040c1c33400035f40730ff000f01c57040000340000c31c400f101070c14730000300000003c3301004340301f310f1c44443f3f33014c103511c043410df3f13373504034d30d01543400c3c144f040000cdff400c45c0c300041001113c10000300f03700c00003300045cc035413f034071cc7033334f0401d0054c10100d11043407500cc0403410043d034c00d00005034010c00ff300000c51f000300415ff07304f0400054d010c4c0313043400d1c431001cd333410040370d3c430000000514711c1c0100030c00034c70d003d13dd0c400000030fc033c04051105371c0d0034307d0c000335c014f040000030073c37f0cdd00100100004d00100cd077305311c310503c1d30310d0047d41103f00c4400c00700d30c303cf0c403c00dc011040310c004df100007010f0133c0010700100013545c0105f473300100001c30400047d03441d4cccd45c0f003444775ccc13c33c100c1100000010004301c10d0307000000004f040f10d070070c3000c7101d0000f1dcfd4100351d000d0005440c4334040dcc1c000010305704074c000d00441c500133dc00170000011037c343014f303c430dc01300f3100003000ff0c00c10f3100f0033033cf00500ccc3f500010010403035100f31fd0fc030400d100307403cc134040531d0f300000cf733030c1000130340cc0334070c500100030301030403010c0000c714000001014100cc30130130433c00c1cc10c443403000100331300000d101510fc0000113430000317d1c040cf3f011343c041c0307cf101304330134303cd00c03c0c43301c000040d0111300130050000cc1141f04c30f3c31103400c0000001037d53d40013330000c07300c500c330304111c0701f1000070cd74cc03303030c0c0510300f5130d000c100031070344137c0740034d01000f0003000cf3c005d00000403000140047400100f30301430dd1000c03307cf013403341c0c44cc310440003c11310c0c3c0000000000f304300073303000fc74c000000c010147100ccc31c30034140131;
rom_uints[684] = 8192'h703310f1030141000000d1c1c0133103030041cc005c050030310003df0d000001330000000010010cc00010103c40570000401dc4000130c3400010013000000103701010030000100400000340c001f33411013f001c4340000033000000001033c1f530300c014015700001f14000000000403f11f03c04010f00c0c3130030033004c05000000301134f0301030700d00000000341ff00703007c3000301cc03c0003cc3f0030d1000c0c01000003f43303003c004d0c40010430051d303c31300d000010f0c3003f1330f04d3431370300105013d00001314130d100000043000003f0031000f000d40d1401010407303000300011c01c0403100001d0303007005304000030010000311c000011fff1c100dd1300531c300010504000133730000413010000350c0001001104041030003500100400013100300000f000c0f50101301401050c40fc0104003033100c000003301cc011344000050003403340c034001130300330101f140d0130cd0100303034303101500000041400011c0f03c30dc10100c0033301000c300c0030140000050710031cf03c1000000001100c0013c53003400104073c1ccf040340f1040004300330370f1d00df451f01000103031010004003001c000010730fc00030304c0c001110010334050d754d101d403004f000dd30133c0f0310341d0c5013133001001c070003010040131d04c407cf00f1d0003070fc001c33f0301f01130000001cc04c014d410411030df301133400000000fd007c303013007347000110303030050c1300003440310dc000cc30005430c1d004f00f00134000113030000000cf34c007300d03f400c00001050400d300501403c03005400f3010030000c0000004c0d00c5303000031301000010030000c0011c00303001f3010001000345c000373300f1c00c11c0010011c007031f430103330433503540c000031c0c00c0040fc130370300405130000030001000103007001040003300f0c703f01050f1c04300c03107c030300c31dcd00c037d0cf001000c1f01c0c00113010330430000034400fc5fc00131000041030c077cc331c4007043c33700003300001f3330030000f1c010c000fc0c0ccd0030443343034000000c53030fc3441041300131d0300001f1c44400d537c43133014101304000313f07034400c3000034400354110c10041cc0010c1010d30c07100c30f01001101013f100040c0103134c11c10040030040000010100d7003c00034030403c0535300350003003df000007000530111c04400037303010313130010f00050030103000cf0051114010101c00000334000100000311310c4040340f13103031300c0000004310c30c000100010101141000f00f0c1c0c00570f30305000053703010c0003f100013c300010fcc530001003000001;
rom_uints[685] = 8192'h11100000d000cc00c300030c3030d10cf7c000400cdcd1c30003410000040c00007cd0033030000c1031003300001d3fc014c03c00070035300dc000c000000000d1077000000001c100c3cc0c00c303033cf4010c000d0c040cc04c1303000303034cff5303c0003000c0000014d3c701c000d13407400c10040300cd03400010c00700cc0000010f0303c33300f50f3c3f003000100104d01300000c0c40300cd403700000f003343774001d4cc000c000f300000400000007003034000c400cf003403300403074c3001103007343000407c30700003030000000cc1f0000000c00c00d0d303033dc00440410c0c07001f430433c140070004c04100000000101c1040000070000001c00303000003f000c0c001ccc03100100470ddc7300033103003444000030c0301030f03cf0300c134c30f5000030030100057000000130000c00000430d0c0003101413700034c43030310301001f40310033fd0001043c0f300430c0000353f1c501433f0014110053700c3300f0c531301000000705c0377030f00000d004300f0034f070300300dd00003030003043c00c0000d07d31c7c135c00033034000014f00dc1c10003400c0c4f03304c013d4005c1003100100f44c310c0011f0000c00c00703c030c04330045f4303030c30d7c30c3001cc10003030cd40c4d034003d004d03000303330c0307f1c0404040004c0d1000000c4140413f303f00003343c4c0401030c030313d40d00c00300c03f03c0000c303c313003000c0110000400000013c00000004c3041ccc54374100300d004400340c707f00000403144c0040413000c30c140430c000c1d000334000000033c3030fc001050000c033c0c0304173405330c00013414c31403730cc0003cc03c11f03d4f300c0307074c3cf413000d003c300004004d0034130cc000f7c31d004330030c0034111003307004040003c30000000040f43c0c0f11103140c0f03c0c301c0000cd0003000000c000000010070fc0307c00100000310334cf01f30040033cfc0331004c00034010000c030c003000033c0000cc00c00074340174c01301340700d07d0010c33043007d0c0040007330144f000001d01010cc3000000403510000500c40313d10d50000040100403037001030400cc10347013030070c40000c11c30005c7007c30c00353c00c4f01d400c10c03c3003404300010004010010c00005000c0c003003000730001cc40f4f0fff300000005f04100c3033437303000404300070034030c04100c03504c300d0314c1f01033300043701c0c0337011014041003431c70003c0030004014000cc010300f000000c0500033003030040cdc000c01337304000300300700000c073c035703100010310c041000c073c40407011f043030051304400f3c40013131cc00d0301f040c3770;
rom_uints[686] = 8192'h10f10030d00c701173ff010d03003104f10c011110303c0000037c04403040130005c0c530030000f0001100031000333143074510750f00400330300003fc00c1c440050010411030000014030033c04d31c0c00d0c10003003033d005430c1033c4500031003c0c03d40f33c0f30c410c70000105cc300040c414101c003303c003d00100f000f041001033030c00343f000000000f4070d003000fc317f13c4fc3c14f013715f000c01500003700000104010004c000010c3010413307000ccf000110d00014714351003003014c100003f54040100c105141004fc100000010c3031030330001c30001103050c1cc40c00c3037d10014000000470d30010c14c3c7005c317510cc3301003100400f4fd00001003f5005030003cd0ff155103004000c31100cc04c010f154043103051030331540000000000730c0010055f00003014f31c0003043010f403001304c510f10501130411004400344043c03cc7f00400700013000300005010307f43c3000003c000c0c30054d013503157c1010c150034010343001400cc3000f300300f00000000404014d000310c473c0d30510715051100c0000010c00103030c03f40014003004f440133301400cc01051030437c14000c0000011430000000047c0534000c0c13c00714047043c3100f300003041f543c70c3310014500035c0003c00400000044c030310100470fc70030733107f000400f03c40ff17003c30000034100cfc3001030dcdf37115054054f03000cc0040000c11010c010c03c13c04d0c030cd1d00c7415431000cc331c33350c0000c010c000004fc001043000d00c0cf00400c103017c11004c4f0701700403f110c1030000150400030030370010c001c74f10010c314f0d4403000fc40140c000430c1c73f703fd35c540c0033000010033c10003c033fc7170c303cf43010041fd030c000fc1100d413003ffd07001c3333173000034404cc33d031c40000003d0100047000030c4014330074c7f3f14001110d40f303c03cf001000104c0cc000004500100100101733d3fc0cc01c400303d4c101c00d3ccfc510000c51005000d4440030500501431f070000014001d710030033c0c0010044c1c00070345300100cc45000c0004001304133f040c0c503c0143000330541410410300d0cf0010c0043370dc000c1004f4000c0cd0f00f30553140c00000d0c4703cc5104c0c430000000703043c00503040f410fc30c357044005c03dc001f101d3510d00fc001c103c30f010cc1300304c337f03001404c7c434005c000c47001501c040404c0031414c43c0300001c3d711c10143f000cc00000c004f0110d10444010f31c01040534d00c30033044cc004000c5c500333c103d47c01415c0c403001c00c017c00304033305040fcd0c10000d0137c303000104c0c0000;
rom_uints[687] = 8192'h40d1000ccc5004cdf1040000030003d4013704c30cc00f4700c71c0030c40cc013030741430700000033004040041cc0cf010000301f03c100001000cd033517015170dd03030f44000030f701304dc0c300001d0c43110f010000c30013c401403105001440001d43d00701d333133100c341134013510000c0040713003d3c3047300000d7004c00c100003700443d074000030014c454d107f314c704003010c07130015c5d00c00c00dc00700fc700c05300000340f0c3500300c0dc0100c0034400003000cf000f00c0c3c01d00174410031400001710c10c34300004300003f00001000005000500f4001340033cc00000044401100000001403400c0dd7004400c04c50c0c030c00370033003cfc70d045dd7d310045000c7030c3d01103c3c0004c5403000000000340040c3c31303444f0403c1c0000003130040001f30ccc0304153000070004cc14114007133c0cfc30100c0c037344303303340d000c334ff1c300c01144045cd04c3004003004440c31000005c070000700030dc33d3c0c150ccd700c7000c0f13f0d030000700d3004c17044310000c1450000313000303f0c040000cf0c000044030004fc00c3fc3070400004041d3cd447cc40c033311040c4130000f3014000004c5c3c30140cf0114010c4000003d003c100c0d3300c3cd103037310343ff03040c00001334f3c010c70100d001031310c00c000f033d0ccc7c073dc0003000437405c001cf31c05555f340cc0f40d7100dd4000c014000c0c000cf000030c4c40177c00d110041cf401143f0d40d0330040100000703030000c00014c3c400040033d04cc3000c00004c00c400300140c054010000003c0c5040400000000030d743cf00d0700c0070c00300c4430d00c73d5c1000c0710f00cf55c05cc31cc0cc0700c003150cf0004003007005c40c37000103100fc00404001300f01010c044c3c0c40c0310300004300050dd11044f0000c14000471010103441000ffcd071c0c3c341c0c04340d0c70133c31d0440000010c07703430000003300c0041cf10043030403100c113f0f03400044ccc1c40515005000733c00030140c0134107c00000d030000003103003070304150100005dc013c04c0cc10007c0d1cc0100707430400041c010c10cd3d010c030c3010055004150d00447007134cc3c4c071700f10044037dc43003030c0004c3c000c003cf0f007c04cc30c70c03dd0c40c3c30c01005c015c01c000400f00100dc00300c000f300c000c1cc1c001300301103047013c1301c40d017c000cc01c10cc01f0c1110f311c00001410c4c430c4100000000d00c0c00cd000000c3c3000c34df033c10d0000c330cc0400070000000c300cd00c004040c3cc113cc034c00d40400040050000143f4000dff40f0000001003003010c4c0110c0003041;
rom_uints[688] = 8192'hc1f101104004344000c0c00c7003c03000005d0154f001c100073c0c44070001000cf10fc133100000f4430c40050040350400c3c00534403001c4413700030d040f0f010d0400c00700100774c0444dcf334f334c00005430d30d7300d0103c1c01d3c0dd004001f333040d0c33f1130003003010c04000001131c00301437447c0103000343100004000d0c0c3000fc41cc00c00c1300c1034000c050000c04300dcc70c5003030043c30000c040c0c3c40500001001035001c4fc3700310c33f304370003c044000400c4f300450100c4cd03c5cc7400cc0413f43354010fd40013f0037030007030003374451440c4017140c1001000040001c1710cc010f0d00c0000100400004f00c04fc43c004447d000c400f1304c01c1310045d140c1300c0034700010001010001401c301f5043d04030001005c4c370004cc0040cd43074050c10c04340403f01c04c0770004010c003103c44003c3150570cfd00307f003c15d043330cc440103d0c000004304010c00500043d017400144f4005714405c001c5100d303010334c10310403001431000d0c01c11000003c00000dc0504d0330001c400c043c0c00f43000110c053c4c5c040c04341c34010dd0fcf5301c44c010c1fc30f130000c4d30f3cc0374700c347f0000104000c00044d000000c333310c44c44f000040d403c7445044c70d00fd01d70c010310c4d31d000003c0f044003d30cd070330d43340c040c05005430c3c4c04304cd710cd404003030400c0003440c00c00c003000030c0c00c310c0307d3c000040c00c530f0c004030f030004340c0ff5f04040013400403000311000471c0407074010f3303c00d0010010f30c00c00045034000730c031041400dc001041400010c0c0fc1331033c4c003c1040f317300c0010f00c073400370d040043d0d404c30c300c44034440110030fc0c4f434c3d1c043010c0100c050350300033401010040c01000413c00000c003101000f30140335004301d041f0c0c110044443c4007d43f300400cc000030000f0f05444d000ccc743d3f00c0c0110cd1043d43040fcc000000d040305c3c7470000110140000000dc000701c0d00cc0300030c00c450c1df33010fc1000c4014c10031311500c4c4fc40f043d0100075cd0440c34030001100300f7100100c00300c0cc04d300f4f44033031cc0cc040303030004f0c311000c10030700003f00c3cc7005301c13c0d771cd0350cc130001c00c30303c0c013010000000450353c000f33000c1f00c0000051df00000c0000040500001c55340f04041fcd70c0410003340300500010014c000113034000000470300340353f3cd0004c1cc0010114c304c0073c000070004f04fc303304440dc45000c00cf0100443010cc4c5000000000100043100030c40344f3f1300c004007d04c;
rom_uints[689] = 8192'hc537030001041fc17030c4000c000cc40d0f00030c0c343cc01d30300c3cc10400c0370003034010c3170003703c07400c3010030c030013030410005f04500c1010004c430001313400370d5000100011100fc4034c40d11040731c0330043001340c0331040304040370000450c034d0400007043300dc000c043443cf10c03c40104004300000c13401d071030c040c00003000c00040300f03300f00f00130501d15010c0005033000013700333c000f00040000031334c033500301030030cf33310f0031730d7c004404300010301c43310c031c03413030000c43c0001c130c3c7d0000001001100c04371c03c00dcc0d00030c00010104cc070c000c0750d3c04030c141113000130113143100d10d37000300c3030011c3d103c0000414f000ddf104107000011300f000c004043000300300001c004303c03c000140074f0001c0f0305343311070c14f0001c403100711100cdc3c00333c34040c0c000cc004cc401c4c01ff3f3100314010505c0050d0071d31340c0000010d0c0404f3300c30070cc3c3cd3c3030100d37100cc700000130000c13103300001113340d3330d0f031000c0f0414401c1007030300d4c001fc4500070c03313d73cd01101511cd305007004000dc4040043d0014000f0301110c37003041017317c004000707c44010040411100c300c435044c00d550c403034031c040074701704010310f3000cc3403f00441033075c43044300f400400010f0c07f300f3f31000700410c3c30070471c000001330c5000300c0007c000014003003510010003c114d30c140c0fc301410c103d01401c0073070301c4300001000010c131f0114000cc0510100151007350d04000003c30305103c1444300cf00504c000c3fc0030035151f00d43103c003414c1c0347c30d7c03031103c0003dc001003c375d751f4000040ccf004cffcd07d110714cf00fc1c33050314050d0f05030c4c5470000f003000f01c3301000000400c0100110004033300df37070341110313104c003303c00c13000031103505100c00715435cc00370000cc1030c0c000c00c05000313c0fc001f1300000c03c10c0d15001000400000300330404c100000000010000c053f300003113050000c370030010c75000d31011134303030007700d3d3c5310401110cc0350c0c34101d0003304030d4c4334c0004d4003fdd0304300f3c1f1073004c0073010c3d303cf404c403771c403c01cc004000300351010100f000300040cc14f000000d30c15077f430170cc55100330001005d33000c300c040030300034003c31000500410f00403300d00007c0000c0c00003000f000341700f015f30703004003000303444340011c03100430c73cd000cc30c01334c0400dcd000d4f0cf0c000010df000f4f04c4400c0075c400c003303000000;
rom_uints[690] = 8192'hc30cc10cc30c10c0040010cf13000c00fd0004045300340c30543000007d0300c003dfcc1044c110dc00005041c1c0f4c455c01d33400034340304000400c0cf0300c44f0050c1c040003030dc0000fcc0033cdc3753c3041011c3ff0cfd033c0c3440d43c031433df3030cc0044f03c0c0430011174ccf303f1001c3431c4d03d0ccc000055000c00c30000100000004400000000007c54cd3c41003f403010333030d7044d040743c050d3c04c00400c0d00d0000077c0f4cc1fc010030000130010430c004403d00000541501f0cf0c0000fc10f3fc3030701c34cc310f5c0051000000001c331c04007100c3000100fc34fcdc03000050c0013010100705f100cc03f03d5cc40000430100013400000d30c31104f3ccd7401c01051340140c33d00030cc034d407c4cd00c033c3f143004f333340400cc003c0341034c000c0c104013c003010010cc0770100d70c000040154d01030f03cc13c403000443d1c40043000350c400400c017c13044034001000050c0403010fd0704134400041443c1c03100c47c5007d0f000c300100003033300000073d0c313ccc440043453c000cfdf0c03c0f0c0f0f1c0c07c3300004430033cc3130c0c30300040330400014c130300f0f0fc0c0043007d04030c330130c030f0c000c0c0ccd000dc301cd340004f03d03710f04f30c40c3314004d0c341000fcfcc00cf1d0500dfc0c300c03010d00030030304c0f3103400ccc0300c0000c0ffc70000c4c003340001151033140c0000013c300cc001fc0013cc030c033434000100300f00010c3000700ccc0cf3400c004700700044407001010c10000110cc3c3170000410007017cc03030c0051c0710cc540d50c03df40010010c40030c00c14403340004c33c3f000030c0343c704000c30f340c01033c03c3d0f0001c00fc400000330d007d0c031ccc3dd170c0fcdf101331d040c3401033c00f0c01003010f300c00cc13330300c3c00c000f0003000304040f0c04f3070450c403cc0100c30040cf7001300c0317d00c0040cf301341010003073c3c0dc005300f03f0030004c01f100d4f0331c430c015f33000030cc0100004c30c03c0300411030cc0000cc43340131f03004070c30c000ddf0030cc1030001450053043430c44c0400034437c0003100f010c00007cc3140073304000030ccf40030100d307530c70044000dc04c4000d37104cc000c103f00334303100044334d031030d053070300003c03105074c341c00c000c0054c130c14cc10dc1c0c000c0c0743300cf0000300c3d0003031cd3fd04003f100000c01003c00c7300f10000c0004334c0003300f030011010030030c054fc14c33144cc050cc3f01000140133f010c0004300401130ff01c40030000500f0c3000040fc3405d5305100000c0044c0c0f031000fd1000c00;
rom_uints[691] = 8192'hcc04cc000f0d5c4ccc404c37cfcc1c00cd3100cc4010f34f31f3140001f4c304070150c531c3004c4c3004050307430304c0400105000c37d10003d040c00444c05c373500cd0430030010000400fc0407100c403434033007c40d070f01354c0000cc7000050403100cc70dc003474003303c700c3d044c00130030034cc3f0c344000000c300c1c404040030000d53c041c030000400c0000f3334503343f0c17c7034037cc3c030d00cc70337f1cc0000f30c00005c01330010f31344001100fc0004110033410c01000fc3c400cc0037070103400744c4c00001cc1005010400000cc0031000000c00f40ccd00004c3cf0dc50f340f004f00100fc0f000034414c4044307d57c4000ccd1c3c30c0f03343c3303d000054000fc1fc0370c004c0f10030040c5ccc0ccc0fc00015d405300fc30c30000103001c0f13dc11300c40010f00501c000303c0070310c04f30dd03cc0fc40cf100f1f71c003dc710100031c143030134cf07c00d10c7d50c03c4c3ccc4334f07fc3c0700c337ccc70dc3030113cd0140004f000fdd00c330f3000c3f000001c10c07000744c130f44f00cc040f0300cc000101030303000013107c5f333d0510cd733f1030d330110c31713cc731144110544100fdc0c000cc5403c03044d40000f0110507730cc1fc007cfdd170140337c3cc000d3034c17001f0c133c340f1d74003000fc30c1d50c0f15305d004c10100105310fd0410c445034f0cc41d13030c0411d1c3d40d07330300037fc03700ccc00140007007104c00000c307f4301d30537d40c40030000c134000f3303000d347330333337041f000070f30000ddc451103c145f0143c000000cc40c034c0fc33037c0c0473c03cd030dc3c34ccd5c3f004311cf054401df0c303034143070040043cc0cf3f4103301f0f7cfc401344700d40000c0c000000cc5055ff53f3001701000c07cf00014c0f30fcccc3044c05f100000c03d374f00cc00d000c13f00301c131ff700c3010d0f0d314c030cf0d3700007140300030dfd0d003000c0044c0f41fc4110001034c13000005c13cc3300c40050c044430c35310040d4010c1c04c0005040000530000c034f00c3c0d15440c1005330004c7010cc00f30f30c03c70030430010c0c000434043f003d00c1cc1300c1770101044f013d4330c103000000cc04f10007030f401fc01c0c0001f4f4340f00cf0c33030ccc0700cc0dc5c1c10d310cc0cd3c031c0143c30004cc15005c5d47f3040500543c3300101c030443030303000f004101301cdc0c01d0fc0004310000c0dc4315f3000c040437f3040300cc0f410d05010d0c000000f130cfcf0c4fc4c104301547030d7f41071314030330030100cccf440f0d1c1c313704d433000400340f07c700175014cdc1c305c000cc37f303ffd40440303c300010c0;
rom_uints[692] = 8192'hc03401c0300f00c03c0c3c41110004433d0000040004470d000d0000c330300400070007173f0011cc1400030d4000c00400400c100005d03cf103c030c00001d01c430cc04100000c00000f4000000303c00433c4c1331100dc10c500053730c00043030000330c05c00001000041cc1004100f37030470034c30000c43010051005c004030000300000c110c000330000304030000004d30004c10010041100d03003000100d03000004c340f0c071c0c3d00c000300000300c0300c04cc00f043000004000041f103000d0400c0d400331d010300000434440c0440cc00144430001dc11c100100c00000c7c0000c4000000000040000000101c0033000400143010040c03343003cf413cc0044330c131c303c00040103c00c400003c1f001340c00343470100303dc0c10000404000030004410c50000010033300d00c110d0343000053000010f040f0d040c004100040413c31d771000430000c07c4c3000000000400c0c00100cf1173404dc00000003d11303c0307c754003040000d0c40f3310000400c1c000400400c5401c000000000140300740c34000c30000c1c000040d03005100350410000d3f0c031304dc3f1001300470dd0cc14f30c0043003000000000000001001c33041f004040700c13c30d5003010c40cc00301004d0f050033000f130343000d33000110c0cf03400d040107000d0fc30c03c144c0004c0130003300100000500c30c04c0c73013304701001300003c401d403cc34130ccc4001c3000005035500040010030c0040140300103105c130003f0f00041741040003c0037110050f100133401c0000043c0301030cc0c34030110700cc0c0c710c70c00c4000000000c001d07f003400f1d014010c00c433100d4414103000c4030c00310c03c7010040030014333c003003c1003c000300c10004c4c0c4c044530c0047041c011470354c0c40c5030c14c0000000dc0101000001340001003000000004000cc0c04f00000010371003c5001003c0f300c0c00007000001c300000305100c0405300000f00007010c01c0000f050c0d0f1c000f00c43101400433433ff000001c00fc001501404000000000030fc00300040040c301c0401010100cc3004440300043c300304030f0013100c0d0010f3343c5000cfc0c4100d0110f3010004d3d03c0030014013ffd43c10070070740000004d4c4000c400100c000fc40c400030d0000010100f0000303c304c10400034c0d0000d000130007c010000f0000130004011004000003043c07304f000700030c00f101c007310c03000300c3c50c0c05c01000cc00000500033c0000c0000cc00fc301f00133000c070c0000054004c000000400000000f4c003000001137343104100000001c14c0c00c0f0030101407300700cc0033070d000137003d3c3c00cc1;
rom_uints[693] = 8192'h54300fc040070c03300104070f031531f405004d3d00100c035ccfc3cf350c143041c40400d300c0051404417513c70175c003134c10d0103000c11cd7000f0030d0003007400050010004510c0031c000304033f110d1333110414337f4cc0734cd13000310050100c0340c0307f053c001f0f4cf03033310040000d05310003cd011305301000000400c73d0d0431c1100004400000d1030305dc000043c13c31500101d553f7100131c0014c1330c00075f5700003030f4c00035450c1303fc4004300341dcc01c04000001001cc300101330c5000337dcdc0403331103000110003c700000000000003500374104c004cc0300d7034304034c3034100000f4c50404f3307c7300cc00370034001110f101343400f300f70c050544dc010f04c330003d030005c01040c0370041300101c01cd00000301303d0dc03540c030010301000c350300cd1001c0f1003c1c43ffcc001c30030034c1007c001f01033c40d1fc5c0043700004307c30070751c551140c7001d00c3c7f70c003105cc05303d300130c03007340c114000031351001cc0d00cdc00041010440303411cd03c0300330c305f004d3fc007d00401c3cc71003d1f03514000030003000c03403c0d74cf0730401113010cc70004004d0030014434c7f000030000c03004031300037c303703cc0c3cf73f030700c04070117733010000c41c000403d14033103300f413c0330c00f030740cd00047d7d43f430030d0c0f3411d0040317443c000535107d100010030c7011730030707d4000000100100cc110c41400005c10113310030340f34d01703ccc04030003040030401f0cc0c40130034c0cc1c101d3000c01100004400003314c4034cc0000071033071c30300303300dc41cc13300c034c0300104071c0c000dd413705043f01000c3015c04004f03013070100317d3c0c3c44301d10117000d700c0040013440133400c50040147070f3000030430d10000000300f3f0c0130075034c00003c40d1c3151000433410400c130310000c0717000fd000d73c300300c7030007000000000100cc330f0450070001470f400340000d13103000040c00f0113c3f01f4704004d431401030f34d4014313400c30c70d10c0003d00f01370004345004c10130000041170401c30c4000310400dc0401000300013fdfd33730cc03c0f031101100d4003d0100000d01010100c00413440030100f1140cd00100030044103fc1d3070300033d740070300340c10130000343d530010cc00c31103d3100cd43c0000300f1df0c0410100c00337000000547004cc003371f303c0030033000714013d13000403000101f1430070303c0443cfd5100445f300010300030c11043dc00004030c0c4cc3f0104400370403335d0300d3030403cf0000100d4000c3010003314115000400331304;
rom_uints[694] = 8192'hc000000170c300c0333d0070030f10000000cf0c10d000030f00f010c31c111f00f330d0100030431000010111000043c0413cc0d000dd3c0c0000700c710c7043c3c000000000000c0f1c01040cc01f1003130d0100040400c0704000f34103f30300307010044d03c04cf07051c31f07140000171700313f4153c0404c000000400cd0f0c400c01000103400017c300300000003003c045c0000401f40103cc333010104c3030000ccc0000c01100050000000000143c03040040c0001740cc30043400001d0313000d3011000400030413f3d435005f005c3000370000c44730004030040f03cf0011c5c10440c03d3013030010001010010c03000000053c00401003140400030401c000000010c503014c700100cf34003034050003041000000c04001003c17333c301030d0070cc1104cc000004c03dc44514c440c0011d01c00700300f1031530c30000340f1044135040301c1cf1043043003c313d0333000cfcd300110304734100cc10000f030dc300c033fc704000c1c041000c130400f0c4103130100c003000743cc0003c50d0cc01437440010341000003001300400fcc10300440c400000c40d000f01c0f1d3c400c3013034100c0401300004c10d001c10070000000c00000c0c17f13c13034d1010000d401430cc000000cd00c0040c00c0300c10030d410000043c0d0c30104051000000031c0300dc04ccc00050000131030c40f01310110003000031101d03074dc7070c0001d0000dc13313c5000cc00004000400000007c50c00003000710c0c4315d31000104007030330104104000310010375010c11310c43001300034c030335003004cf01003700d040407110f00000cc010053005400000700004711030100074040070000330510030c00150cd00c04c0407f0f000000005d0c0430c0040314003031343c0470030c40dc0313c0500d401ff0c411730030310030f1d3c10000130f13c7000031000010300003000030d10c0cd34c003100000c04c1053c04144c0f07500033005030f01401fc330000013c50010c000100301f0103c1410105f400003c030401c00fc1013d007040143fc307571001d0c04040003734033004c0300f30040007c5c500440004dcc00c013c0010c04f0c0013cc0001cc3df01f4000013000cc007407031140000313cd011011035303070110300013f0004001c10cfdd0c0340104400400d3c30000c00040040304100301407003100c00d00c00030403d0300c00001001cd1c00d04d44030000300001040fc3000033cc40000004003f337d0c1c00014d000d01f000031001000f00304400d0010110000001007d0107c0c0cfc04cc330000010c4400310011407030cc0400c01001dc4300c0c0007c000c003400c401f30100000033c0d5001c0c00c0030717130100031cd000d00;
rom_uints[695] = 8192'h1cc4040000000001340044540c3c1cf00000040cc0cc70001c1000d00c00c40040773f7c0c000034d03f3c00300004003400043cd00031c1000010304000000f04300c00310000300070100400dc00130c5cc0c30340f0c1c03c700004c0570c101300500030104c305000303040100400005000c71c3403704073003403005070340cc00400001030101c43304000140040000034f044005c4c0c0440140004300010540700100ccc10103c300c0c000c51cc003c010003430000151c00000c0c0c0000403c01101004c000cc0c7000404d3040305f5cc0740001000404314005000004c01c04001c0077c330003017441c04f047000004040000004000c43040700000c00014013c0c0c004004fc000cd00c33c4000004c000403f10cc10000003000c000007700000004c0ccc4c0030c310403400003c000c40300c0100c000cc0c004010000c000c3c000c3c00070cc4001c440c30c3001400d0c3003030d33c1034c01c0000c4104c574cfc0c0c00040000003c003c4c5050c0100014f0144303c4040c00041c50004c0cdc00000000cc000400403c14c000cc001004444013d1c00c00d4004c00010c34100c00010dd41c300c4414400440041dd30d40f030000c0330c033dc1104400c0c001004000cf0401c000010100c40000ccc000c30050c4001070400131c00000040c01f3f1c0040003010340000000401dcf0040f3cc30c101050f01c05030000004fd414c010000cd00c00140410005c00c000100cc0340014c00013404c4c440c00440ccc100170000c00d404100000d03407300003f00041d010cc140c40300400c040303000000000c4000ccf1c1000c10040c44000000000007c50300010303700c03c0003000c01c54c00100c1400500330000003001000c00430000443000c3c070034040014001c0000000040cc0c0c50c0c03330040704401c013c04004c400cc40c00c04c3040cc04d000000000000c0000000030040c0004d0c00cc40000d0c10400035403103c1f04f0cc0003000c030c5cd3000000cc00c35430f41cc0304d703c10000010c04040000300001444334cc04044cc1000cc00300000f00c100c440c3c0400c1141c410000001c0304c004113004c000007c0000000cc000543003001004d0c0cc30005000040337f00004cc344034070cc0000030034c40c07003c43034001700040c00c400001c04000401000007004c0f07000000d000000c004cc040c4040c0004013010c00040cc03004011d430ccc07c1c3474001004f010f40000c0300000043f000010c7d034dccc00000010301743c03010cc0c00004300c01c0ff0c000c030001000304c0000c4007040000100c43000004c40140c1c4000450300030440c4c00c0430c00c0000303000504040001013c00c3000004c0c00ccd030004c000c0000;
rom_uints[696] = 8192'h404d03040140500cc00000c3005cc0c400f50030700014040c03c10041f110505000001d544c10000040c00000cc500370f0730330750001c40f144030004004014553400400c010130010315700cc001003f151f0004533001cc000000404100041cdd01400100000c0f300d003073d4300404c50515000000371007000cd0040004c10140d0054341000730cc043c3031100c0000140cc000130003044301cd55c011000140c05700330f00cc0f07c00f0030000f00f40d0100100430403c300cc010c31000070cc03001300141070050c170071014c05d000f00c0c33140030033030c01300c00cc000f3405440f3c31030f007c04000440010004c1001101c1010c3c4dc00c40c30004303dfc0304f33004153d44000c04543c00f50c3f1c000f000c1014c0c1001c031001ccd4003d4c03c4130c000f3c0070035344c033440c40c0f0c010050c001030d040cc01305c04c550104f030300100300000c00030300077f4303350000dc10104033c005c001403404c00005c054104034533454053c000c74504cc10004cc40000d0c700c7c004000030c4d00050c001d0030051f03410014fc051dc3110030c3503000040030c344407c40043f105c0103dd04000030c30070cd1010103310003c3c3c70030034c4df1003300100004c103500040100040c04033d0c013043050014003ff350c0cccc00103070403c4c040d0f03003c31c054500c731cf400010c0cc00c00cc101103411c40700f40c5773c40000c0c0001000034c043005000111305f0c0040c44c0000c4c0c3f00003300003c4c03c00d00d04f0f037fc0c40c7434cc3c0c000c003c0c10f0070040d0f10d3000050401d1441101055f3c040d4300f0110c10c04f0cfc04003004003c0c03d00010501310047c30304500340110000043c00f4003700c004040300c034030c404000d04f3400c44073cc04c00f00c0f4c00c415010cc40f40417d000010130307c3000000c0000ccf0004c301400347000133c00401c4df0c0537c000f0c00c0c4000d005700c4343c40f0c0f44100c500c340cc1cc34c500140433040c4c0030004010c003010d00c07c000304313330d04c000c00070c000c4400101c00000c00034004cf40000c3304004c050c0f03c1f430c140f31d040c40003c0ccc0c0030000050407000cffcd00c04030c41dfc51fc0310004101104030f01dc0400034c5c10cccc0f001c4340003c04440d040410c04c000f51000c7c0700c3f0754f7fd0000405fc0003300c0d4d4d000c05310d000004000f0c470f3c03050003cd47440041340410000c3030054303ccc0f33004040c010f0000000c1303c0d0dc1f45c1354c1c0704cc430c0410403000301010041c4f4fd014110cc05c300050110f0000010c3d0c301040d131c00405403330c4c10001001f3040c00;
rom_uints[697] = 8192'h1410000045c04300f13410041344740333c100007c001c03044404004f0c0c00013443031704001fd0df3d31c00004d3c400003c3050000fcf0314011300030000d50005cc40310013000d410f701df30c010c50074000c0041c743c31400c330031450103000c074007d13400cc4c5430c3303530d3c03401033040100705c0fd0c14001c0c10c030040cd00c0044000343c03100130c41005fc03000d133c00cc30f000cfcf03144307040150d0c4400141c400000030ffcc0010f1cc10c4743f11000f0004471341c0044cc00f00010c4c500c300401d43d3410f01101070fd310030f1000c0cc33730cc1f550c070144cf0340d1003000000007400001c155c1000c310df00dc03cc03000100f130fdf434400cf45003300040cc0570cc00000c400cf4300c00310cc3000001c1c000f00cc173c04000370103004003403d04540ccc0f01000c30c733c740c000c00140f010403cc05c43c003100c301301010073cc0331d304cc0dc1545054fc0dcc1400070f344307df4010110cc30005001c433d33000100c1030004c41ff4501c33c5014c0f000300100004400010403530d0033343044103c000014450f1c4110c0f07130007777d1f040df0c03010100001c71033113111101ccc3000103700c50c1000c5750000cc00001c040cc01cc40fd0c004010300301df0d01145030c0cc1300cc400001000000334c00d5100c0c0013011533fcdfc0c4003c014101c00403d010040703cfc0cc5d00c0100c10c00ccfc000c3001010051700c43003d40103040000000100ff0cc100cd74df034003c0000f0010fc100000c0c404df007001440cc1f450143044c00f00341d5f0000010c01fcf44444c0dc04704cd3311740f74c3040f010f10301347010d14031440141cc0d0337c7101300c00cfddcc0c3303400300c303c30110f3f330f0c0f040130c34f07c540df70c04073000005300030c0dcc3d01511c04300003f441c04c40003d543000070c005310f3c3400431413dc1455100101100044043000071c100c03330c00f0004013000c41400c303f44331004fdd001d74370037401c1c13300c3100d00c00c0c4ff0031c31035071133101030d00410dc4c300dd0d03fcc30000d30033404c0004305000c1d37100fc7030107415d000103033f03f1030cc00c1030f30fc007710300070d0cc41cd10000000304301331cc70d00f03f00100d00fd040c00004c00f300000d300004343f0dcc370030040d15003000cf0040003dd30304333f7000001d700403130f371c00041033304fc34070070d030003d443cd7010413c350c3c010070c013c0013d0303354c00c340f100004400f030cdc7d01101d3fd30cf303150c011dc100f00ff00740c74f301050c3c30000140303137110c000d0030314c4430000010c3cc5f00140cc100131010;
rom_uints[698] = 8192'h300c030010140c0f43301c0c000f330005033cff00334ff0c00033cc0003f100000dc344304cf305f3d54031103c000433c7c033340d0c303003cc04040001d105000c4c03000001000070341000000010034d14753130013500ccc00350d7cc00c70c4000f00041000004cc0000f1014100300370004000501010013f030030010040000c005300303040cc34010001700000c0001300000cff00070f3100cf10004504c003000303401033c50c0fc110000037c0000030c1010014000d0f00000300d300100d0fc14f1000f10c3c0050000433fdc0c100c1f1c0d0144c0313f000c40400c3f00c13ccd1001c0534c1011033014450430001c31f00510c40031045150303304003000100c0403433000001cdcc0353cc0cc0cff00c04405c0300f00100534530c0ccc10007f10dd0143400f45000430401f1d300111700000c0f37000000c0030f30041040330f3300073010003005c00040100500104c0300000d530030c073f300c7430d04030000074000005c00137300c074f13310530c000104c5300f053000c130300100f030c0300151011437070001fd0d30710c430300000033000c030c00ccc0cf0030f03034410d03c10030034404cff010031c040c303030130c1005f0000504c03100040d0c0cfc001401000333f404000307f0f40c0030070000c3c13f50001144071035103c0333111401440331f300000071453040c00030300000140700f300300100040130003c33000100cd00c7d04030030c040000005c0cc0005140033d0130003331003d31111f04110c040001fc53c1010c0001000c310f0700c001301111cc3410500cf0c0cc300034310151c70cc440400330000330c4101010d070cd001033000c001007c03c01000c01f7000030004443440d0304fc0c300100c004c00dff003001c04000030001034c3401d000404c10c0cfc1070c174173373cc30c0130c0331000cf10c00d033c0d3f370100000030cc010300000c700c00d304343cf0c0fdd301033003cf04330c00031110c4000100000c14131c703cc0001d0d03c07100c0340c030f500c00070000c1cc0100000f03400100140ccf3f010030000070c3ccf4003c0f0cc30100cc003133d301c01c0f55300f400530004001dc000440f03010304c0cd051400050100c051040000c010007d000500f000d5cc70011001034c00d4000c00c0050c0cdd3cc330337000400403c010f101040003103c7004101030004000fff3f44000000300000f47350c434000c1c4df330100cf04d330000f1d70cf110000001001050400400430000003cc00000c00005541ccf00cc1000003500003c4c03c351c0013071f34100400144500300000130010cc03000c03500c000c00304403400040043cc135c00500cc001cf0300c050000003003030c007110ccf050004;
rom_uints[699] = 8192'hc40dc0003f100001c403c5d0fc0031003d0cc11c0c70c10007444030100c00001c700001c3c30400c4c711310100c00770c001d5c00fc0c34c014c3f3001400c0374010c10c4c1150000170c3340330000330304fcc3030f4cc0440fc04040340405c4340c5507c010c1c301001431c743404005c40c0c04305703143404000c00c035030043000100000041010430400f040004003c4003010740510c0cc3c30c4040c00013c0304340c0010057000400fc3c00001d301400033003574c0000003503000100340401000004c3133c303031331700000043cc30140ff4040c1017010000dc574310104100d70c011cd013014c0001c000c000004030f015000c0100c034d0d05cf53c000c0f4410334003050100037300c4cc4c040cd5f310d4070fc0003d0cc51cd0000730010fcf034c3c000340cf000003c7037003074c104c0c04fcc43534c343300c4c0001c303c0c0030070044047000013034c4f0750030f417fc5c001435c30c0050100400d00034500000f001000c51304400c4fc141117f0c4d0140000134001043c0ff04d00c0cd00000c7007700000057004300171cc300004030c3c01dcff0c1d43000f010444700300c134004410003003c0704130130f03f00f40403040ffd00dcf40003004c4074cc4dc0d40300c0c3130003c5c4c00c3004403104470c001513030f00f40ff00540010034000c0547cfc104030f00140c04000003130431140440f15f3443000004000143354143c0100c30c3c443c3c4c30d00001041070000130431c00030003c03c0005c13040105043c0400d00c031cf03c150c3ff3cc10000c30d7d051401050400100000011734c4050001045100c130004d47f03100c041f3c7c0c0c400c13050001301340c0c01034d1d710d0141400c74303f7d00000cf4f430004000c10000c4000c4cc47300043cc33010c005f0c4144cf301d0f003300c3f0000d0303000ccfc51f430c0744c0c00300003000030fc0c00d010f30044d007040fc0c04c0000c04c35040030f00dc03dd01007dc0140f011105407c0400030700000301c01100d44110cf40010030050c400c3f010cd040000140f0000c40400c11d0f0040c4430004103c00cc4000cc4100031c0c4c400000004000c410f010d0100013d0d3440104c04000cd01330000330031004300317011cc0c04c10c400d404500c33300103314d0000010005c1cd00c0c0401043c30c40c040c11004003530000fcf0000c045354c7d30054c0700100c40074c470303300f00c0d00c034000040001c340430440c043030c03ccd040c00033103fc4dcc0fc00c3441435057c0000c040003c000c0d0014cd3110c00cf40014d001cd0414040c040045000300f004f00c030431cf0ff4d00303d001d000030703040cfc00c03014c3cf104cc033030004c30c331000;
rom_uints[700] = 8192'h740473003105030fc70100000d0c4000c0000400450040401033c1000c0d054c001300044011000001f0000440004100c00000ff7f013400140411300c440c403c00040000040344f00000cc010401105003000030033dc40030170c711013300cf57f714004dd0003c3570003c005300100001431d1c3c0c30c0134c04140017547000001c00004033c400430000ff10401d040004c0c000341014c4003034000010f0f3c00330000040f4300300dc3001f5410000001fc1047100000073c30c00011fc350030c0d3300000c0000000001c744040004010410d03103f334c4c03f400004700404f3107330000f100ccc301130077440000300304534c00c1dc01c04307c3f013430cc0000c0cf00dc33cd0003d0011100040140045cc31ff4301c000001410c0f01c4c004050000400c703007c0c40c000cd003030c13cc000403cc0cc03374000070c00f0007fc101405d0fddd4c1041c1c00c003040c3007c0ffc000410fcf3d3c1c00034300dcc470c007014c00040c000400300003cd03d4003d13004c0d1037031c01140000410c00474c0004000004100cf0c05001c54cc4001c4040c1f31c040f000003cc0c0000d1f000d31140c4c07403c0c00d14500f00f3444c04f000d0100c0c10030c030400c0c4d00cc40003000f000001ccc0c44ccf000100f0074c014043d00000f40c0c10c031c40c035040000c011047301000000430005100500d00703030013004100017000140401c0404c00f40c43000f4c10c000014000c0f0310c01c0030350c003000c1f1104443000300000033001010003000003cc00374303c30000f30c014051d00001000001c000c35f3310c0000f40c003c00701000000c11501f3010050c4d31400000030300074f0350f10034cc00004000c044c37c007333ff5c3c1c0000013c10c40000054000c5c3414c400400cc0c40401cf0fc04f00141f000cc03443cf0000f034540c004440100400c000007000f000c0000300c000310d4103000030000c01c0cc0c0300030007c10430433c44070c000d0034fd001c004d00c0100c04030c1004c703c30000344330000001cc00000f050d0300050c3000d3c040330404c0000004001033dc300d030403001003100c04013f001c10c1c1337d04050cc0d00c11300c010dc031114d000710d0000c100300300011c0303f130400030d00c0300004c000100c0400004c30c34000000d00010c0c4c500c0350100f013fc0400000303fdc0304044000000030cf10030400010d0100040c0000fc40c0340cc00100c0f00c0c0004c04fc70c1d3000c03cc40403040c031000c370014030cc3c0000040131000c01cd710345c0500000335c34303303440300f11010d0d040000741cc403cf313f40530c040004f03014cfc300d004f0340ccf00004070cccd0100d004f000;
rom_uints[701] = 8192'h410703c0100cc044c000d01c0c003301cc0d0410040004d03c04000c0000c51004cdd410c10170303c0c00057c04071cccc000000dc10104cc4f40c4330cc43400c0c4d00cc0c00c3004330fc0030c4000430c500003d5cc03705301034004d3c450c4c0000c0000d01000077300000404d10000044000070cf0c000433d0017104c33dc010c000c04c0c000dc3c11304c000f070737000700170014000c0144400031000700cc000c353c300d00430cdc000000d04df1dc0444054ccc01401010031000c404c0040400c03c30310040d100d0f0000ccc0c0c00114000c704004c30404c0c000f50037d40dc3f0d0440004f11410cc0d0000300040c4100057510317f040c300c40c4d050000f3ccc040fc00107100333c703c0500cc0cf00c00007c000100d03000411c0f040c400030cc0f00ccc003f40c0c0cf07003000417401030fc1004000c100000dd40130c70115c404143c010574c4c10040c0030404007c1ccf4000030d070c0d4fd00c015300100303030fdcc30010cd03010c07c0374c01c00f040003c53c0c30400000d000010ccf0033c050340d3c00000003300147000c01003300400cf07004000d0044d0014001140000cc00030040c0445d0340d033000770c00cc00d0f0d03700000544c00310c100c30000030c0c700cc0cc3700000c0c000cc010c40311c000d1c00000f01047110c01fcc0f140d30d40c4440c007400005540fcc433cc0cf0341c00d4003c100117cfc3d1c030414cc40134f010000003f1c03050c000473000c03430000031f3330700711cd030d4c03404d005007df0cd01001c340001040074c013004430304405001cc145000cc000000007100c3f00fc430403c40d4c4343f4cc035073d130001d0c301400000000c0fc040d40c1033f01040030c0173cc07001c0003c74c03fc010c4c0040041011c0cc0c0574c0104cc01d00d40303c101000cc10c015300c10c4c34cc0c03c00000c3030c000000010047c004000104400d0443c4000c3c050f134c000301000f0001c03000c00400441573010305400d00d00400d100407c0070001474405d073007107000ccc30c0044c7010000000000354000f000047110101c3c00000f0f0f400304104cc104710340073100f307c3070f0300c0000ccc4000c33f050000014103c0031300c57100000cc000000c400f4103c3c00d0c44c0000ccc015173c000f00007c00f31070c010fd50c11c30dcc0d4dc000000f1044c33374c00f00040c001103c04c03740ccd00003500c503400cdc0f00033d40444c030001c0c0cc0403f0400035300034000fccc143340c00000004400dc030f4000430c0dccc1cc3c0005d03130040030ccf07f0400741114133df04040410034c003c0047d0c0c0c44c00d4401041c00c4d0c000c000c01733470300400000c0;
rom_uints[702] = 8192'hc0044c00c7c311c41c000310c41c00f04034cc0c0043300ccc31010c4c00501003c0c70401454c1450c03100d0df73c4300c0043cc01f070300000003c7c15504104000440c7040000c10c403000300c034c71131d103c00050c740c040c053100f4c04f1dc0c01c00f0300100c0001000000000301cc00000040047000c10c43cc00003000c000000003c10003c03305005000300704040000700740300c07c1000dc4001fc10c000c3051f40030000373000040031003c100dcf000c3cc344f34c003014cf0cd0004050334d403cc40300001c351400013ccc30c0000411030403400d00110c113030301440034c40cd4fc004300130050043400000030710c0170f111c50c0c000c1411cc0f0c0734d44153c431000fc40c330433141c00c30d0010c000543f030f500c0010cf01c03030034004010000304c00c0cc04c0c1ccc1070c00010010c1f0cd0001007041f001cd0000030f0dc5d0301f7311c4c13313cf00c40001000c0c7d00031000001f30003c013000dd400c400304c0c1cc74c000c300141c000105c34c03040c0040100004cc004770c4003004040047f004317c7d00c34dc0000c00c0d4440ccc31d30000403cc0c40c0404c0105c401110c4330c30001d003c00004c4c00d13741330c0370f40c1300cc0c0304110c10000400c3070c03404f40c10331511d13c4344c400c14f504000033f4043f7000c4c000fc0100cc03511040cfc0c000c104057c5d05c040c3c1004010c103d0c4c000501cc00000c040404dc03040000c0f000ccc5071cf00c0400000fc0500c0000d000c05400ccdcf530c70000c000c040131030045347dc0f10000040f03d70c14ddcd000700004dc004000c0304437530c0030c31103150000051c3d04c150c000c00141c0300c500c3001300c03f000307f4ccdd03000c003113300c07000140c00030f400c5ccc00004034f130c07c34c00c4750404003300050130c000134c0c001f0400440c00033c0cc7d00033403c001430000430d004f1f37003000404310001f440045551414c03003100c1c00035c3c000cc114c0c00300070004fc0f0c1003f000c004433c301fd040c00c004030331040100000cc4001734f4004414c400c0001003c4c4c00010c30dc0c100c0100007c10301040c000017330000050001c004c1d3d04dc000cc000404d07440400d101c03000400334d04c0cd44003400cc0dc01103000003c4040cc0330140000710cf00401c00cd30500c30300100c0c0044010100000c10c0fc130c4c010cc03000cc004c44300cc1c00410c3300c10700d0c1c01100013c0053040c1f00040400000300f47f003cc00300000c0f0c70140c073c0c00014c703cf40000c300c35543d34300000033cc430c04c000000001cf45000c0f3f00000004014000400f440134c030400010;
rom_uints[703] = 8192'h100300001003c43050300300f4004300000004030000c000003410000033430300d0cc110f3300001100010100c0d01317100411c00340430050001010000100001330c00000c0c40000403fdc00c504150010c34c0100045033450000c10110000703d00000050f134d41003140401433000f513c3110030070005c4303c11141cd0f0c11700030000010130040003007c30000003c003414000040dc30c33030133c040001000003003004004c10300074f704004c04d300cc4100440c030003040003130033053040f0004030c43000000000c3d30c0130000131d113000c014d00000d0c4f00cc104000df040043004400350331c0130000403f5014010f00000070c47100c3c00130301001011fd30733d00cc03370043f134014c0000700433300000000033003304000010010003c00d0cc000000c000031300d000c3c0013500051014301004330100000040fc1ccc0007f3100310c44104010cc00f050033f07cfc0c003c10033030c1c153f00c4c04030c00303c010000000410101000c33013000000033100000400043300000d1f00004500cf00001033340c0043dcf0000000c070000003c71001c303c05301d70040004430004f300005cf350c00400cc10301d341047000df0003d073005c030000c30010c00301310301000000c0d11010f40fc01330d030010104401400003f43343005103000c7100503c0010c1303311303010c0010c001c000031c1010030110033000c003003305d030c0331530404000000cd440000030010c0f05001003300000000000300453dcc0d303030c4c700400000000c0000003c0c1300100c000041007f003f70f0450d4030030403c0410031300401c3010015034103330041000fc00cc040c00000301001000310000010c0300001c000303f0010f030000c03103c054000430cc0141dd0f30030077f01000c31034cd014f0533c70c03300c104f003017c10000001033d1f0000000040c704001011f44000000d00f10f00f0fd4037cd010c0371f0100341c3c03f0c0000c134000003031340000cc03300033c0f10040300f010004000010110fcf1c00c0413000340030ccc0c03cc30041044ccc00c0c0000f00c00000c5130004c44cc3c1ccc1044030011104710335330400f0400f03c305c0005030f1c000031000100004731fd033010300c1d0407f0004030f030500c04f30013c0c00070000300103100d000307c4003010300150510041000000d3510043d0c0330100c013c40400007d30300c00d1000cc03fff0030010000cf4000010c5c007134f0d04100000d0d000001c301c110031c00100300011000000040404004000c3014401c014330003c5f013504d03303300d043010f1501000130310d540c034330035700c47000004d144c00d0300300c0310c01f730000044c0001;
rom_uints[704] = 8192'hc1004c11004474c00000400000000500c00031d033000003001f033cc400000040c044400000c010000f40001c004c0500003cc303d43040001440300d0001400df30134400000000c014f4004c045003000c300130000f07140000310710c05c00400000f0000c0c000c0f4c1f070010400000500ccc104400d004cc11003c0c100c00000007300300100c00000100f1005000300101310cc000000cc01010343c47010c5c003004303c0400004000070c040000001f001f00000130300000500035000041030403004430cd0fc00d1f3cc71000000040010003f03300000cf4000000c0000c005303cc000000cc0dc031040054000003003037001c000c34141400f0fc04030c04000f0003c301411130000000d0000300c030003dfc4c30043100007fc100003400570300300033300c330003030001000310000f00d01c00000000400c00000c340cc000400110310cc0710c1050030c0d0000005704041c1d40c000033d001040034d303414014014043c0d040f004443040c00cd000007f5000001300444000c000000500300344c000000304c144c400003343000c00d1014d0000004003c4104c000f0c0314400000533030c04000ccc00000003c743300c0d0c10400c0c040044104f004300cc000010000d0303033c000000310000000700c0045714001331031f30000c03000000043c3040f03105403050c340000d40000000300000030753f4000c5c0c04000c00000c0000301534414d3400330c000c00030000c017c10000cf00c01504000c303c30040000004400040040500003fd0d0410fcf03001000ccd4030740731c30cccc0031337005400510d0c340003ccc05000000400000c0c44000000300c0000c0040007c00411f4004f00f0c30000000c1c00010304174434000347d00401000430004100000d307000314cdc30000c010c140003043740c03331300c0004cc400fc03310f04000040001370030000030000c130100301434c40701000000f0f00103000d3c030030c54000300f0004470004c0430f0304400000040110300170100040d0000c3c000c4300100ccc003010cc1c000000ff0401c030f0000c350010041330040330c0500c33c0003c0104000c14040500d0010034cc0f00f430f004303000cd04c007c43c0004040c0001004001000d000300010c0c50f000040c0c00400000f41f0000f331500c000f404c0c0417000c00c00034041435035053144c000003330f303d5300cf310030000c010003cc0007c43c3c0701470ccc0c054004f400cc0d0000ccc337f04003000300330003c40001100004c4f3400014040f000000043c0030041313c00000fc0c001c00404c00000d40500d0410701003004000303050031c044400003000103d0c0c011c50fc5c00c0c0c3000d004100c00100cd410c0c30;
rom_uints[705] = 8192'h1000040004000010000003030070005000000c030051000001c0f00434000100c3c0551c0004000c7d00000c000c04040000300050300040000000000c300010103340d0c0000000004030301044fc050c0003100d0c3000005400000c0004000f15d1c000000034c05c0fc00011c1030000004cf40c4000044400440000005c0000300f00004003400003c01040403010041000300000030404040503f000000cc001000f0030c00004000c004000000c0c00000103040100540300000c0000d010040000144000001dccd104043340c00000003051c000cc3c00d000cc40117000003c3c000c30d0000400df304000c030073c1103000c4c0cf0000000000d0405000c7c001000000c0350c030000c40000c00c014c0003c0040444d0300004c03000c00000440000010cc00d000000000300030c00070400c100f0c0030c000c404000740000d0101c00c00000000000000004000c5cc01c4cf00001010005034003000c00c4000001004c1f01c000340440000030c00041001cd30030004000040f404c0000d000400000c00c00c00c40c0000c00000000c3c403c4003c0000c170000030434300400004000040d300700300000300447300000000000c111c030010140cc004c5000dd000c050400014c00011c0c00fc010041300c0003000c300c000c010c0d30000c0d0c10430000030000000c03c0330034fc041c31100c14f000040004f000000c3c4300000000004c00003000303444f00003044000000000040035400040003004040c0343c00000403c0c003000010c0004cf013034300000c11000340104100c0305000c4000310003f3000c014400010000d03040403c0010c0333c4400001c0000f0000440004c0c0400103004f0000300070000c030000110005001000400000d300c00000031300c000c0000400030030c0c440c00000001c030c00c00037c4030ccc00030c0104034301c000300000007000030c0001000c000005310100134000310000c04300010d00c00303c0c4d0000000404701c30000c0c001100000401c30334001400c0c000034000011000010c00100c1000130110d013003000033c00c000301010040010cc05040033000c0030007033000000050000004400000c04cc007c4700340c00013004010c40000040343303000c00000c40c0040000c00010300130300c00004030000c370001004000cc000043101000003c000140030340000000403004c000000001010c00010034010000003000100c307040300c34040004d03f0000003000700c104000000cc05c000411401c3330000040000040300404000310000000004040100010000007030000100000c004001000004c00000000c030000c0100300c00c0000500000000001043c00c0000c00c1000050000004c0cc01033343c3030003000;
rom_uints[706] = 8192'h4000000004c00704c310c0713d00c305000040005070100300c70400340004100f4cf00c3c0300005140000000044003c0c403014013004f00001310d44f00c03c40cc0c301100001000010714003dc03c00c3033cc100cc0033cd040003000000003013030110f004303fc070431404103100401f04000004cc343300c0303317ccc100d00700000000000c10004cd0d00015000040d0000305074054d3c4c5c040cd0004010fc0030000007c433c7300c00c00000004044400c0434400070c000dc004f050c0000300141040414c000701004c40c0d10140047c0c3c70100043c4c00041c000c007c1014300410c000054000100010c001c000430400000f00001030040000434301c001001c004d0000cc00340440544f04000d310c30fc34030c0000137041001000cc000c410004000300000000f0000f3040340000000ddf301043cfc03000304304003133cd0c0701003000330c00c00703013fc00000030cfc511033310d7cfc004ff01c1000004c000401010c003dc40c4100000300c001c400003100070430000040300cc4300004300000100040300d4374410cc01c10000c03000f0000100100c40400040000d40c47305001100d0005003413034001c33f503400c0c070f0070000300444403304dc1043d003004000d0400dc00150003400401000c03c010104f00c01c035301c34040030c400400003400000c00c0c0003c0010c10100000103040d00000000033c3c0050030c3000100140c0000f011004001000f0030fc3000003f4c40401303300000c0514437000d40cd0040100c31000001dd4000c005301001cc0000d30004f0c0000c030c140040c4c01370c0f00001001034003c340c001470c4d00000014003c141000c00000004130001003301003150010000000335c50ccd5004010110000c00330003010dcd3c0c010c10d0c40cc450700000101c340001000c040c30c0f40443f007000400000010000000300000c007000004345000cc000c30100c03000cf334040c0307100100000c3001c000503d0001000710031dc000000000010f0c03011047000734034000d0fc000110c040f0000000d170d40c3400000000000000d0100c00f0c50047c044c1000040101c1400000000000dc110f1d0000f30000cd44c4c4000300c04543005504104001c100d10f000dc00030137d10c0c113d40000074c107d00c0cf01400040700c0000f400055000c030c004004c01000000404400037003c413d0004010044000c07100c3140014310053c000040004c10044c30300c0c14400410c00004300044030710100d300730cc0330031f0044c30000100030350c003d13400c30f00404cd10c0000030300c30c0400400000410000c3040000040300c0140140000101000000707340030030d7100043c0031410401fd0cc30;
rom_uints[707] = 8192'h405000000c40301300cc30047000030d100c4000301000000cc003004010100c000c0c4010c00300001000470c00c00000001f3030001000000300411000c0000000c14000000f400000f340000004000010013040c0c400100040d00c04100004010013104cc0500033c0000000000000001f030000c0100004000c0c010043100030c00000000000000001000030010000000000000c00cc00010300c03cc300100040000430000000000000400000c403000001100000c0000134c000004340300c007001000040401030003c04000033400010f00010001000000540003c0000300000000000400041301ff3000010404144114000000001c003c0000100300c0040c0103047c00000013003005300100410c410400000000305031144001000700000100400003300004000c40000000003000d00000004000f0310000040003004c0403000d00041d0001010301300000c00c000000300f000c040d00100cf300c0000c000ccc0305000c0000004c0f01000000100c040c000c0c4c0430000500c10434000d0004004c3001000000000300000000000000000404040c033500030301400000c0040000040cc33500475c300001c0040000000c0f01040141040c1d00000cc00300000d001010030000010000100000003304000000000c0c333000004c010c714330000d10000040400f0c000000334c0000400000340000000000dc0000c4300050370000100400400771000100010000343104010100c0000f01000030000000000010100c03005000001c4d000045c4031000070c0100000004000004000f0000000c00000d004c00030030005034040503470107f104c0033c0c0d400004040c0cc040300c0074000c100c04130000000f07070400030000000000000000c5000430d33d0c00cf34050c530100030d0c0c04c4000d4c053000c00c3100c01040d30c0100010000000000300c00001c343003033040100c000000300130000c0030001000040c3000000003000401003c00000100000004004300040000000c0f0c0104c00001700004000000340400000010010001000040c0100413400001d00000c0040300100c0c000103303c00011300074003130000000c00c10007000700000010001d4c0300d40000c100010003f0300c040c3303cc00cc0000300500f3470c00000003000144c0cc0c0104000300c00000100c3c0f030003c3000000c0003700030003000004300700c1000000010031c000cc00040000000c00000c00040c000c0cc00c000c3c00010030004c0d0000c00000c10000000c00000400300000030040001000004c000003400030033c0000400c40000cc50c0000c0040140000000000c1000000003000c00030000041c0c00000000000000c054000003010c00430003000c00010000103c010030000c;
rom_uints[708] = 8192'h1000000000010330004000000004c000c000000f000411000001c400c0c0040000c10411013f0000000000030000031030433000403c00cf3004c000f040100c0030400f441044000000d3d00300cc000cc4300c3000f0400f0000c3400c10010000c100c0000300000304000410000000000044c0530400001c00f40030c000034dc0400c430030cc0300000c0000d0003000000004f030c010f00c070000100400400c0d501c130c03c110000c0007044010c000dc4c0004c0000cc300f000c0000031000001000003007c10c03030c00341c0000040104007c70000c0400c00000000000c00000014140ccc104c0000040300cc440000003040cc340400354cd500000030300040074c43fc0c004c0c05000004f001c40c4004000001300c0034c30000c0000c0141300100400c10c70f30300030c4003c00c0c433c70430010c000100fd00001000f00040ccf11c0d000070004c0001340001144000003000000c0c000070000c4040c0c5101350400030010000110030fcc00c50003c000c0004f00000300030c001010f0000c3000004004000040400013000001433004040000d000c10f00000010000c0f0f0004d00c005040140c50053c00003003fc17cc03000f4cc00033030003410ccc0c000000c4000041400430c000030003040c0004c4044000041d01c0000000170040000300003003000f40c00cc00c0c0000c004300f3003003500030107003f000c0000000c030100000c50130000c040c00ccc40403cc1c00047000c03030fc0000000001cc70000000c040130040040000013003000c00040d0004000404010030c000000000000071c000500c3014400000004c0304dc030c30f03014504000400430c0c0004033f00c0005000501d0c13400c0001c0c7040000cd00000c3000c10f0050450c000000700043c00cc04033c000c10003000c004f141101431044c00c000400000330031f0003330044c00000000001000c00404703050c00030403040c040ff07000300c0000cc751400000000dc0004c00c0404c000000c300c030cc3040030043000000c01c000c00004d0000c00034000004300303330540000000000014110413440550400305733000040c0c00001400000131c3d00000c04000c00000c0444d0000404c30003fc0fc44c0040304403047005c000040000404074043003000104c00003000c041c00c40100000000003c044c000070000300c40401004d4c307400000c30104400c40000d30010010000c0fc0cc0c0140c00510004c4000c0c03c000c0000c0c43400040010001c1000000340000001000030cc0c00003f0c00300003504000000f00c00077000c0f704000004030300c01c000000440400000c0c0351400700010100040c000c0445440d300054000c000000040004c0dc00300300040003c;
rom_uints[709] = 8192'h3000c003d0000010c01010d10c001d000004ff0047001001c0001c33470000013740f0f0c000000130001c303001030c000300c0c400000050040404000303f00103001000043100037c000000f03000031c301c00f000c0000010034c00500300140744001004000010400103d000f0d0300030137310017003300010103070030000017000f31c400410440d075340000d00040c04d04f0010104d0f0310003400040400c0500004100000300000100430000004c3d03c1003300000c00030d4001310003c0030003400c300130000511c034300003000013000c103403003f0043000f01000011043430d0005004c710c030c5100403000330130100c00404000300070cd1000703c04dc0003300c00f005103000030300143c040030c0043700000c401c70330000003004c00c0c000470300100c00cc00403031000f30cc0001000d030004400001c00000010010040f0440f1310c704534c00c00414034340c030103003c010dfc004344010001000000430701004000300000c00133d043000303530000c03000310300011300050030001d000040400c40c000cc01000f400c000c50030c00030371300403700d0d0341000440000f011444400df30300303100c00340300001f300c341000710030001d35c000c00004000000300000073033040c000d43003c1130030c00007c0c00000c103c03040003000c01100033300300000000740307030000d41f031003c0f0300000f0c00010701004003030d0301000004004d0301c0003100000003000ccc03044031000000300c4f410104000c00c00434cc0000c01d04000000040003034400030030004130141c430000dc0f03310000c04103c00300c04c0500c0010c343033c033450001d0140d05400000000d4001c010411001030307c043c4000400000003c0403c30000043c00000000307030341030103000c1040010f0003000003013c0004003000440100000000c000d0c40301c300dc000000330031300cc000034440c1f403100d00040334330c0c0000000300040001000040013c000c0005000c300c104400000000300f0d013430010000300000403c0f0130000303010040030045003cc0000300c000003000010d0040c0c040300011440400000014000003dc000c0130303530030000033d00010040100400303001305000030340c03000000c0f1c03301c01171000007101000005310d1d4340ff730f0cccc0c000340000070d00003c307c10000003c3400000000000304344f34403c4003000c0004305f00310004000c31c10000c1011c000040d004030000003317300000c000000000110030704cd0570301c0004310710fc0045000000c04000000c0040000003000f0111000100300014001010004403c40cc0130043003c0000cf0f031104040000000001;
rom_uints[710] = 8192'h7c0c000003040130010000c0030d054d000c0433000f010000400d0c437f0300010cccc01400303000300c0045c0044043000f0301c0140d03000d400000000000170c1c0c00000f00033c7000cc0df0300d03073000000030cc043303300000c3000c010c504300033c030450050d07000cf0131100000040f41f0001d300430310030f44001130000000030d04044400003000000000040003000300141003000700100304d0000c0003fc03000c0010cc0d00400000010001044f001400700f0c040000c5c00f000c0d030c000c003004000c010c005000c010004000000005003300030003003f0033100f004c040001f004300000000444110000000000030401000c4130070c00000000710c14330f0010000c304004004473003000000300000041300c111df000c1000501011110041c00000003000c040d0fc35c04010110c00404000d000007010cf1300010001410d4c011040c0c100c00000041000000010cc17001040013043300430000000000300000000c0010030030000f0c0c0103d01000043000001004010c0301c00030004c0001140c0c004cc43033cf30d000c00010400000d0000c004700000d00c00003c4dd0c3f3040044c0c003300000031f1cc0c040040000104010c30000003001dcc0400150fc014fc0000433d401f44014c0400334001300504100c030d00c1001000070000cf0000400300c0004001101103003c00c001040c3c30057001030d070001000c0000c001101c00034d0000070000cc033000040004dc300000000410cc3400033300303c0c04401c030c043000000000300313000401000c3017031300000100010005d3430000000c03040c30000c000310003000340000000030c000410c001405004c040c0c3c01000c1d410400410c30d50030c10001101000000101000c0c000c0f0c0c000c3003310f1003510c1100001400000f0000031c0c17400044100001100f0c03c001000c000000000d0001403011c00c0400cc0000311003d0003003000000330103000110300404140000000100013cd0000c03000300cc30100c01004003c401730c001103000001000001c010013344443030000cc03f0d0310010c1403000034c00c01001c30c1300133000c0d000c0c1030330001300005c501f107000d1110c3f4013d1000001c00300c0c00030c031d0314300040000140173ffc00440f0fcc00330000010d33004c000000c00c11403c1300030001000f0c003703130c7c000700730c013f0c11410100001c0d101c000c001c050000003000333c354c0c33000000000c0701000c04003c0031c000c11000000100403331400c03000d3d4450c30c000403333c30101c00130000001010f0030300000c0004000004000c30c1071c034000003c0101cc11310310040cdd000014fc4300f300;
rom_uints[711] = 8192'h400010c00500004300400300000010f013000000c100c0003130003000430003430001f030001010001000000043340000400c003000101341000000c03cc10000700000000140010017433c0000c010c0c010340100100c03100010003000010033000000004000c0034030400340c05d0000c00000000040c00001033000330010c05000000000000001d1000001d000000000000000004300000040c041100fc100010013c401700010030030c00030d00000c000c000d0000003f001c01040003003000140030000c000103100000c000303f00710007000c0cf31000300c000030000c010c04c003300430c3000000001105100400000001300d10000c300c0030c00c40c030070004100004131c00033401000c03030000300d00001007030000000000303c10040030000c1430000c1c0003340000030000c010000dc0000400030000330003040c00c00c0cc330000033140103cc0101003c1000000c0000050040110001300000030c043dd4000c0000010014303070000000c000430c4430fc0c10030d00340010c4d5000000000000031c00000000100101000054000d00300c0010003030000c03d3000101011170d000010001000c00000300300003000000000c0000700c30044000c0000c000f0040000001040d001100300001c300013004c0040004043c0000003000003c0c30330c00c00000040404f000000c0400003004011001340cc400c500500413330c0100300c014f4031310c0005041401000c000300101f00100303000404001070374104133000000000000cd50000000001011010040001350000c034c3033004000f00040cf0d01c0410f00300071300300c00073003000c033001043c30301400001c00000c133d10310000d00c03001c000140f305400000300000000300000130003d000444000400340c030430003003c00410c0100400cc3500000d000004000000c0000000000c000114000004310000300c07c003000000403000000700d4c00c0010303c0c04d0000100003cf030010000000010311330c7010330d0000c300d0c05140c0000300c000033040103c0000010000300c4000d0001000c00100003000c0000070fc40001000031000f03100c000000000401010fc03000700401000001303500004c0031c00001000c003c3c00110c00000000033000100003fc0010000004c004003c0f0000000d4403000010c03415310c3d3000000304300310340004000000010000133305000410000004c030344c0d010ccc000ff003001000c0c3030c07040000030100003400000000000000000740004010000000000000040310030040030c30000c3040000003010300000c0000104334000010300000000100c01c5c00000c340c000010100c40dcc13703000300000c000c07015004700000000;
rom_uints[712] = 8192'hc1330c007100070300505004f300330113300000300050000000c000130300000031d30004c30030033000c0311000403c00300000c31050131154c010300400c70f45040cc0c14d310000300030301000c40c00011c00000cd05010c0700300000000073300500000fc510000005000010000013010d014c0473000114710c30070030c0100000000000001c7047511171000c0000000040003004013000010307c74040011003114030000040300000030040000d3301000c70040330c0000000300c033101400000303100000004030c3015037000000100f4014f340030000f00000f000f50c00cc0000400c00401000f010c300000000101444c01000073c0130d0c00040c1c0130300400001c30011100c10100073f00000f3401000d000300000c0c400000300001303001000000010000c300400145300100ccc300040cc00040010010013000010cc00030401c000c00001000310d0d00300000c0d000f0cc0d310c0c30001f0440001140114001030f3d0c0d050c004ccc00000cc307100010c0c0003c0370040400000300000130100400000100d0f0300000030034100000cf00110000033043cc0000000103100040001400d43c00000340c300410003030c00004013f000c000000c40003310003500f7c1010000000030301c0000001003000c031353000104000000000004c00300043740000c0d0000c30c0100f0010031c0000040c01000f300c030000005403004c00003000000050c00c00005004d00400313003003004000003003500401070000000c000f000c43000101050304014300044031000f0000000c0441033300c40000400f0000403d110400000440040000000001c001f100000c001c00c444010001430301010c34001c00301000000500000c30043010100d4c440c0000f30d0003400000003d400c110f001304004d304033000143000c5371000300030004004005070400003003c00f00000003c0110000040c100033c03310f00410001c00300c010013003000000041007003030004010101000004c000300010410000004300c0c1074c00300000000003cd41000c00314000000000c00100000040000011003c0040430000040003001000000c0003c073c00010010011300003400013140003010d104140040000100300340130000000104f000031000411500001300c0d40011000131c4c01010404c005013101010300040003c0340031010404003d00000040c00000300303333003c003003d3c0100003040c0000333010c0001004f000114301400000000010040334000400040c0300c0004410500001300000000000000400001014033f3070730030404000d0c04000003401401010010000004300300c00c0113000304001000f0000000030300000c043000f040030000000003000000300;
rom_uints[713] = 8192'hc000000000000000c0000105000000000c000000c03700000300000300070000044c331d4c00000003100300000003000300017000c30000000000010000c04403c1300030000030000c0000c000000010000003030001003030010040c3000000000150c00000000401010707103000c440010000030003000001001d0003041000000003300000000000003300100300000300000300000c53000003dd310105000000011040c00000c0010330000000005000030004c000030003c0000000030004c0000010000300005301000101000c01010030030003c100c000100303c300000000000000030001c014000130400c3100000000030400010300030110010000000c010340301000051fc30d00005003d00303010c000003041301000040c100030f0070100300000c0c0000000303030c000d0000000000000031010c00000300000c0003000ccff0c307c00013c00000000c00303001c0013040d10000000f004003c440c03300000000701004c100007000000003011034000000000000003c01000340303000000000010300000000000011000c00c000004000041010310000011100004000000d03003331504010000000000004000401030001040000c003030303010101000000100000c301404007000000c10001000100c000010003000004004000371d4340030114c00101000001010c00000d4000c001000000000000c130c14001100c40c003000100033000100000430010c0014000001c40040030000000000311010030000d1000001000040000310103000030041030110303307340010040000040500003000300300001300001000c04000000000000000001000000000000300303000007333100110000000040030101010000c00000000401000010430030010c01000130000030401003000004050c010004030010014000300003000000000010c0000031000000dc00000000100000000000003000000000000001c30000033001010100401303000303000000c3031c3000300000000c00000000000000013003040c00c0003000000c000c000010003013000041000110100300d00030c001000330010043000003300300d003c0000d030000c001100000c0310030000000000c0cf00100000301003000404d00031000000000d000030030c00f10400000c00101005000000403030000000c30000300004001000003c0000040310c000103cd00000041000400400000403000001c015100c000000301000001030000410c0d0301000cf0000000330000000000c003303010003040c4000303300000000401c1100000400000000000030073310003003003410c0000000100001100100100c0000003110030000c0100030000000030070f3000000300011300004073c1030300034000030c10300c0000301;
rom_uints[714] = 8192'h300000001000003100000010530000103f04000000301c10000301000011c100030f000003000010011c01001c03c0100000c03040330003430113000330c510330000000ccc00d410000000054343000031130033310000c0c0001000400c400011400344000010c30503000001001000040c0030c100c100000040000001000053f40303c0003f00030001040300000100000000000f0334010040d100031000c001041400100400000040400000000030100000011c0100000030100c0300003100003000030003000050004c1f1000001700100001030000000030110000300000000c1001030031007100c04000c00143110004000000030000000000003005013035000000300103300400c0000403014000111c01000000301045034c40c00c0043000c00000050c300030f1300003030000340000030170010f030104f300000000003000004300071300300000370c0101400300c003001000c030000000100c0003030cc07c00050000c001c0100000030000010030400000013000430d333000c0000317510001000000003000030001010003333001c03301030051f0c400000003000000000c400350030000004c031000000013c000100d0003300d3000000000330000300330000041000000030c0034f03000f000007040330003c1310000030300d000000300300000034030c0c00000000140440104000400010f003000000001003000004004404340010334000004f10303000000000004c570004300000000003010070f13000c03300005300100300300005000430000500c0000c3100040400003c030000040040003013000000c0300010001305000410000c000310303000000300f00005c0c000114cf3c000031000050040000035300c30000510300000100130400010d0c00003000110304004304c400310c04301d000010cccc000c0030000040300000d0301000000040070d000430003104011030300104000000030000030c00c01330401101003040404010c003c3cc0000c03400030030003cf000003034070c0d010000c00001c000000c030c00033000000030300100400004000f000000f00000030003001c00c003004003000435f00400c07140000f03000000510003000c040001000000003c3100300000044c533130000000033030c334310c000000030313010001000043010100333173100003c0c00000003c1000331000000400003130030300040c000330000004001000700300000100000300000f003000700c004003000031f0030030000003301000000c3000c003000003001040000000c00303130300c0c000000003000040001c03000000107000000030000000000401400000004101300000300014040070010100000303c0d31000000f00c00000000c000100c031004041000001001;
rom_uints[715] = 8192'h30000c0c000000f0000c003000300030000017d01030000030000000147000000c010000000000010000c40000dcf04c000000c03033100000740c00000000c0040c0030400000000d000c40000000001000c01f0000c00005000000007c03040474304000000000c1000040000004100000000c004c0000300010100001404000000030c00000000000040000000c41000c000c03000000700cc040000000c0d004040400c000000000071000c000300040000000000000004c1c1000000034003000300c00000400400c00000cc0000040104c00344043400c01c0d044c000000c0400040000003007dc4100c01c0040003040000010c00000d010000000000c000001040c0000030c00c0000400040000000170000c00000004010000fc44d0f0040c1000000013000000000c0000000c0c001010000400007c000000c000003c00c000c00700330000100030c03f0000c00044037400c0c144000000c0013cc00d400034330004300c104034030403030f0000340030010c303003c004c0c0000c00f0400c00004000000100f0c000701000000c40301c007c000000000f00000cf00c00000000010001c01c00330000000c0000303000000310cf03000710400430500000c000000000003c0070000404c00c4cc000c0100000000c00300000d00d00c03000c4cc00000000f0000701cc007000000010400c00000100c0003044040d00000c44c100000000000070300d4000310000003000400040301d0000403c4c010000001301304c00c00040000000030000c41c000700003000000000c00030c031003000003010000300000000c0010000c4000003001141300300000730400100100000300000000c00300400c4103030001330000000400c4c170000c0000c400000000cc00c1010100010301cd034000000403030003007040c44003000000001104501c000000c4040003000c004000000000c01300000c00c00000000c00c400000000000007c0000300030000d000000c4000410440100040001c000011000c000c40000040004000cc000000000000330004001c001c010000c00000c44000003000003700400000000300000300c4400000000000010c001c00c0000400000c0c0d000300000c000000000001030c00000004030000300c050010010004c0000000000000c04303004000003000f0000c00010000000001700140000c400000040c0004004cc00c30003040104cc00000000003000c0040000000000400000003010004010003c0000030c00000000100c0c30000c04000c0000000c00000c00004000c040cc00dccd30000003000000000010004004c0000c000c7300001c0030140000007000400330003c030cc310001040000010c04000043c0300430040003010000700c0000340c0c000004004100000000;
rom_uints[716] = 8192'h40000000000000005000004100003c03f000104000000000c0000703037f040000000f40300000314c0000003000434004000c30007040000001400c0004100c00d14c0400000000000c00130070000043004000d0007100f4311000c07000005c40004304f330003c10c00003004004c0303c00000c3c100300c343d044401f000c100434004400500001d000c00c00000000000004000c03000c00000000c004f0000c0140300c40000cf030000c00000000000034c00000500035100000001004000400c0030300c00004c01000000010007000001000000000000c0004000000334003010000c000c3c03300040c00f030c00000000300000c330c00010000f00ccf400f0100400000004000d0000400300000000c07cc0c44c037cc0000000000d01c0430c000c010000c400001000043070000000000003040000c300000401444dc33003773004007104430044000307dd040144033c00c10c050000c030c31cc10040004105140040000000000000000c0001c000cd3044300fcd0310044c00c40440003430000c030d03c00005c700c00004000140c1044004c00cc1004c0f000000c0001040000c00300070001300000000f3c0001000000c00000330f00000040000004000040010c0f4cd041000004730100c030000c330ccf01000034000d401000440050000c00001000303cc0700000000000001010ccd0c400300f04010004000c400010cc4000dc1004301c000001440000100410100c004430100c0300c0000050001c000000c03000004000000000000010010003f0440f100000000000300000010051313c4004000000f010c000000c000104340c04c3001010340c030000003f00000000000000400000034000000100c030c00010000c0073040c034400000000c40c31004501101030003c00c00c000000c04000040001c0c0c1000000440d14000110400015c0c0c0005c000000c050000fd0c0100030440000000440330300100cc00000c0c003003000c041000c5c34703c110010f0000000c000c01000004c3000443010fcc000c0001c00304c01000c000000c000c50004014000001c10000001dc00cc0030000c0004001c40dc000400400c00000300003070030cc0040000000030c03000c0000c0500300400010030001001010000000034004030f400000000c00003040c000c0c0000007414143100000c04c0c000f330430c001f00440030000c07000050cc003c00cc0c00000010c00c044740c04c35001330000400cd00000c0000cc100c0300c300c4030000304010040c3044000440000cc0000010003cd0000f0000c000cc10004407000344131000000043000300101000c000c0503000c00000000000c00c0430cc00100030000003c00cc040cc0003c04c0cc00300000404004100000fcc3034c40030;
rom_uints[717] = 8192'h50c3040d10014000f41003070004c005100000403c0c10000500000f03000000000330401d000300c0000000001c004040c000cf1000017100010005c000100d0ff3c0000c033c0000003cc41000c1000330300dc01c0400540000c001f000003055c1040000c0004070300003000040001c344000010400100010000410c110c430c000c33010d01000000400004c1000000010040c00330103400cc10103010c00010003c03d340cc0000040f00f0000003000013c100dc43400cc0f0000001110004400d03130510010010cc03000101070c4000011331f0cc530004003100011000001101000d04044cc0cc00003010334400403300010c0100dc000010004000004000c10400c0d0003001c110103310c00c03d40000401c1f51034000440c00000001c0440005c0000c40100731f0400300c0000c000100103037000000000c10307011000c00cc007000c00300f4101c003031d1100cc40400041440000cc41c7c00c04c0c03d0430051d00304000f010c500300033040d0000c0304410cd71101c0f1401003001010c30001c000301c00000440105303100031100041c4cc0300c000030500cc0034000000dc170c4cd0001100c0000f00c01000331f1005310c1d00000c030300110000030010c304d003c0730000001007010cc00c00fdf33000500c00c010f1430c400033000f010000005c07cc0000ddd03403d0c000c04c00c300c11c00411030004c4d0c0300d00004000000c00004000c1000c040cc4cc30310030cc4407140510c04d04d004c44340c050fcc0304001100000f10043c0c1050005c01000011010400100f30000003004000000000003007011100400c0000400000340f0cc000001d11cc00440c0c34051041000300005000000f014d001003410300c40000401c4f47c1c10c0000030d0440010000100c003d3000000040c0347001010000405145004300100c300c1700700500fc4003c107f400c000040003000030000300040430070013430100ff00011c03c0d0400c0000101d10000010304c040cf400000104c430f3f0c00003040040c00170401103100d0133c0730c00100300310477031010001d100000000000104000cc03071300030130500000003c000000d00100030c00045c40d003001030000700300030cc140030003010f001000c40000c0c03040111040c0c03000c000dcc13d000510c13c000300c000003410d0001d030300310f0000c030330000000c00003151040000100000001000103704c014104040005034303000400c0000dc0000000030c300000001100100000c4003004101c00414100000010000000c1000314000035007000450f000304010340000341100f4100031100cc100004010300001104d0404000000cf300444340410101000110c03c040340000d00041c000401;
rom_uints[718] = 8192'h1c40000300100001010134000c0403007c0110400c03d00000003400300507cc1100041cc1010003300000100c050c04500553040130c40304570500100c00000000000000140010000000300000cc030003c00100f0000000004037000004000040000033000130100700403300f000010003000003030c0004c10030c004c130f01700133400c00003000c00000cc4440000010004440000300100070cf40003310c40003001400033000000103c000304030000340c04040003ccf0040100c130000130000040400000003400300f0003010000030c03000300344105000c000c03000f000000004000f3005300400000003300400000000101400511000143000041030c01000033003710000000103000034003500041c000c400d03010c04000004003400400d330304000f10301304500100c3400c30010140700004300000000005c1c00330440f0001030c4300034000c010000004000030f00340100010000005c00000c30001100c43040000040100103d00001540f0003003c0000000c40000300000c0f00003000004c000007003000d0040000000000c00000140340000000000400010103dc10dc0400040013f10700004000cc00003c400c01300300f0010000003030010d00303700000c0100c47f3c0300000043000070c0000d000000400c400cc000403000000c0300004c3001f0030c300004000041000000003700000c0000403030430000400444400400130044300f00c0003300000704034c0000130000530fcc0c00310013100000041c03000330000400c031330731004001f40005000140003000c04001000004040c0333c00d0740000c0030000c004cc000000c000c3434010030c01000040000130330000c300400c0010000400031000400010c40f300041c04f330f05000f0d000000c00000c0d003300004000010130100300003c04000431c0040000340c030034000100000000301c00530300000c00340000cc40000003100f4040510f0000014005040100040001004000473330000004001003c300000000030300130000030004000330cc014500000c010c00030040c7010034030000c00400300d331000c030000c0030003c33000c01001300031c0c00000003c0000000f003410000000144000440400c00cc140430030030701040c007030300000000c0001f011000030400000031045001c0000000000300404000000040500c03100000017c5030130000100510000c000c0000000c7c000000030000c431050410c3f007004013440003d0000401343cf034c0000003304040300000000000433030dc5000007000c00001c0340300000000013004000300415dc01000000100c1000004000100000100c170434030c0300040300f000010dc30000c00400000000000013c0c3000f00700000000;
rom_uints[719] = 8192'hc31004c01001004000000300c3c45f0c000c0cc040c00000000030040cc0000100c04101f00c000340000cc30033c0070f0c4370000c0c0001140310c00300c1c43000003100005000450000007d440041100043030440407343c00c0100cc0f0f3170c0004004010400014000c30000030c01001003000404c13043c00400c403000f0000010103000041300c530010c003c000000301000030104004c30001330003c0000000030000004100001000000040000044c003c040c30340030001003003c040004101c0000c0000c04300c004010030010003cc014130400000433000c340f000c00cc000c40000c000000300140d40000c5000040343c000000000000c050100300f03004030c040c301d00c00010000047c000301c043cc040c4310000000310000c3c1c00005434100c0c1c0003d0000007c0f0c5f01040500430000c0f0000f0300010cc00d3000c0c0050c04cf4501c1404fc3c0310f0004c010000010c3000104040700000c0000c300c04001c000c030d5cf4001000d00c0100140c0c00c000001440003c4c30000010040035133c0c4c300414003c001d740c105014300000003000000f00d70004404000100c04013000000000001c010000000400c444000c0013003c00c110130c0440f0000003000004f0c030cc04d030c05414033c10303d30140050c5401c003c0000f00c1000040c00040c0400c0300430000403040000000030000c00000440001004f4303400d0d03010001c3434007c3004001c34000c104400303004340c30c00107410c00c40034100c00004400c0cc10c430700100fc000000001004400c00000040400000003cc010100dc4c00400400c010c000c0000000c3001000d00000d3c510c40c30400001014cc0003043c04c10d343000040c00c0040c400070000000f400044003040cd00000f5000000003c30531c44d0140c000701403c3c344c3c003c1031340c000c0030030000000030d0000c000c001000000c3c00053004500400034d0034130000011031000010000010c0510c00c0340040300040c000c1103400044c1500100003014f0040c404000cf00100c004040000003050104000401c17043030cc10050000401000f004f004c01000000f044c001000051410d40c000c3030cc303030004400100c4c000010000000100040300400c7c40400100000000030301c00c00c0c3c000cc400340c040c3004cc0030000c000cc1c00c040000f4040ccc04cc443d00000700d000300000340c404c500c101cd00000f1f05410501c0000c000440300045400f435040c0030000c040700003c040c0004101c0000cc0c004c01000c000c0c000000c430040c0000700c0c4030000041000501041000c400300c000011141000003030041c310034c000c03030300d1300450f0500303030;
rom_uints[720] = 8192'hc0300003040d001050400000000c10c040100043330010101c00c04001c000000000403dd050403340f00001000034340040f0100040c0400000c0000cc03000033110c0011000f0000003170000000c00000d00c003137c004000300041000014010cc410300010000100100040544050000000140000100700c0000010f00003003010013010d010c000f030005034000000000000f04100c000340010000000300000007c304000c000433130004003013300000000101030c43400000000701c0000c10000003003101001f0001040104400000000400000340073001010401000000000000010304101c0c0000104f1030000400000400010000000001030f000007170135c03040103700000000c31000000f00300c400040000f0107040c3d0000403000004100000c00004301010400051701000c0001003700000c000033000040010073000d13c4000000c0c00d0c0000000c0100070000110000003c0004400401c300d00303040c00041337710c070303000033700004003001050c00014cd0c0050413403c0010000d0000301000000000010d41000f0141000d0f0f03100c0c4c00010c4d07c0001000040c330c0001570100430301104137010000013401000000000001110c30017703000034053010000c1303c70f3c01030cdc3000c5c001cf0001043005000000001331c0010401c3cc330000050030110c1000000010000004000504000004000f010000c50005000000350010cc00000004030405000300003c140000000100000001300104010000400000000cc10001000f03000000100100000c003c75041001c001000400c0000c00003030c7f100000c400d103dc00000010d00000411011000030c010000410000030cc00103c70000010100c4000570300000010100000501003c0c040c0010003000010c00000c700c00100014000c34c534c0010414310011000c0000330d4d0407000c00c0040010000000000000030000000f030031010533050001000000003c0000000000003001c000010c000301040000000003300f0000000fc00c0103300404000700000d001d13c300000d0011030304050c0301400000040010000c000c000f030004100004130300030d000c000000c000000574000407000000050004001f0c0d000007030070030000c300c4030c000404100000100003000000114000000c000d03300000c0030000c100040030000c0c0034000f040300000300030004300f00000003000000000000000d00300000c0030004007c031001340000010700cd0000c0000000040300040003000007030d04000c0d00030000010410030000000c0cc04fc00003040c0000000300c1000400100304400100d4010c3000c4031d00000c040f0003000300441130000c01000c0003100040100040000004;
rom_uints[721] = 8192'h310000000040030400004003c0030cc00f3000110d11443100030000334103030400001c0300000000c0000003000c01000000003c0f00c001000000d1000000000c1303030100013c001000010700000010034101300f001000000100013107300100040000000000011c00000c5400000013140300c01500c1055f01070300c30047000101030000000000040300100400000300000d000d070001400c0307000c03000003011dc3c30300001c00300304100300000000c03004014001c000407737000700c001c00004c01000330c3c70d0c005413000013d0d1031000000001400001103100030330001030c001c0140cd0000430000000303000d330004454c71034030000313000004000300030dd303c0c000400407d03301000403c00010c0000001010000c00003c0070100053004331c1c0d000303003000130d00100141000c0310010c01000000000104130c00030c140005330130500003030400330d3000040003040000130d00041303c1000301c4073300041300000c30043c030c0031c30301014001340c01030400003301010001000014000f04000101000f00003300000300030d30014101013314003d00cc00400040c003010100030301000f03c500010105100103001000307300030351c30f010c000f100000c10441330000040400011d000dc00f05300000c0d0000000c30c000100c0c01d00000d0100040303000030000003d000030344c73fc700c000c1c0c1cd0c0c1000010cd700030303c100011f30cf43440300c0c5000fc1c0000000010011000107030400004303014000030000000f03000030050144000fc10147013041010000000c0100c300000301001c07000010000d040cc40d0c333c03c40f004101310340033030cf00001300c7030043010001004400310c00040000040000c0cc31f3cfdd33cc43030500334c37c30301000731c40304000c0000000d3303013c03100c3000c300000000010c000003000c0000133043000cc111733701cf0d0c000000000d033300011f0013c001344c00013000c051310101007c00030011030000c00c070307000340410410c3000404000d00010400000040c0403f0040000030c01000003d1003300031010331410c00000034300130000003000300001005040f4004110c0000010001000000330500030c1303000103c3403d031001030d11010040030c0c00d130101000040003cf03c100c000343d4101cc000300c0300005c3c3cccc00000f00000c043040040004043003340300003100cd0100c003004c000100cc0000100000c1000100000400cf00003100010300000000113c01030003373104c00c1000000d00c003000040000000330300100c01010d0f070103c1000000003330fd0400414107c000010c00000c030130000c41000d00000000;
rom_uints[722] = 8192'h40c30040003000011003004303000000300000311300004c00000c034734470000104103043400c010110030000300030f7d00f03140c3c4c00004103000000000000444003000030300101040000001d0000034400c0000cd0c443400cc00f000030c1107c0304f70c1100000400301041044103044704000334050000c100043100000004c00000040000c0040c0c140000000000003c00013cf007031000000c00300c40003c30010cc0110c4034f00c1c40100f0000100340010000100000cc000000f03330011000051f0c3010043f0001c403c0701330f0c000f1100c03c000000c030000000c004cfc100c300004103100100000010300001c000400073003701400d0000010000c11f0400c400c770004400030fd011403007070000000c4c00c010030c00c10300c0003000003300c007011000000000004c30040004004c3f000003004003000013401000074030040c03c000c5fc30401010001f033f03304540010050f43c30301010c404100000c011100000044000f0c0cf0c100100400100c000000c03500000c0c0010000000000411c03000041000000030000040034000c0c0303734400c0010003c04cc11000050000004103340c440310c0000d0333031c000000c3c0000000430d0000c00440dcf001050003070030033304f51c01c147030434c0c03100001100f4400303000000100000050101c00400000d00100100c0001f01cfc50000f300045040101c00370c3cc300c0000d0034315033340434000031411300300001000d000c070000d000440cc040403d410003000000f011003df001c3004040c0c110000100054104c000000007c3c3d110100003003075cc0003c00c0c010430f0c0040010001301114f030470c300010f4f0070010034003043110503400434d4033010001034000041001f4000030011005d00040c001110010004c00d4013010c0000003000c0000c0333c31c000300c013000000000304000000400cc3530000400f5c40c50310007100000000310000000300c01100070d11000001000f00000004330000131033c03140300000c1000000000c11070000510030000000c03d04000100000001000000400000c1c000003000000000000000000000100003f13343034c00100c340f03030000350c10030300c0003003c3030f003003440400c0301d00714000703043c00000cc000001000c0030c00430003d004000c0000003403411110171004000c000cd0550d030030003000d003000ff001010c7014c000710f00040000000c131044410000100500000cc0331100f0307c0300154c17440000000000c00000003040100c40103103043c50040c040000003001350001000f00000004c0403c074010dc00c010004cf037003100000004331c300400334030000000034c00000000100;
rom_uints[723] = 8192'hc0c300003c0030cdd4d000014d00c4101700000030c3f00000030300f300df00c141cc1301000070030d00104001c0c00f0000700303100c10c0d113d400c0100003c110003400000000105ccc507000100044cd3c47040044001f14000000000c004707100057000040d44004d3010cc4004040000100c000033d4313c1000c0344c330c3370010000300003310410c04cc00000000c040c000010010c0010400cc00c00340c30f010300007003707f404c10000014310c00c010cc0340c040c004000100001400c301000404411f0040f3543000300050c3334040030000010701c040000401000cc7007330030304033c4310dcc540100005010c040000050400311000404103c03070140301cd0000f0340007007f4001070050300c070001000000400c0003400540d0c0004000000000c1c740c00070303003001010c0100c00c000d0040010030d000cc00c0100cc00353f000003d4030f500000000500c37004001001040dc0cc0003700d10310c143003110d00f4d31030000031003f0c001313100000c030000d1d00c00043c000cc004000003100001000404001d077f40300fdc0040040c000c3033f3330d14cc73d00410c4001c40300c003011d0c0f303000010707511000c1c104003040c1344000007000000413433001300000f1013400c11c00cd0010d1c4010113007040000040000cc01013c30c4f43c4004000050000301cc400010407c000c0033130d00d4004040440cc00030c0d00f110000401d00c003014000000000400031003c0030c30c130030000c3030c0f100c400000c17004440410000d00000001010001010340c0cd0c313101010310403100130413d5330000540000c01000000d01000c00cd3001310c03410000104003c4c040c01100100000f0440000100131c3030030000010130030001f300043300341140003c3430030050c000140331c000170030001403001d4000c400030000000000000004134300003043d0000030104c0301731c043530170cc0000000010074000400000c10001cc003030000470304c4704040cc4004041001003000d0d41400014c00014d000c0004044730004cd00540140103303400c000c304000403043000000003301300033310300c04c03000710c17100300500010140c00d013070000d1074330d00c04001f0400044c40c000503f3c70003040000c010c0f5300c000f34c45000410000003107303041040f400300004cc0030300000000c400014130c400c3440010004501010000f05374000f00c030004300c30040c040170c3314c000700c4dc0300000130011f30033c00100300000031000000100730040f0040c004c300010400307030430c01000000140100301000c410010c044c401001330f300cc301c100333c041cc010131434f00f04f030c0000;
rom_uints[724] = 8192'hcc00000cf0300c0110c3c0003000c010f00000141c01100000c000000400000000c30c7017c10001c3400040c0000440fcc00c405001404404000104c050300000ccccc0f0000c0d000100004004700000300c5c00300000010030700cc000cdc03030c0400000c0c400cc004d400000100030001c00400034330c10c0c340c04070c001040004c0040000000043434000100000000401005400007443c303c0c410ccd00040043c000000c100000c44cc003110000100000000c004173040000cc00100c0007000403000100c50cf03030000c040c00040404003c031c0040cc000341040030000003001000f3040c00104400010000000000403010100030c00c1704c10540c03004003c130700001441000700400c000170400010d00001100100004404001000000ccc3000300370010c10c103010c04000c000c0044013c14041cc5c00c0003040044c0007004303c3cc0000c0c4f0104c41000300f03000c000410d0000c30300030d004044034131300400003000003c000003000000d3c00000003c101430003c1000300c004000400040c04000000130000c40400130c000300c500440004030000c4d40003070c10f0033c00000c033000000400c11c00c13300044000034c0c0400000003cf300107031cf0000104040044f0000000f103c003d40ccd050d140cc000030010444c0010000cc005000000000c3c140c000304f0030004040f40c5cc003400000100c400003000404703000000000105000c1003000000011000070000000cc3100400071000c0c3440004000c000100401c3743453c040c000c0000011000000d030100100000cc0100000050c405704c0003500001000001040c00000051004c0410330c000c4c0c010343040c044400040300000cf4030000cc000c0100c00c00100c00344007000c00030400730010c00000003401343f403104410c14070f0c0004100001040c1003440c4007c0100043000000000c40000430000040c01c0d00c05c03c0004cc40400003000001000110000040430040c4c0d001c00000f400000400003f4cd0cf730140301040c0c00c30100000c041c0004c0c00c0005000d00070000314003000c3f0c34c00003040400040043c00000d10c00040c000000c300c000000d01003c0cc044150034300000001011404403ccc000000c0f0c051c00000c30c0000400fc000104000000cc045400000c00400000000000000f00040000110000000000440040013000c304007001d004d545301d03000000c5c30c31000000004034140030040cc04440000c05300c04450304040c00d30103c0000c0100c400000000010c4000c04c0c004711000010031003000000cd400c0c050030040000c00dcc003c000400c00300044f0350030400000100100c0c000c00300003000044110c0050;
rom_uints[725] = 8192'h300c0144401c00ccf4400000c040007004007034104500c0100401100c113c000040d0f003400000000000c430104010d00430003c40c41004100000004000000040d00f14700440000031004c00000c141000104cc40ccc30c43d50401014ccc000c00000cc00c0100000c00070f040000000c04c01040000c00000143c001001000140400c0044c0400040d0c0c0c0000c4034000000340cc0c0c4400030d04050c040c1700c0ccc10c000400010700000431c00c04000400004415130000cc4c400000000c00c10700003044c504c00c1044c0000cc5400c004140030003c14c003003400000000c00100014c400c00000c1034040000000070c00001000f04010401343c0c03cc04c050410040cc10d0c010005400f04f44404c4000700fc0d31c00cc1c3040004000140c00000030000000004000c00c035000404c00cc0411400504d000001010001c000000c00010000c1c10c01410000700d05c00000cd4100c40c44300cc00304cc03004000030d140000c4410c0c0c40400c040f450005ccc0c504000c710c0105c00c00dc000d0100000030000c4040cc0404cc0715f00043c001000c0f007004055410030c0044dd00000d04000c4003000cc0f000cc040c00300170040c3000300f00d00340000cc01c00000700c000010430cc0000f0d0c0000040400ccc00c0400405000101cfcc0f053140c00000013c400700000c000d13000c000030c0cc030cc11000001f0c010000040c00004001340004050c004cc404c100034001311c0cc30103c00001fc00c40300004c000dc0440000001ccc05c0c3c000c0000000dc00040c000000c10c0d0000050cc0001cc07001004c01cc0444040d000001400005d304c1c14004300404c5c0c00ccf0c305000440c000005cfcdc33400040000c00d000cc44c000c5000ccc10c303101100000c570d04c050c04c1c03000000f00040c010014c00000c00f04c000000004004f00c0000d0c0d004c01100cc004010c01000cc000c30000c00400400f4c40000004000dcc07c004003004cc70005c00013110000000000040c0130cc41004c7030003c003c111c003040000c00c407000c0c0c0005011440001404101cd0400c00400c10000c01403c00000d500c00c04010c0cc3000000040cc303c00c00c1c003040104000404c03c04000c400004004c000c430c0040c000000c0044300f000044c444000c000000431103000401c50d700cc54c0510300400040000c0cc00c00cc00f4134d0033400c0cccf0501cc407df000c000cc00f001c00c0c04010003310300040c010000d0400110c0c0c000fc000043f00001400740c3cc0000c00cc0040004c000c74c0c40cc0001000c0100000500040300000c0c0440000040400031c00f445c400110070300c14400c301c00505510c1040c001c0000;
rom_uints[726] = 8192'h310431c000000c001411000c0300010000033d340000070303000001300003740001004000340000303000300403c1300000107037030100070410000304001300000f3500005430033100ccc30104051130005000001300000c000001c031010c040004001c00001c30c0010003110c010f00340100013000011c0404300c00001400000110001c000010340c301000000c00000c1000000100000000331007300034330110413000003405010000300003010430cc000344010c4c003c0053303004100000300d00013000300030031011040c000cc00004050000c10c000004333500043f003c04c1340c00343153330c003c00000000cc30000c3c030400300d03f70c040000531400000000001000043003c000000f730c003311fc0000300c0000003111000003400005030c0303000c011030003300007d310007c017003700001df000c330041000000300c00d100cc4100400000c000c300cf30400333c0c00033000170000000c01000030c00000033c330c000004541c143303f3000010311c000001100401c000003c100000001330300000001000050001040003f40000030c04044303073c00033354031000300001130441014003007300001c00040c340d00000c00000c150c040000301c0101030000fc03c00c04010d00040100140000044000f01cc33000f003040001103000040004cc53f4003011000c110c04000000000c31001c30000c00f50304000c00140c040c0c0137111003103c003003000000300003000001300c1c300c111014130301003301130400000c100000000004103004000c0d01000030003000000003043c0000003003000035313030340c040cc0040f00003100300f130d030c0010030401040d004410000700033013003c05303f000010700c330c000c00040c000000100f04701303530100350000301c00003c00003100000030050014310033310c000c0f74000c0003000001001c00040003000103070c00301000003001f033003400000c004000743034013030030c04030c0400010405030400000d0030300f103c01040c010001100c003003000000c000103d000000100100041c003f003000000010010c003400004c04040000030014000000001000d000030c010000f000c3000d000300105c3000303100330400010500110c353d010300040303000000030c000c01350000103300000000010330000130c304103333004003000c013054017000140033000001000104c500000350333300303700010003403734010030031000000c0001003100000033000730c0101400300400033104005300304030c1400000070003c300000000000f04000030001000000f000001000000000f0d1100000001073c03c4043034170c14f130043000000c0004340004000c00340000;
rom_uints[727] = 8192'hcc000040300c040100001000000030000d00000003040cc00000431000c441000043140d000000c004c400c0400030000c00c0c40c0c0405000004010004010003040100001000000000cc01c1000c0005c40004000004000300c00400c03000000000040400d00c0003c00003045041000c0c0044c00000000c0004c00cc00001000033c4cc00534f00000fc00003030c000000000000100411000001400d0000c00c00300000c0000000000403c0040c00040c00010004010000040f040000040000030000000000300010000040000000041004040000c4f30300c3c0000300c30504030044000003003400cc0000000c0c00c4030c000c0c0000c40000400000000000000c010410300c1400c3c0000d000040c40100005000000043400400700400000400000c400000040003004c00404300004400000104000c4300040000040c0cc00f00000400f0144c033000000040c04533c004c00441000c000400000400d0004000000400300004c00000300500c00c0c0c30000500000033000701000d1000000c0000003000000dc00000000000000004000400310030c3031ccf00044d44cc000000403000d4000c3f4400c0c100c40000000c0000000404011100000000030404000000400031c441c4000000140d4c00010000040030c00c004000000c0441000101004001000c400100c01000000c31c00000003000000001000000c0430c0c0000c003300004c000000c41000000000cc004041410001400000000400c000400c4000000000003c4000000040c00030000040000c0430500c301cc4c04000c00000c04000c044f40300340000000000004003c000404c00000004d00010000000400000001173000000410300c0000000c004400004000000c000c000001000c00d00404c00030000030000000000000000400301403c10400000c000c003000000ffc000c1c03f000000100000004004c00000000440000000c00000c000000001403000003000000404c03000433000c0500000000030000400440000000000040100100001c0c00c00010c00004c14004043c0000000000000000000404c00044000c0c04000000000000013000000000c400003000c0000000c4000400000000000004000000040000000000430000c0004cc00000c000003000000001040f0414c30040c40c4000403c00003c0000000040000000044454030000c7003400000000010000cc04000000140040000000000034044504040001000040000140030400000c0400043000103000c4c0c00030c10001000c003000c000c0000103000000040000c000000c00000040000000000001000000c010100000040000000c40040400040004000000000c0d0001cc000c000f04000000410001d10000000400000d000001000000000000c0c0000130000000;
rom_uints[728] = 8192'h30c43004f044c00010000030c400307c301000c00000cc3000cc1d003000000040000050c0dc00f000113050010000c100fcc0400044100700010004c00100003410c07030300000c00030330c000051000000c00450430040c00000c03c00000004140000400c000030c10000000000c0004000000000003030cc100430000404c00000400100000040000003000030400000300010c030d033103001c03c303013cc00000cc00000000c0031c0c0c000f304100033c033304004f00c000040404f00000000cc0040001044003050c003047ccc0370c330300000cc0cc0000010d0f0c000300000007000303470400c300100300c10000000000003010000c030000010000100044010f300005000040010d0044000340c31310030001400c0001dc000000400044c0000040000007cd0005410445000000000c011400010000c303c0400500040000000c14704000430340003040040c000001cc1007c0001300040405c1304300300004400013c400000c010703100001c473004000cd0001c340000cc3c0000350010003330050000000000000030001401504cf40000c0c440cc0030000c01001f00000f1000c004c00c0c0001c03140c030d0000040300c0000cc30d40051100c300cc300f00cc000030000f0300030c0304000003c10000000440010300400c4000400010c340150010f0000104030cc0000c000f04033c3700100005040000034000100401010101000d04034001301d0c030007000c0c00300c01003300010001000000c100040334000001004034310c1d40030000004003c004030004000004c00000c000400c300000050cc0003003004c31040c400000040c100000070004000000010c010304000c0300000004c000400400000c341000000430000cc0f3000f0000014f00300000cf004300c0100d003300000c004014003f01030030010c3001030114000c034007000f0301000400300004330c000400000004c10003040f00000400040c003700140140400c00010001000000470c070105000000000001300c030304000000000003000704400c000c00000c0001c00000000000010301100403c001c404000c00000300000700030d0033d0010c000000400004c0000c000c040104000000000003000c043400430f001303000000040cc000044003033c300004000cc04c100104047300000c0000c005004c000300000000300301140300050000c40000000435051000000341000c0000100000000000100040000700c1000000100340c000040700000d0c100c00d70405c0003c000300300c0007010000000cf300400000000001000040034350440c450000040103300c00000000000c0c011c0004030f07010c4c003403000403000000c403001010d00004000c150c030034000000000000c00400001000c;
rom_uints[729] = 8192'h5003000000011034c14040000cc003dc033c0c0300d4000003333d0c343000d000d04c0c010300001000000010000730104703003c43c3500000cf03d710001c0417c530030040000d0004cc10300410000c00d0373113043c0003c000004300c173c500cc0100000f000400010c0103100c03300c0fccf00003030103017000070444c01c401000100f0c5307003004030c1c0c00000000000403041447f04040c001010000040c03003d01100170000000030000c00001cdfc001007040c00000470303003c0000034c043000000c400500fcdcc1730104050401c03401000030000300147dd00015d3001007c4000000c0c01d10400041004c0cc0040003340c003c10031c000411003440433003400f114cd03004c0c3000c4f305c00371c3000d00000f0c0d00c000000000141c000d7010c04000030000500c00100100500040144141d0003c0030000110c4c0034cf00073c040cf000030300c40f00001c40400000c04030344c0cc330150000310031c03030c00000d33cc470443005dc03031000c300000030100c000330040004c0c500000003f00303033c00f00c14c10073044000c00000cc0144d04330403c301030013400dc0134000c30031cd0d04c1435c0d500130000000300301c017000007007c40401000c0000ccd71000003400d0407f0000dc04000c00044c01040313c30000300c50c001504d003000030c7c0f00404304300c14403c1474001f104c00114100000f0000d044c040103c000c031f05010c00401100005c50457110c004c10f0c310c040410044c0f31300300337c000000040104033000004d0c10104c001c1c00010004300374c5010004304f30dd510c04c704700013100030cc140c31340c001c3000703030c10d00cd03030010004f00000d14030cccc100f0cc00c000f000000010cc340031c00000d034cc04440030000073011f000434c0ccc000001f003401003004000450014000000c0000fc0040100341001003033f037440c5300003c000300030003004c000d00000c11cd044011c00000043c40434040000000c33700500300000001c0100003c340000001f00030005c4003d00430c0c03414103400570703c0030000c011c410c4c000440f000000434004000d104c03011730c1430c030c0003c10c000014000c430000000c05f30f00303c01100000c4433d30004003430c10c000314300000d0441cf00000050010d4430000343d0c1c14000401d13d0004401330400001300000003c0033030074c0c0cd0000003004c1c1000043100004d0107314c0cd00130004001c000004300c105c30000140100cd000004000c000105470003c043f1000000000c0500040401f0450010140f000000cc0037430700ccdc000000cc0f0047440c300f0100c00c30007300400c0f04003c40000000;
rom_uints[730] = 8192'h403000000010510c300400f000040100f0070f000c00000d401c0000140010001005004004003100100d00010010004c00c0700104c0c03400013310cc000400c40000000300040001000c04003000000000005c101000013500100d5104000cc440410c0000040301c00303144c001000311311311450001c10007000000100c10c3000001c00000004c10000003030000100001004c3100003030310000000330001000c0030d10010dc0000340001003100000404003011430000041014004c04000005400050400d00300010101c00004011103d000000000404300040c00000000000040c0c0007103040000001004f10000004100450000030000000013000401300000c00100104c300000000340410000500003c0411f0100310c0c34100000300401000100d00004000c00c04040c00c000030000000c0010400000003070f444100c00004070500cc4007000300c340011300c30d00c0405003000000c01c4000400c40404403d0c30103c1c3000cc400034005110041000003cd410004c010000704000100000000410100030000000040005040c010100000003003400000000140005010c0004100c3030341dc03000c0405c000000101041401310000000041174004000f0000404c0100030003c0c70100000400c00100c0000301c1001010c0000301710001033000c0c10013010010c000000c00031100c0000000c00000030c00410301100000040300141000000003000310043000000f000c000100c0000300304c004451000140010410700000000001400005cfc50303000300000140010040c03d01010043400000070000c0d000000300104dc0000004cc04030100404000040f000100c00400040f01400cc00000000010410c4301040000404cc11c0001440011c00d03c000000003c0040400c00c01c00001cc0301c0c300c011c130301304000001000104000c000f0000004000400100c04040000000040000400c3000000c000000500c4001014143040c0000cc00403100000441c0d0c1000041c404c00c03010300c00003000001000010330100001041400000014003c00000050c00000000c044000110034000c3031701001030c300000000010103c0cc011001000003004c0cc30000c10001c30300130400000030540000f4c0000001100cdf4cf3000c43040300030030d000000000c30c004540c334c00300410c0300031000c100c11003100003101000030000013d0000c00001300000010c0000004fc300010c0000300343000c0100010000000300c300011100410000000100c00000030c40004c00007004c30100300000000f0300000100c0030003110030300500000030c1005c00003000000144000000470303000015c031400000c30cc00000010000400000c50000c003cc01c03000030000;
rom_uints[731] = 8192'h140000c0010050d00100304c00450005000001c0000000004c00001003c00000040011000f00000004000000000cc05010003000400c010c3000000c000c000000c00c30404000000040000c000c7000c0004001000000030000000c00100004000040000013400c3000000c0040100cc0050000c3c00c0000c00400c5000c0c410c0000000000000000c00000003c001c00000001000000c100000301000000c0041000c0c74000c0400000300000000000000000c0000000040000001040000040410000000040100041030040c010100040043000c300c00000001000000400000c300c0000030000f001cc00141000430000c00030100041000000c00000300c44300000000fc0000004c1c043c31c010030c4c00053c00000d000000000114000c34000041000c0000400300c400000000c0001000000c01000000000000c0300000001000000400f0000c1cc00400000400d0f0300004330000000000000000003404000c100c05040030c0400c040c00c0c30000000c003c00cc00040410040cf0c001000014000cc0000dccc000000000040000300010f0000c300c04330000c0c0044000100000034ccc0000000c3f000003340000c0005f0c000444000c4c0040000001040000500c0401100c00c00d035500304001040c300430c0000000000c000400000cc50c0000000c0031100000001300300000cc40000000030000000004000c00100000f00000000000415004100c0034c0000000c00c00140000000103c0000cc0144000c00000c440000003c1500c0003030000000400c0000c000010000010c004000005000c0c00000000000c400030000000000cfc000000040001003c0400f000003000000c00c40c5000004140000c041000003300405100000000010030000000000fcc440d3000f000c00c000000000330000c0004404000030c1000000000000050c0000000000000000011c04c0000000030c000000000cc0000000c00000d000403c1400c00c000010510c0300c00000000000000000005000000040401400004000c43f0040000000004c000050c0005003300c0c4410c40000000400000040c04000100004c000000c00003000c00034c0000000000c100c000000000040000310037000500040c101c400000103c0d0000000000033cc000004000004000c3001000000000000014010000c100300000000c0000000f0000000c01000540000003c1040000400000c00040000110000300f0c10003f00c30000c000045001400f70000000000000000c00000000000000100044300000001000cc030000c00004c0101c0000410100d000000000000400c000010300000000000000c40000c01000000003001d00000c10d1c00034000000005040000000c050c040101000f00010c3000000040000000400c00000;
rom_uints[732] = 8192'h43003000010700d0000003000504dc5033304004c33300c000d003010031c3300010f1f400dc0030d04400c0030dc37c304c00c404c4c0d40000430073d3000c00c3030000410740400005100f0000c7130010444f1130c4c000000300d0c005000134c0cc000034c00003000370c0100400041110c010400100c0f04400c3d3cc03001dc0300000400030100000403101c0000000033c0104100c704310040030431014010405d100d31101000000010031d0000043000400c0c034330101300000c00000003001d4000040030010c770000c0300000014013c1c034041041000c030001c0000040030000331403043004030001003000041030d0410001044404050040000111400d03dc400c01000c13f000043c33000d4d000c3733030c440000000cc100004010000d401000400101c00303410700003f100000cf41000335110f010300000c000d3050001c004701000d00000c4c40700cc34c030400000000000cc04c100100707c0c3400050000c300000f0041030c440010001c040130003000fc404c04310000003400f0c0d000010c0000c33c03c0500005000cc0430100700100403403003d04d110c7c013000c017c1000d11c04003430000d1101100410000100400c0c300000300c04d00503100c0c0c00030100304ccc00c0c0000001001c3004313c4c00d43003050c0100d03300000c0c0000340c100004013c0300c130000c074140000cdcd0003c014cd0001000737300c7300330301d00400f00300374f101c44c0d0004cc030cf000004300c10d004c00004000c3330307400f0000001c0c000cc004300004000c00cd1f103030301c40001d33cc44300d1d031330000f30010001c0100004c3f03004f00010131001010040d00004011107304c3c4c470f03f000030300313d000cc0cc044c00030f0031300010333c430d3c00300c0c0c30001c43410040d031700700033100031f00030030130404001044000000000000cc0003300dc0100c00c31030d0c150000034c1000040c004cc003cc103d000104101000f00001001303000103003000c00030000304110301f000d001001c003044000000000c0040000030001143040c000010c00f034000003130000003c00000000043300000c010004c00500001470c0001d0003033c0701013fd00f04c000004c000c0c31034013341004400c030033000030c10c00c34c00704040c030001f1133c00c0000f31c0000c00000000304000d0c0d0000c000000c001000004003fc4cc100501704000100100f0c4110050010000d11010000440135c4000c0010d00d03000c04004400010310000000040003003300003d1d00d310f000440000704000003c0000c0037103400314040303300000030430000c000000cc00c00d00003005000000300010300030000c3400c0010;
rom_uints[733] = 8192'h1000000001054000400000000100c004000c000000000003000003000c0f01040004f303300c00000400000000000304c11c00000000300000004000d0c00c00c4004c40000400010000450fd4000004000c0044050000c0010400000c00300000400f000000000000c04c00301c0300404c000c00033400000f0c0f10400c00000c03014401c4070040000040000c00c00300000000d00c00cc0000cc50104c30100000000100000c00000010030c000003000000c0c50c00004014c4cc0000c043000400030c0433000040000001c000000c04000000c0030100000f4100010f000000000300300030000fc000c00cc00cc404c70c0000000000c710000003030004000c00004c00000003000c0000cc15c4030c0003004030030c14cc00400000000000c0130000000c4c33000400440003cf030c0000000c000c0c0700000004c000c30fc000c0c300040300040000c0000001cc00cf0000333c00000000000cc17c4000000c00133c440001004c0c00031c00f0000c00070c0000c0400444000000c0c0030030000000c30040cc0c00fc000001000001000030030000c04071000433f0000000000c0c10001f1011003000d00f00c00400010c01d00340030404414c00044040030400c000000000004000c0070c050c0c00470c10c40cc000000000000510c0004cc0000000300cc403030c00000000000000c3000014130400c000030f0030c0000013000000030000400300000004000003000007c0001044003c00000400100005310c00000c4000000000010c01000000400003c1c00c00000000c50c00000c0103004000c010000000c00040004f04000000000f070000404c440000c301000f0000400c05000004040c00000d010000cc00040040040c000c00004c000c00000400c0000000000300031000000c0f000300000004053000000000000c5f00010004000c0c0c4000c000c44000000011c000003107c0000000000400c0f0030400cc0000004c0c010c04010c03040f00c400100c03000040030c000007430004440c0c00040c70c000040300001000000300c40000000d00700100010400000c0c040005c013c00c00400040040000033c000d01cc4c00000340c0c00c100400001000c0040c4c04003400000001001c03300401000004000c0110c0070000000f0cc000303000000401400c70c003001003033000000000000000000c40000000000c0000000000000f30000004000000c00c0000c000000c0000300100000100030300c0030c04c000c0000000d0000000000c00cc030c4014c0000000000c000000c300300c000000d00000c40100044000c000000c0000c0c0000000000c3505300c000c000500c4000300000d100300000c0cc0c0010000000310043d0000000000d00040000300c000011c000403000100;
rom_uints[734] = 8192'h10300c0340014010000005c003004c133150003000c014010040030043400000704110010000003c1c0011c0010004101001130c500df0011000031040000030010040c0003000000100f010c4c000400004d0000c050000cfc0000400c44300c003004001d300cc0004000c1013300000010007404110001341000f0004341dc000c00000030000300400c014f34003030c10000010c44010c400430100003100310010010c30010d0001c000c400000030000307c30000004dc3c40000300140000000c00011c34000c000cc000dc10003303c430001d3500131d330000010033c01c3c0000001000c001d1113c0001105704040030c04100005c3100013d0c00051011443000300100f00000410040f0533530700400d101310010c4cc01100000114700c400000c0300c13000000400c40011400003003cc004c0030d00134c301c003040405034070004000400430000c00c3d7000101d7410000700401f0010c505003141d0cd10010c3d1400c1403001340f3c00000000f00c4000c0034331c030000010000000c000003011000003000143040010303130000010c0d043000043100700310c000110303cc140043703000c0003500cc3404040040030010dc00000c3014d010030407300700003100031701c0000d00101401101003040001c3404010050340011d14030100713104c0010300c0300c00000c005cc031cc130403c30d001c0001010000000c0403005100c0c0000503c30013c400030d00040003100100c010100d0000130043c0000033050034c33000000303004c0cc0310013001034001013333000105403300303000300704c0730130401000100000110001010c030304001c1001044070040003300300300100c000400400330000001cf10105f10d00cc0c3d00100c330150000c01003c05c00c031010c0000710403c01040cdc30d03044d400330040000c00000130000c30000000000040000030000004543c030010c13410c010000001130131000000cc40103d00c00003f030031410303d10c0314040f00000000c0033000007c30040037d17000000304100307140300034f70014051c000c0301071034000004000034000300137c410300000133040011400040003310003010014000000010000030300574c000330013130071310011040c000040007000c000030d7100140101003cdc030300400fc0c000103000000101030d000000104030001000c00000c041014040f0c0d300300000000000c100000001010000440030f330110010103033110000c01004c0c7c030c0003000030000040100d1330c000030c0001300000c0c014030041131000143d000d0c0004030030510301000000003000000400d0000000004000000000c10cc00f103001040010c1f000031050003333341000001c00000;
rom_uints[735] = 8192'hf0000000041000070ccc00100000300cc004333c503404c00000300c00000500000443d403000010141000d00010343010cf00000c00445030700040307c0004c0031ff0013030000001500d00000434330300003cc0f010c00dd0000c7430000c1000400000c004003400003043c1101000cf0c00000c140dc0000004cc1400d05c300000f04c000c300000400c70c400000010000000c00010000c0304c0ccf00c5440cc0004100c1440300070403c0c00004000004000c4000c4cc034000300c074300007cc0d0300003c3000307dc000c1304530c01334c33340c000401050300040000c000c00004c0001c000300001cc400000000000003000010013c00045140c300c04c0cc43c0d150000430043000110001300430100c04300000000f000000400431000730300000300007030c001c001000330000400c30001003c40040c4074cf0000014000c04000101340007001010c404001300001cc0300004000000470330c000c000c00001cf00cc0d441431c50030000004100000103050c030001000000cf400403c400430330000000000001300071470f000300c1100fc30c00440070000c040500040110000000501130000144c00ccd1400003103130000004000040430340030000c05004404030010c00c00304c0040404007c00047c004cf30034030000c0f030000c70010c04d4401001f4100040070040c10c0030c0004004041110000714300004030000530000300000300000400000004000100000c000c00c003ccc03037010d400400c03c00c0004341f40c00cc1c0300540000c0100000030c4f00c33c01004000000030c01003430000430401c00d010000cf01030c00000030310001c4c0400504c300430000003001303040c3000c3000c003100c03410350530331cdc01100740300504c00010033d43c1010000000c50c03c000300103330010003c000000005cc303040c0c0000cc00000013004c030000c001c0c301000300c0470000400000c00000400100c040070c1700001003040c000000337010030000000043c00171530300c04c0c40070105000103cc4300010c3404c0000300030c010c4100000000000000010040c5103d00c1c000000c0040040001404304d00030d00c000000000100c133430c000043003c00000000044033000c4000310003000103c0f00303003f03040000033c0c00000001c400000004010003000100000c34004040001fc5000c030030c30f00f0c00031030c003000d5110000133003310040401301000d000000700000000000d70070c3c01000030cc000c14100040000c030010c0040400300040000c01c0003cd0500300301340000134103030001310000000003c00d4300003040000000011041304043000f005000c101000303c00000c000333000d0000dc3c1c00000;
rom_uints[736] = 8192'hd0004000000000000000c000440000cc300c00c00c0000000003c000c0000101000040000000000003c000430000c0cc031003c3c000000c300c0000040000400c100000c3000c110000c4c1740000100d0040000c3000000004c434000300000cc13041c000000040cc070000400000040d000c00007004000410c00301000030c0000c000000c00000001000000c040c00000000000c000d040c00c0000440c000300d0407400000000000000030c00301400000c00300010400c0c00300400000000c00000000000000000c000040000d440000040001000c0000f0000433300300c00304c0c4000c00010044000000c00000000d0000000003c00c1100040300040004c0000103040040000c000300440000000c0300010000030040000104c40000000c0041000000010141034000000c100000c000000400010fc00cc01000000000000000040000030c00c30c003c000c1c040c0c0c000000001030000300303d004000000000cc01404001000044000400000000c00404c0000010005001430400000000000c000040000c000300004f00001000035000000000000000400c440d0040c400003f0c03044400c0000044cc000004003c440000c33100cc3400c0000c00c000000000cc0c000000001000f304030300c00005000000030c0cc0f410010103004c0000010d3001000440030000000000c34000c000c000000300040c3f01003000cc013c070f3001430c00c0000010c00c03c30001400000000500300fc0000000c00040000000c00040000cc3000000000011c000000000c4000000000c0c10303040000040000c000003000300070cd100000c40004100c400c30004000d100c03c04300000003000f03000cc04000300c0d00c300004034000001000105400003c00001fc00c05c00003001400000000100400340010770004300000100d103000301370430c00040000003000000c000c030c000004700000000000000c00000000040000c0c3440001040000301004300003307004f004000010000c300004004000000000000003c0000000000000000433470000000000c000c0c4c40000c0340000c03c000030003003001000000004000c00050c00000004307300004c00003014c00300151000033040c0030010003dc000034010000000310000000f000c11d0300000000f701100404040df0000000000000030001100000040000c0ccf000c0f400000003c00c40070304000000c3c340040000040000030c0000c004000400044000040003c30000001000c000000000400c003000001c0d000003000300000c000f100000001c00cc00030000000c0c0000010f0c000010000003000440030000000440000c000000030100c0000000000c000000cd000300d1000000300130c0000c00410040330c44c00000400000;
rom_uints[737] = 8192'h30003c700000040000007c100000000000000000c00030c00c0034000011000140013c00000010c000100c0c000404403000000050f000300004d0040000d0000000301c00010100c4c01000000030001014c4300000000431c00030000000344c04000000001000000000340005ccf40030000f00040030000000cc00400c0c300c0000003c1030003c04000c0000010000000000000000000000000c3c00343000040cc434300040000cc0701100041304000cd0c400403c04000c0c0034c003400c00400000000013000000000070003d5000041400040413000400c0000010c0000000000040000400f0c00c000040040004000000300c000434000c0040000000c03030001430003000c00004f000cc00103000000c0030504030340004000000300000000ccc300300000f00101000000c0000cc000040c0c03000000470140050c0040040404c100000c010c00c10000c0000f000400c00000c0010400000043404000c00001170040400000400000400000c00500c00c4c03040003c00f03000000000000000c000c03c300000000c000040044c00000c00000001004c043000007c000041100070040010000017003000004000000000100000c0340000300010000000000cc000fc000d54000c1400000100300c40043000000000000c0410d00010c030c000c000000004043000000030300000304404000c110000c000c0100430003c0000040000044c000000000000000070310404331000140c04f0000004003001107140001c10301000000000000c04000000000000001400003cc010304013000000f00000040000c0c00c000c003c3000300040400400300c100c300400000047000004c00000510030001001000c0000000074300010c000c00c140000c403c00100000000c4c00c00300000001000003c004000cc0004000000001000004c0c5404440c1000010c0c00003400000c01004000000000100000000000040c0000000000c0003300cc0010007c0403001304043c1c0c00001400000c0000000c043400300034c00c77044c000000300000100c040030001000c03c00000300000000000050000000000c000c0000300400440400000c01001050071040000000000000c00c0044305c000013040040103c1010100000300c400c00000c0010c0300c04c00003000c10100100c0c0740c300000000004000c10f000040340d00000001000100034303010f00030c00c00000003000031003c1c00000030001000140000001d50004010343c00003304000000100030300c00003c003000403000301030004000000000010000000010000030c4000000d4400030c0000000c004300d10000000404c40000004000c1400003c70300040000c001000103c000400040000000000003030f030f000f430100c00001000;
rom_uints[738] = 8192'h400040404000c0c000304001c00030300000000000d4000000011000c050d00000c400c0c1c00100c3c100004000d1000400300000c0400c0000c000d000000000d4c40000000040100001f00000d303cf1004c00040001000003c101c00c0000040c000c00c00004c4010000c0000700000010003c0c0c0404400001340c00001031003c00004c00000c00000040c43000000000000404004104004040300000000000000004d7000d00000400000405333c000001010f0c00000040c00104000c00000c00c000000000000c00c00d0400031004004000000010400104001300d00004140100000c000004030ccc040000c40000050001040000c30f000c0000000000000143000000c44c01400cc000100134000004000c0d000f00000100000c070000000f04000010000300000044000d000f000004001040000f0000000c4c00000c0c0000005c00010c0c00000407030c0050003d00000000000c0004d504300c0c0f0c014c00000c000400030004000404050100100c0000000005c0170d0c0301000c0004300c004c0405010000000c000400000300cd3030000004000300010c7c0c04000ccc000400010700004f0d4cf000c0010101000001cd000cc00070004000011ccc10c00000000c040d4c000530010704010000100c0014000003030f000c00300f00050c0c01000000010c000003070444010d00003003000cc0000000c000000d00000000000100000c104c03000c0c00c0c00000730000044d0c50c000700000030043000000c300330000001c00000d0003040004c000fc0cc000050c01000c040004400004003d0c1001c01000050c00400000000d0f0c00000c4d000c03001001040000004d403000043c030000000400000000000001000c7c0c0000000c00f4f30c00000d00000c0c0c04c000000000110101000000030c0000000005040cc44c0001400001c00c00400c030f340300000001001000000100000c0d0001000000030000000c040c0c0100000d000041004cc4010100c0c0140c0c0000c00c07030300c000c4047000000000c04000003000040000c0040003000c3400000005000c00c00c0001050000000000000d0d0040300500c500c10d5d0c0000000000100040040000700000c005004c010007cc000f0c030c0c0c3000c400000100100c4c00004004c00400040c01000fc1000033335300000003000c0c010000000030000000000411004c000c00c003040700004100000c71000c000c000100000d050004000400000c03c400000300030001000001051c0f1100044c40000100000300103c001c010c03000000000100000c000030000c01070c00040d0cc0000000001c00000c0000300c4044000000c04cccc00500040000000000010000040300040f0040000c00400730050c050cc000000400;
rom_uints[739] = 8192'hc1440000cc0c050105c037c1130403c0cc00003103000001005400004070010500d310c5c00000404001000100c3fd7c0001cc4141c043300004334cfdc043000100f1c030c0000c04003c404dc05000c04000c0000430050cc010000c04010400c315c0074000c04043c0104ff1014300400403c0c000c100d0000d0343540c1100f340c00d000c010f00400000401000c3c0000000c0000000000100c04c0003cc45100c003c4f0543540010c0c0c4430000000040070070c0004dcc00001000c003d00300d50c000300c00041433400c300004001004001c4000040f0011000030003400700000000c00301f0c107c1004304c13300010001134103c10003000f0c00fd40c0c003370cc07440c4440c0f4307c040d403304104c0c101000001340300c147040000707000400ccd3000c005cd000d00000f040310c1444303fcc0100d00c4d0007130134f4011430003c040cc40c104030111c70400c00340030104c03fd103010c013100000f0000c30100000c0cc304c0c401000001c40313000000c103400000000000700d4003c100404cc000434000004740000000030003c3c0c1c3000410c0c0f30c53cd01cc004003cc17c11114000000350f040003110005400c0000003400000c033300d401000c000c131000c0cd00000c44c4031000c00cc1300c00000c0d050510cd44443fc00c0c01cc734000000d40000300c0000d405c00007c30503001000047c7034043f1001c01304117034fc03141f40010300330c0000003050007000001c0c003000000014003000f00c000d051c000400030700c1000d70050104cc00000c0c00113434001330000d0c33404170c010001d5f300f1cc04040cc0c1037000031c0004040017040cc000c11013c70cd40404410030c00101cf0404c0cc3001437040cccfcf0100c3010405c400404f400004d033c0040070434414030010dc0105000100004c03c0c5f00040140f30c40004c000c0050040000000c100c0000fc70c0103c030d04400000c4343c00100144330c341c0000300cc10030070100f000fc000cc0000ccc503003100005411cc04c0c0000333c04040300d0003c10c0003400103040003c100c00c0f0304030000ddc0c0040313010000f30443001030d4c1d3010000c3440400cc33004d7113c040000c300341c003d7c004034fc047c3cc0c0047c00c00c000003143440000c33c4100c7043000435000140503c00000dfc00c0000c00c0000015444d00c0341430000004000000003001343530c0343004fc30000c7cc4f400107c054730043c14000000c0043400c0000c1000500f01100000000004100030000000005f414c0411000730300c00140000131010075000300c10101000003c0007100c00000d0d400010c011003004c040304030000c0c000c00310cc4041400045;
rom_uints[740] = 8192'h30000044000403c00007003c3d440010c000001400000000011c0c003001000040c31000300f0100000c10d00011033000401030710100000000101010000c700030303400001c00070150000c000011543010400cc000303000400001403003fc311140030400000403c054cc0000000300000071104003100d04033004005304c003000000000004000000000f000cc40000000000040000001110303033030001101c00c1103010c00c1000cc0000300000000f0f31503100cd33000000110000030003035010c0004c4c000d0001033c0105030d400300111c33000000070330001003000004c010c05041000000000410003000000030340414100033005500000017cc47301c0c300c300404100004001010300c03001000c000c0cc4400c000c50040d00000050001003010010330400014300000cc00040d3030000010107013c3400000d401d00c030000740000310000040070cc0103003004030000010007000c0c00003010300014003400c00010430000c000304d0000003700700000c10c0d007000000c10004030100001403011051300040c00001f000337fd30c3010000000300301030000003000010c05400040000030001000d000010100c0c4d001d03d3c110004140010f300040370014003c00104c14000003c30000041000010d03004d003001100300c01110003000000010c400101000070c301003100010700c0000300c30d0000000310c0110001c3c3003c40c400000040c303300103000001c000104c010000734001000010c300000400000000413017300c001f0154c100700c003c0007010000c03003003c001000100000000c01040c004030000400000100404000013d5500144040c40100000005104040000300031050000000004700c1450440500010c300110104000000cc00000c03100014c00000030000c0c3c0004400c00010000403000000010100033000000d30003c073fc00300000000030c3104140004000030400340d0c000100c014001f003c30041001350c00f00f30c00400000010000301d30030c10400343100004000004010300370003405103140c0010404f3cc30040040d0400000001100000030d00c000cc0000404341300d0c0d40030000010000017000050300d0030c004544c0d0000c040000000000040030000f4010300ff11700303000151000010003004100033f0000003dc330100cc000130070000d3003c30100000400c03004010000100c00004070130001000001c0000400c00c11054000c0411000cc005000c0030111010103000500140000044001cf00340013010001033001000000c004100100c03100f0430d01400c00003300c0111101010000c1c3c013400400130013550013404003017c03f0400001c01500c1001c0100004000000d0f1300043000;
rom_uints[741] = 8192'h1f00010010100300d103101011101001d01010003000010000d330001030c0400033331f300000400030010075000000c0000050033133110003000133300000404004c00000001000000c1100403000c0100000f0107000001000000300031c000110033000000000c030000010f000011100c03331303313f01fd300c04430010000000c33003000000000c30000001330000100003010000100c0003000030000c0f000010000c0010000110300400000130000c00000010300000f0000000300401000000c00003000103130030050430301c30c0000331000000f10000033000100713310000110004100cd0030333033000010000030003040001000130c00000010040010300030c01d00300001300040033010000030003000cc00100030300003f00000c0104010030000003001130c1030400003500000000010700403300c0010430030304030013013d0003010000100100300003001110100000100ff0134c010c030c300000033c0000001100003300c03031c00113100101000110003010000001330300c00c0004300001000000000030003c003ff001000000034001030010f30300001c0cc0d001030f03101130000c300300010f00133303133031033003001030000400100100330000010c000403001000000c01c0000030030310010d101051070001000000100010000110000d1100030030303dc1000300c030000110000010000400003000014303340004050103051101100000051c000f0033000000003000c3003004010010010100170400100410001f31c0010300000c30100030050f000300000c00000300000100100300010000040d0103000003030c000010300d030000000000030c0011400030000000000301103305000101000101033303d1011001000040001031cf000000003c01055001030c1051130011000004440cf0c500000030c00010011001030c303511f0030003000004100000000003c4330300104100000103034000001031100331401330000030000004140003303d0030131d00000000000cf00000300001010003311f000c031100c300000003010030000f000500300003303000010000100003f403000300303000010030330003010030300030000100010100100000c0000101044000031010300400000000000004000c000303050100030303401c0030030501000010114743011000003010017030003400003000003300030400000d03010030004c0c0000100050000301000300f3047031c30000000430000033000030100003000c030100000000000303010000000001170d300000100000001000010000000000031003000c000001000300000000010300010000103c010c00003050013000030003c0000cc00010001c03000000000000003003100103000d030000000;
rom_uints[742] = 8192'h401000010401c30c0100004400034040c013000000054c000000000103d04744013303403000301040404043f413c04301000000c301d301c330400100c1c0c003134000450041000000d3050004c0f0030310c101000000c0330140f30c0000007050c0300d1034c03cc00cf0404003cc1100343103005300030333cc3040017010d004410041f0100030d0000001c10000107000400013c340105073d0000f30f0103503cf0430050510003300003000c0c0400330c0c370c31100d00003000300c0c00000d03100c00100000003734317c00303103c150000304c0d0403304031000530c0000040c003014731300d00370033001000110400c4000000003040c500304001f001d000000010104f0103c050000c0050003340030014c700c030c000033c40c010005000c01000c1c300401310000c4000000001003300100001003130c140000130c000d10000000f157000c3470cc003030d00004040100107001303173000103003010075c0f3d0c000430103c0f000301033030d1051040301c04040300303130340f3130303d0000341000101030000004100000000001410000c00f40000000400c105001300f100c01331000100000103035d03400c30d10003c04340000c000000000300530c030003c004474010100700000037010030003003d10400c070010c034000040047140300330070301000000c7003c04000c0c0d00000010040700001d0301314110c0c700030440000000340340010104551400c00010000ccd1000040c341c0d1c00c005100310c3103000101003001001c031000030001cc1143130010304003010300104000cc030300c310500740000001430c01c0017400040040f0344001c3c1314f000001330300110003000000014040401c0c00430005050100300130430000010030001c0f0750405050100345700000c300004410d100c30303300370400001005010404000400000301c300001000430504c10104000c0007000f10000104070c30004004140003300d000400700504300011310f0c300130040c304113100000003000003c310001140c0c0000050110100004310000104000000100f0103301040300cc30000000f40000040000010000100010000c01000031c13000530504101000000004000031003710040000000300c30004010100340c0000001300c0030030000cf13534000004cc040700f0111003c1341037030c10000c0fcf43003c10000703300c10c0300c05000000040100000c0c3410041c0c1310040c0f00130010301cc0000000300c0f40000003c1050000131001f500141000170000000330c000000103000000011300c000100000000003113010340001010413001030001010040000c07000300000003400000141031014330030033000001003c0171c30f404c00c00;
rom_uints[743] = 8192'h311d004430c50100400f001d30010c001c03050100104c30c3303300001300300030ccd503740400100f10000000c000c033000034100c070001000014000000c10110c000031030000057100f00000100000100300c0000000010dc0500003000cf010010cc3c300130c7113040f0410070000404d00c1330ccf0144030c0000c00110003ff30030000c00300000100000710100030300003cc00c0105ccc301d0307300313c017300004000000001103005000001c005003101003cfcc00000c3d00c0c1300003010030331f1730013000033310010c4373f330437005001fcf301003000004000c0d13c0000000cc030030000075000cc0000fc00001001100100000c30003050303404551003000300003040c5c0d30d04001cf300141000407070030003104404100000c00330c3030000001f00300133c00400f1100104d0c130c07f130000c1000c7007100c0d00c04043f0400003403c410030010100c000c300f0c430000f00045c103f01000010035000c050cd0f113040303300d33013c07300040440400c0001f000140003000000000000000c0001c004504f05500031000000004000331007011100cc00000010c0c05c00410cc0340130c0000000c770303003000cc1534430110040400000cc0d31173304000100130343c03c00c00340040500100040c4440040c40000c3311003037103700033030071135d000d0300f15010c401c74313000f73101304000305030c13330011400004c014c430c003c000000001130c010003430c00400000040004001c300310030301300c0001c03003000000c1010d00030000c0030f00d0400033100013000111130300010fcc31040003000cc0c00c000331100f303c311000003140033c300c11004040310004010001300000100333300700003003f004c0001000001c13310301010340d1403004030033010004411cf000000110000030300413510000000000101300000cc300f550c01011000300000110404013301c140303330003cc004000c44040f10000001c03303504043003cd0000c0d3033fcd1c1d00305001034c001000c340c1000000f0d00c3000030003003010010c003500340d340fc04f0043044030400000001c00c000000030000430003c40c03043c4400400c3010d03010300300000c0f34c0c0004300c00c1011140041000d300000000000300004011350000000c0400c0040430040000c01013000001014040c004500c001001c0400001000034000c01f740000f3030f01c04c100333000f003c40030c00000434303000000000005000140011000c00c100d04010010c1000130000040f0300c010cc0003df0340c400f110000001000003000033004030100000000100c13410000330f010cc03c1c00c314013000000000000000300033c0f0d33033000;
rom_uints[744] = 8192'hc440004c034000005c000410000c00404000c000c00d10000c000c0044040000001fc7401040000c533404007c00c3007130c010c04d0c00003040000001000043070004000400d000070100300c00110100004c043c003c001000000000d44000004c00cc0000c0f3c5110003f0000f700c010000003300071c04d03cc000000740400100000c13040010c1001003000040014003034013c3700440004c0c000c0031000004000c0100400cc50003c00010000000c4040400c00003300300000110104000004000034c0c0c03304033000f300000004cd0f4013000d0c001010410000410003000047005010c030c03003000000040000000000004040003041000000003400011010000300000000d0c3cf070100d700000330030030d4c00004c0000c0c0030730000114130c100c0c4c0000303c0000c100000cc4000003000000d03041000c0c0000000c000000c000404c0040015014041cc000010c43044c00c410c04000033c0c4013c110400d00143003000c00154010400007340c003010c3c030030040000c000cc10d0400000000000d0400c00400c043403c03c0c1005330000c000001000c04015303300c400003d04c07040c3044000031011000000501c401d41014400c010d145ff0100c0f04404c03010c00041070000cc300010c0300110401c40033000ccc0041003047310000040000f30403041f004103c011f00401040404400100d40c04c0004c00104c0f7040030011d04003057c0d0000c000030100d1d0000004000c030d10c40c017000000715111003c00c400000d7300c3c03030000000c0000007c3c0000404000cd00d000400103003c300000000f100430000010040000575c30000300c00c030d000c4400501000000074c40040c00400035030d40005ccc4041000d004c001000710004c0103003301044c0300000000c0f00c7c400fc00c000000000c3007000c4003d70c00c0c300d4010000000001c0010100000c33c004000000000c00140030cc030c03c00f0000300410110f00010304f0fc0c003071dc04fc500cc0100004314d0c00004c0cc3000c0c0007003400000000c7001fd00f00000c04004034003000c00030000c000340300003400c43c4000704000004030040000c00100c0003004040c100301000400030030c0300037c7000000c0c04440cfff304cc0170c00c010c3003f045457fcc00041305001010000000c00000300c0c0001100cf00fcc003310034003300000c1007c00c34330c003031c0c04c0047c0c000cc10c7001000001004431ccdf110101c00d440131010004000400003004010c30f3c00000000c030c00004300000300100100004000000300000c4c0047c10344030d00300400c4c0000000070030073005010400c1c0000130010500000c0df0c0c344f00000c00;
rom_uints[745] = 8192'h43000001410040000100013003414103003000f0440011000100030040000100100051c0010010000007031300c33174c03000d300c300000101004000410003304101040fc3010300050340000000003741010c0c0c70701145301300d014c005030303030d0005c3450330000c0100010034c0000040017d013000000000d0c300030000400003c501410000000d03000010000000d00f5300000000000004f3100000040101010000c0c30c30430000030000405000100000433340c3003001c0c10000cd43001c00003f000003030d0100100100301c3c30c40c3000c0013330000c3f11c0400400031430004310403f04d0c700000000c000c04000341f0011c0000f7100c030c110000301400cfc00c00031000303c0400d4307c000013c000000040003410000050304000100010c0f0c103000300030104100300000000c31f1341f000000010f00403000c0c30001c1010070300057130101f100000071050000c00041004033c00f400400c031400d00c0c000c000030c400003ccd37043d0003d10c03300004101d003cc00c410c000001330044340c0c300300031c01010c0010300430304130040401340510404000071040401c04103d3034000030c04d010d000f405000300c3007000c10c30410000c0031103c1c10000000c10c0c3000300c334dd000000f0d144000c03f40c4033c4030000c00044031300c0410001031103040010010010000c0010001100100703c04c7000c00040c33cd00000400301010c34030000101030f10f03331000000370d03000000130043000000040c01007300001c000411040d0703100313303300d040100000104000001000d0000003503000c00c1700c0c4031c03000000100000140301100301003301000004001401003314003000000007100300400c0001001033100d001d3d0053400f00000d03040c713000001d0c0000410c000010043dc0c137000f43c03c1000000c04140c00000c0430f00000113011c040cc000140cf0310000030000c1001f00cc0000100000010c0000c10c00350c0100000134d1310003c34000c00000000040150f001c00040c40f400040c004510000040000fd3000c0103c14340000d00401400014041004001003000c0f00074030004c0004d40100300034110040003f4410c00040000103c0000c337031000400c00d40c314000300000001130c00000c00107010000004101c0010c400100f400000001c3034070f000d404504000f000c0400040330000430f03050c00cf03c0000430d0004c00000041000331c0000f050000c0cc00001100400c40000000030100000000f000d040003100003001d00031400140000011500000400103001000dc000000000001010300c00c3000403114413100330000cf004040700030003050c04301400100;
rom_uints[746] = 8192'hc030000000030c015030000101030074100000403c0000c003c100030030c000033000403030000c030000303017c000d3000000c010000010300000500000013cc400000c00000f00005041f00014c04040000400103000c00001300c40000034000140010111000040100000100d3000000000000000100050300100000004141000c0400000000000100000000010c000000000001004300000003f1043003041004000100051013030110000100000403030004030004000000100c0c0003700000000031c104001000000710030000010010010010030ccc0430f7000131000300000000000003000404d0030100d04f13000300003100000300000041000400000001000000c00030001000000004430f00c3c000001100c103130fc0411001000303110c03103000cc000000100c00030000000000000433300040000f10c000305004000003c3530300000070040000004140004c01030500000000000c010011013300000040000100c047333004000c00105c0013010030003c0104f700050c0300037f0400001300010331000700000010000c0110100000000000350011331000000000030000d000003c0400cc04134c000003100030043301033000000000000401001500730304f03f1104000004c0500000301405c1000003010010005010000003000003050001000330003100004004cc00130100000c043000017d010133133300c100113110001000cc0010c0400000150003001103c40304000013040000c01c00000001000001100310304c30000300000500015030c000111c0030003004000030c0c0040c300001033000010400130f00031c10000100015105000c000005c50001100400000f30000003c30330300350010004100000400000000131010300cc0000000007341000070000000400000d0c0130030c00300000411c000000000044440501040000070c100030000000030000000000c303000000000000000d00000000001030003400c000000300330c03000000003cc0f300000030304000300300cc0f000c3101c1000000000000000007000100000311000000310004c0000100000000400000000400000d00000100c00f0000000c3d0030ff00f000000000000010340010410300140000000c000030010c01033c0010330000d0000034c014101000400030c001010104c0000000000003003030000000c53014011041000c00030000030140000000000000000000007007c00100000130010000c000000151030c01070000300000003330030103c00000300004000c05f00000100d100000001000140000100000041000003004370000000c000c03311001c01101000101400405000000004000001000001c000c340400000133040d0103310400c0440000000000000000400014301c04000000;
rom_uints[747] = 8192'h4c00c000000000030400c0010003000010000001000f0c0007010100303c400003000c70407000c03f010303300001c4c11300030373cd041c00001c0001c00dc43040000f50015000010041d044dc0010c0000cc7f00114000040c00c000000001c0301700440000101f3010c0040004443400c4f400c4003f00c00430003033003100d005003410c0c140c0040000003400000000c011c40c001c003403001030001000103c11000c0000400000000c03010000000c30c00430d5044c001c313c40100000000c034c30000011430d0001034000031010c41000c0035c00000340000040300000030c00df30300740c40444dd03c040000c04040401c00043310000000f0f3000005c003010003c0004000300c130f51c43070005c01073d01c0dc000f0130030000003f01f004d00403000000400c0cc0003000400030034000001303030c4000000000dcd045c1d33000330140040300713140710c34c03003cc030353340f040c00440101001f03300c0000cc0043400f013100000030c1043c034047434300034c03051004304c000c010c000051030fc303d305c04000c3c3c10f030013100400000430110c30000011d00c033c401fc010f00c40401000100301fc00000003f0000c4000cd0050cc1540c0000000030c740c00010004000043d54000c400010c300043300107013501c031c004000d40010c0001030100c0034444f034400011cd00c44014f000f104c370040001c03510111005101d00403c11034000100004c040310003fc0c000040cc045040400d0c01f00301330d4400c0f4cc00000c000043c0dc11400001c003c0000000100c30005100c10341403003404340300d0f0c00c0400000100c0300130f0004300300010040d7000100000300f00003104d0003fc1c0041c00cc00301004100017101033401c0c00140004305300000404004c151710cc10504c0003000001000c33030400300031003f0000000000000c000400010000040f4303000c300300000030407047cf04000070cf0c003400010f000444304004403000044045000c0030f0311f0f00d4000033003005041c00074f00003000f70030400c031f00500c034cc300d11003c00000c01dd0000dd0003540040f03c030100d00c0c700010430fc00c0c01c400430001000ff300c000000c10110001c10000104740430401400000110000c4c10003300400001000c0000100000000c000040040010400304000704005000c0cc00130c0033341100003c05003c5001c3343004c00000040004301c4001c0114030503c0c40040c04004c001100f4001f30cf1300410433c014004113040400c0130d0c41040000003c004300004000c000000004010540cc3011c4ff733fc0103340c0fc130c0400041000003400fc30003100340130cc04034004043000;
rom_uints[748] = 8192'h4741000040300c4c000000003004300c0c3c070000000c030c0df100c03401c3000c03101000000000cfc5d4440fc70d41014004f50004c30000000c0c00000c0400f40000033000cc0040001000c0c000000000c30d0341000030c04010f0040040000c11c000c41404f10005cc3c7f0304044000d4c00f000044c00c4f000010003c00004000c740000c70c00c0c0f4100000000000f0cccc4030c3043c0004000471c0003304c0ccc01700cc004053000fc03000000c0000000173f001c0000c0001d00030d130440003cf0c003c430037c331010f0d0000001cc044cc000304000043cc0000000040fc4c03014040000150070f4000040d3030c10000000003000400c4f0030c00d43f400440001110104c1c000404004d000001044541c0403c000031c0c00404130c30000cc0000111c050013100400100c0044c51400c03000c03c0f00000cc070f00d711c0004c40cd004c0c00dc003003c3000013c00004f00c01c340500f300051d040000c7043d00410430300000f0c1f04407300003cc40c405300040000030053005001c00c000000001cd0d0c00300114004c000103c1f07001000150c0c0435cc0c0070d000dd00d0000410004c300401f040dcf0300000000000c4c0000c40c0c10053003000c4c0507001410150010041c410474040040003cc10c3c140c33c00000000051c3004005000000c04141310004cc04c0cc7d01c00400007c0000ccc7f4c00140400030001000300c00d0f0405cc40d0000cc040f0000f5507c0c0000134c70000001740001440500444033c43c01003c0441430004ccd14c000043004d300000004cd100fc410000400440d50000010740030003f300c0ccc030c0c0044434100000000c000f00100000000130c441013401c0fc4050c04c0c0c43c0c03cc00010c370c000104cc0c0140cc044c114d300c00cf304c7007000c000001401f0000004d57110400440103040c7140cc007000000000004000000c0000300010c0c00c1400cc40000d303c130cc00003c00d401005c0f0530500c7c004c00010000000100000003cc3000c004004d0040045030047dc0000110f000000c0ff000004000300004c000c00c0040010c7cc000c3d14000007f007c300c01070c0c30dd011740100c400c0400100040d7304c00d3c40770000404004c003100c0cc0400044c03f30001000c00c13300c01400c30705000c1cc0004c4301100c400000400030c0d0340d000004040031400cd3004000cc00443000ccc4404c0000c03300000fc010c000c33cc004000c000130000000cd0100004143000d100000d0f1304000c410000c00000000000c0004d010407104d000000003011000d41041404c00000007c0104c0004f004c30c30c00c4ccc3050701403fcc04043c0c10c0c03304000c0310007c500f03300;
rom_uints[749] = 8192'hd000000040000000cc70000c00000000300030100004000c000400000c000000000c430040003c00100400000d040d0403100000003c044d0000040004001000001170740c000004c0000f0010003c00c00030400c0001000003300000000100c00c0433000000007300c000000c00004100300400000040000010300100c400130c0300000c003000100030030004c0000000000000000000040300100c100000100c00003c001000300000d100c070040030000004cc10100004100d04000040000c433000471070f000000c307c403c0c53c0044000000cf43000c00100004c0000000030040c00c000311030400003043100401000400040043cd0030000dc10004000c0300c000000000c00000000044c54000003000c1110000100003c133003003c0404010000000003004c000000400c000dc400f000010040c000f0400c004000400000403004003040c00004540300034cc0c030fc03c400f000000c03700000401040041133401414001d000000c0c00000000403100000c030000000000400400400100400000f00071000004004000000040003000c00000000d040000c03030030003400400000000000c40c4cc0c40074300001000000dc0c000c1000c3c4000d00c00c00c40003007000c000000045c0001c4000000430000010301d0c00040000041040000004034d000030c00000000000000cc0043c00c00000031400030330c4cc01f00000f001c7000000c0000100004400030070000c010cf0003400000001c01000000000100030c0004040340030000cc100031044400000c004c40000100044000400000004000010004c00000100400001000334cc000c403c001c0d100000400000000001040000003440000003005000003f003c000030034c3f04000c1c00c0100000f00c0000011410000007000000c0040100404cc3000c30013c370430cc00040300100c00004d000403000100003001300cc0000000000040040000000000c00040000000000d00c000000004c01401300010007c30000100c300500003000c00000c400c03000003003000300c000000010040000cc013000014040f00300c0000000034041000007000001c1c0000c0c0000300700000000000000010c000000c0000013300000000000000000140000300040c0011040000c3000000303003303c00c50004007003030000040014000004c40d3040c0000c0004c700037000000c0040000000044000300100c007cc0000000000104000044070040000c10003331c4c0000004000000000300000f000400400c03000000000cc0c000c0000cc0c005c001c0d0400000000c00010000000003004000f0c400c001000000c000c104000001400004c00100400c000001c0c0070c00000000004000005000c000c00000000001000101c0000000000;
rom_uints[750] = 8192'h30000000404000015cf000313c0000c0300000c0d030cf4400c30000000c440100100071000000000c4d007400400fd3f7040001000340001000c0040301f000040000400000010000004010f000001001c03100013c0c000c307cf0000d0001003701d1000003003000c70300c000304004000c001c10303000001034500440300000003100000f00000001000013c033000034000000001040c0c0f3000c00005f03050010001000cf0070cc0100010040004000000c40d0000100330000000301000140000d3000040c00c010000d0340051c1000300014c41c10000000311030000103400100400400d140c00000000004f005c000010000cc103400001ccc000050c0000040c00330c0000004000010000000c30d3c10000000010340400003430034c50010304030031010400000000000400000000030400030c00004c001030310413000c0030100c000030003000010d040310010004000c004c000040400030341c074430000010000c3c00030000030000300000010430000c031ddf0c110ff001000c000100c0000cc0301400000000000d400010000001000c030010cf0044010100003004c0741300030c00310100000407500fcf0c00c37005400034003003700000010000100305044c0c500c01c00f00000004400400130c000010100c03c43c01300cc14d3c004c300c003404000000f53c000100000030c10003cc00fd3f000303c410045400000111000010000000cc0c03d00001000400000c3f03000000040100051100c0170300100000030000c40401030000cc4307340103040c045004000040ccc0104c3f110cc0c400c1ccf1050000010c304d044004103701030f0c0000100030040c4c0f101c0f000000c00004404003110c4305407000000110043033071c34303d0030314d0c040000040c010004050c07c01c00010d0000300c0110000c040401000c01c0cc0c003d000c000040000000cc13000000040c100040010d400c0d000c0044003300030143000300000300131000000d0400000000301000000d00300c000003140003000400000cdd3000c31c04044000000000000c0100000c4f04c03cc300400c040003000030000cc04051c400050c03030007c0400001010c0c000000c00400000304103c000c0d3000100c0d300c30010c000c300c110304000010c4cc0504000000101001f00c310c00003c1c0000040cc4000000c003070400010300000134000000000000030c03d40c0c000003c007c00703c0c0053cc000c50c0007c30000000000030010003c4104411310010d00000000f00000104004310007000c00000000000030cd03000cc30070330741d0000c04c00c000c00001501140000150000303305031300010c001000000c040030c0c000000d000c01310000000c00003000010c1040030;
rom_uints[751] = 8192'h40030040004010c1000003d0410003d030300000000000000000000000c003010014007c000400000000000003300cc10000030000034055500c0300030000000100330000d00040030000d400005000011030000003001030310c0010030000403000473403031c000033c030030001000000c30003001300c01000034300031034000000000070100100303430000c0000000000003004d004300f103010000c0000013000100100000530010003d00301134000000003d3000401301c00c00003300133004403014300340303000300400003071040000030c0030310c03003400000000000000000c014101310030000001100400003000000d100000000c000150100300000030c0003310000331000004300101004000030f34050000000330000400400010000003004c0300000000043000003001000300400c043035315000101701001c030013c0110000000000003c430f00300c0f13313333000003003003c00000300000313c0450103003c034010004103004007c003030040c01007c0c00000000014300031100510c000000300000004004000c0001410130cc00000c030000100000400000510031043001c403f03000040000000005003100040333100000000c033001410033430001000000000400000003000000001c00010c0300301004040000313c300000f00d1004004000000d000f00c003000c0003000100000104013000044300f7040000000000001000000530001c0c00040010000011300000000c0003004d300004330000030300000000004000003c0c000400003304000004c000f003000000000c00000003300100011140300000334100030100f03331040013000300000c0130c000100d00100031000301001f00001000313c03030030f4030710751000330c001000341100030c000c1c0c0100301010000c30000003000003000300c1500003000c0000303100050730000403011000000000000000000000003c01001c00700100100431030003110001c474300100cc00300c310c01031710000000000313001100000c14010000300010300001000340000300c00030340c003040310133000000000401c00030330003470000040000000000c00000030d00000004070c10001001000103000101000003cc000430040111003030000100c3000000030004000030030043300c000000311000033c000005034300000000000001000000001100000013c000010c030000001040c0000c000d0c000000c3000f330010004300010003c03101000c00000010cc1c0c001000300000000000031430c110000010010000000000000000303003d7400000330f10030f000c03000004700c0c00000003010000000034300401003030010400013000100000430c000c000100c00030140c00000c33000c001;
rom_uints[752] = 8192'h40000074001134300c4fccc00014c0000100034cc000c7300030430170000400cc0000100004004000500000c000c0c0f30d010043070000011000000000000f00f00400000000d004450003410ff0030c3004105000d030340100000c000c10410d00000d0300d01c30400c000003c0c0100c00000311313cc710c0405d30c40000300030004001000f0000c3001c0000000130cc00c13d003100400340000040000103040004030004c30c040017000000100c10104100040010414000030004000000000c0000043c10414000000144014300c00003003400c44103fc30030000d4000130c3000f4000050100050430010c00000040400130000011c1c0013430c100c00000004c73c0300405d0100030c0c1010045040cd43010400cc40000003100000c03dc0000440000050000000345100000403010c00c00000c073404030ccc00044c00004050c1000343131131400000130330100500c3c300700010045dc0443c003c000c00000410401401004004040d0010004d1030400040001070730000c030010003304c001000010000000000030c1c003001041000c4004c0303000400000000000443413110000700c40000353000cc10004103104430100c303010c3301000cc1cd34000c03c14000071c0000100000000004000000c400030005741401c4cc0100700541040040c1001400000000000f4001c0d0003ccccd13d00f0dd00441c1400000c010104d00017000d00050403030c0540d043cc00f00403043f00040000f000003c0100003c00030004c10cd000c1300f0010003c000000041004050c003c0000001dc0000100100300350f100c043c30140010d50010000c000c0040030300440000140c3000000044000000f040400cf300c1c000400001c03100300100000000f004040003100000d0004c4031c0300030400d0fc33fc00c3075041c04500d30013d100070041c000001411003300004010000004c00010100000c070071004fc054103040f00d30031fc0000d0cc70001004d03000000300403441000003c1fd0030c100500010003103070c00000300000c03503c04c400c10000001000110000350001000c003d400f000014450003000c00000000030030401c000c000003004003c01000c00100c113074003c030400f0003100014001c0c100101000300cc00c1700d00300040000dccc30000c1c100004001430c01000000071d300073000000f50c0530000040100c400d0007010c00000010154001700000005004000030001cc0104c030c0031000c0054107c4040103000c4005003300f01c0031c040dc00000000c4030000cc1000440430f101043c4c4011004000300000000d003400000003003007001c01c10c70031100053f1000000cc0001c00d030cf10c03000004000f000000100000340;
rom_uints[753] = 8192'hc0030000000003011000000100000cf4433300701c01c30000df4400d000030400c1000100400003307f00310340300430430000400000cc3014000300031000010010001300c0c0000031c100000c1001dc3035510f00d0004d0311004013f0000030dfc00330000404c100140300cc0010030104c001010004043530001003c330534330040000000100d301000c040331004000f00040c50000c000330053000111044030400400c000000000003000110300000310103400010130c001c0011f0041300044370145001c003001c0031370f703101010037f30013c00000000000000000c400030100030000c1000c100f0c0300000414c300ff1070000000140c004053030404100401000100000030401033c1003c0010c5033c0c3c0030014f00000c014c030c0000c030101c00c0000143103000000004040300d053031d110400001f1030f40005000c00300c01000001301101fdc000103000400300303c00071000000030103300400400c0003300700c1041131c4c00013000c11071000300d01f401c010000000000031730010c000030c00300011130cf0c00000030d0401000030003c00010070010001000f10c4000d003101d0003030c30101300040400c005c01013100cc000c30cd0005130300031f001700301d4430040000c00000c00104040314c301c70000030017330330003100040000000f000310c0030100114004c00c4004dd05400110000043f300c00d0dc0c0410f001f0000300000033171c0007c00000300053d01001c03013d0000c30034000100c00001015c00f04f0000104000c00c0010c0c000340000404100010104c01c000fc5c0430c0c500103c0000101f40f400000040330f1d41f3000100f030404c10300047110cc00000000003c3c4101000d30000c370003300014000404004100cf000310c40000013000000c4f1000c004040011034c030c045330000c3003730003f00000000000f0c030c0400141c0c30110010040100c3c4cc0100301000c500000000000f03040c13c4011403003000000540300000000100c1000000f00c00c0701400000300010400300000044040c13000000000000000040500d10f40004004040c04101700003010000010000000034d03000cc00041c503003313034f00304f0030000000000300040430410000f000001cc00010111044300300f0004c41000030c440403030c0010400040c040d00440000100300117000c000c00000d30300040004000433300707003000037d0041000f10d004f003110110400c033010100000150c700000000401000cf00401001d100d30001c003000330030000000000f003337000013710d010000000434c030001043100c3cc40c013005c700000001000c40040d00310100cf40000000007070c000c000030000000100c;
rom_uints[754] = 8192'hc0300000c0c44000014000003040c030cd100000c0c000400010c000cc000300000340fc501000400344000004053333c050c000400004c000c4c0030100000070000040305000040000c1c0cc0013c010c07010f3d0c0c030400c00000c0c33003010c00003053010000000300c000000040004003000c0c0c13000144100c03c400000d0100040004c0000c0100050000000000000f044503c04cc40511c000c0000001040000010c00040c00c30400040000000cc0040c0c003000f0000007430504030004030300c0051000000cc0000300c301cf030403000f030c40000d0000000100000400c34000c000f000040c0c0c00cf40040000010000400000ccdcc0000c0000c0040c000000c103700004100c100f0ccf140140000c030010000c7400033c0c30030401000c01040300400000000034000000030140cc3000000c0000000303c00c0300050000000001c00000c110441fc00000ccc003003400044000400c000c003044cf0000c4044040c00000000c050300ccc0400000000001040c0530cc003040004c033400030500070c04000003070040000c33c0cc00c405c003010001400c00000000030000000cf00c3040040170c0030000d0030c40c00100cc0c0000030340030000c00c40004003c0ccc00000000c0c410cc0100c040500c4010d0170cd0000000c040d000000c304400000ccc0c0010500ffc0c03414c10d040c0c07c0cd0401c0000f4000040000000000000c0005c001003004040c0c0000cc00000001000c010c37070c00000404050004030000000c0000040400cf0c00010000040c0000000c0c0000c100c030051c0000000000c40c71040000010d0000000000c000010040000000f00040370001001c033c0c000300040d00000c00000004cf0000cc0c000c00c0000d000cd00004010c033700000cc1c04043000c04040f040c450000010000100c3003c00410c005430003000000c0000004000000003000000304c0c370000c0403000d34030041004140f0004500000300cfc001000000000d00004c0c00d0ccc00401000000030c1101c0000000000c403000000c000c00c40000c4040f3d0c04000f000000000030000ff00040000c004000000c0c0000000dc00000004000cc0f44000007000cc4040000000000004c0f0000000c03440500c0d000c300c400050004100c05c00440c03c3c000004000c000305000004000000010000140f04000c40000000000004030c040c330c00c00f0c010cc00000000400000c00000c0403000cc303740701cf0d004c00010030030c140100cc04c0c10c30003400c0000030000c0000040001010000cc0f3000000d04001c0c000500000004004000c000000c000cc70000000c0c4c00000c033cc1c30000400340050000000030000c0c0c00301400c00100000;
rom_uints[755] = 8192'h100400003440000330c0400000000030d0400400ccc0cc0340cc04000040404053005c00c403c03000001cc004000000c00f10cc000c4013cc10010c40700000c3300c00003440c00437100c00004041c0340010cc000d410110000c030400c030100c0050040047cc000000000400300c0300330000730404474430c1004f4034000c0c000030001000033400010c0c004400004010000700d04403f40c03d300504003c100434000000c3f0c0000003cc00000010700330004043000034313040c0000c300004010ccc0404f0010c40d34c0000443130c0c01001040010040c000104000000000c01044130c00d0cf0c14440c000c0c400c011004000030d434340470070030405f0f300010dc10143100c000c013010c03005000c001c04f70100f005014100c3000c000c00100031400003400000c000000c0fd000304c0405040004c0000ff300000004104000d00cc000070c0ccf00300c0c4c0c130c00740d010003000000000010c4110c0030f00404007f00c03d040c00f030c0440c011c03040040c300040011000f01c40030d00c00cc00ccc40100000101c00c010f400c0410300430113404c4000004001074c0c00004cd4007100cd00010c000040c1001000000001c00c30c00003507c000f0501cf030cc03c1010cc00d00003004c070133cd11c0004f10f00003c0400cc0cc404cc034cc0003000000100d40d0400c07c0c014d1c0030f000c130000c3c0c000f400c0013411000d1001007140000330c1000000000100070c040c000c10000033030140d37c001440cc33300400d0c033000400004304c303430c00000740000140007404400d10c311000400fc0c3c000000010c00000100003fc1d0010c4304001403c00000000f14440f00d0c00015c00c03314400003000000400cc330030c000c000c0cf00100c314010c01330c003c30003c0000c40c30f0040003104c0000000340000040030105000100001c04000c0000000cc00500c011cc0034d00d3100c0003400100000000401310000f5303cc45347000c4c1000d00c017003007300f0003c000000c400400000c0110c00000c0100c00000fc3000c00500034000100c0c440cc0c3d431004040c0f0000054f031004450000040000c3301c40130310c110000d01c0140000c37033c00007d3c00043010ff00c1c3c0000040003000300003000401000c0c00c00040000c100001c10c00040d00f0c03300000041c70033f000f4c00070c7100500050000c050170004433000030000000c03001300c000c0000000f00004f30c05100001000504c01000c00010041045000000000051000000cc100c5000c1c0f4040001004c0040500500300c030000c0000400300010c07c0c00000c0000040103000003005430c50c10000c0000000c04001775000104004400;
rom_uints[756] = 8192'hc0000434330700310100401004034fc00000000c04040003000000c30f4300014001045000f000011c00350000010c0c000f0c1c00031404304fc003100400c0c000000c400f0040003000004000030003c407070000000c1c0000000c0744000050440400010005cc3d00c0c031c1000000304734000700400cc00000400305110c0444030c030c03000004000d044c04014c00000041033040100c10410400c00c004304c0000c00101000070c00c0000400000000040c000001f0300000c0410003c01003000507030503c0c000003001cc1003030100430d100014040070310000c140000003f0001c04f00103030fc0d00001010400400000000300400053013000c04f1040400104c0c34c00400300000c000700700100730404c01100013700000c400003010300310034040310010004000000030004033100000f10000071400144033003400cc0000000005c000300c00c33430013c00c004304c01000000c014010030c00050007300c00c10f000c4405030f01004400000f00d0c00400d03703100c100040010001000503c00003014000703003300003004c33c74c017000041000000704c411c40701041c0c4c43400004000010004034c140cc040f0c0300000c4c000307430011c00103133c337000000000050104010731001041000100034c5043010f000001000013cf0300000c010000c00f00c0f10701000040000400c100005c1d0d30c1010c40cc0000011c10304017f400000410071400c04f001000000c10031040400400500c00030030103030000000730fc007000cc03d070344440cc130d0300000400030004f00000300cc0300003f0400400c00750c00040c401c310c0100310000440700c030010030030004700040010c0100030c00010c0c00000540441000540fcf010004040000000fc1011c0f01d0000170034340050003cf1501d0000c4501034000cc0040cd0c03c400010030c0040000000010000400310140c070010df00400d1000003000300c00c43030300000003114c000000f00500c3030c000c341c05000c0301003f300000cc001001340047004004030000030c0031010c000300030300000c030000000140c0040340c400f004043030004000530300000000010c000000440d030340350070c40c43500c010003004170004c00cc300000300004f500470c1003000cfc0f030c10000300c000c0100000000330300000c0c0303104cc0004c400c001000300041c14000300310c1000030400030015001000c003040400004007030700300003c0440c3144c30000c001003130f000000500000000001000c0c4003c0c001300dccd000d3c0010c1010003000000010003000000c30054000101004303000010000311c040c000c0c400033000033040000c30034000400340430303000000;
rom_uints[757] = 8192'h440100000370030c03c000000000047035340301f30000f000000cc0c00100040071c010303300c0c004000c4133f0c54401d0101030dc0300100000c000c30004cc4130000010400000f433f130005030130ff0f411000c410500c400000030000c0030300000000c0c50005dc4001fc0000004c00300040004f30705400300f0d0000c7c0100000100044000000741d003100000000000d0011404030030000000410310c0c030000c0040c1c0c3cc004c5003000403c7c004033c0001d0f03c3300000001c0c01000003500c000c104c100050000000fc00c0040c00300300703000c41000400000f000100040c0401c1dc050c17000040000030010400040010000304c1004041cf0000430c3cccc033410004cc3410f4300000c410000134d00c000c4c4030301c00003303000f01cc0410c033c40000040310035000c01c00cc40c110f0001cc0001dc00c0300000000c010034033c3cc1f00c00104040000c00c4d3400040c0c3f5310003c701c00044000001014c004070303303300f433c1004100c0001400c0c003c0040300001310000050100f101003411340c0350d0c400300301000310cc031d400c00c433d00fc0000004c00400000c0dc433f00000400d0c3510c40300044004413c04000004400030d00050000140000c03040c04dcc3f3000041c300d730400003001003400303030000c0040c103404344000cc0000003c04cf040304c0d3c141400c3c0c300cc410401dd004c01710c00c014404010013c0000070100003000000000003d070d000310403040003000cc1000300101300450000000c44030130000370030cc4400000c00000040cf1000000c0411c010330c031354d01c00c0c0000d000407c3cc003034301003000000001040000110403d3040034000c104d47331c01400010000400004070405c3300c0000700030c10000700c1370013400433440000c0c00070407130301301001041ccc01000005000410c34040143c0070330c0000004cd300c114c4c000044000f400c0300000004f04303004000003005c4100100000000000034c4700010000000030044c0f03400c04000d005000300100350003040040c104030d3cc443040cc00043011c000301cc01f0c00000c470300004004071030400047c303701303c1f00010003004000030400040003004101105c00100000014000400145007043000c0300d413000c0cc0000400033001fd0c00c300301000c40044100c3500400cc010030c000700c000703070c00f0003c000cc000000cc0000c0d0000000000c0400000440004300cd00100300340503c10000030000c0004004c000054004000040c0140c0404304003004000c0100030100074330c00401300440400000403030000000341000000cc045000000030003f030000010040000c0100;
rom_uints[758] = 8192'hc10000040430c00410000004000dc0d50c004000c1c10000400000f00030c000f414c0c00d00004cc4000410410004110010cc0c0d0030d300c0c0000400000440c0c000c0000330000070010000c0040c0401041400d0100000440c4c0cc40c30c0040c000003400310040c04400010031c4301f10c00001040c0000104c0c4003400040c00511034000400000000c04d00000010700c0c010c00300cf4003c4c330000747030003430303c03000000033c00000c00040c0001044003011000c0c4c13000301103000030c0c133c0400c444000c0f000001000fc0c7000000c50003050043030c0030040c40000001c3c4f001000000c00000c00c30000c000000c00dc10003000100000040040d0c400c3004c4c0d005f30040004c00c040004030040400044ccc00443000013c0404cc0d10c3c003030c030305c00000050c4000000c40d044000014400d00000c00301017044cc00cc00d01003f3d000100003030114d000c4c0c030000cc04000040007c000003410c44000c01000003034c0000401010050010c00004c040d1010f040c000d0004cc400404000301034c010c4f0400030001100404cd004000c10c45000d000000004c7030c4c4cc0004c00000000400cc07000010c1001300c030000c3000c100f000c000000f10c10500010cc4000d50010cc0000cc10c004c000140000d3143040000000000040c00000000dd0c0c0c4000c40001040010004c05c00d000430403d304003004c00001f0c400cc0000001004c0c00000c00004c10000001050cd0340c30c0004000c0407c003100000cc07000000cc0030d100000000000000010f00010c3001f3c0104030d01cc0004c00000000004017001d300c0400cc44c34c34000300000000003000000300c0d10000033400404c0c0030000000c1000000cc00c300000000c4c00000c00d00100f011001100cc00cd10303f03c30c70010f000350cc440340000300000d0d0400c0c040011cc0000074170c134000d00f00c0404430c000500033070000000000c04034c1001cc0c1f103700c000004700300010c00000037c070cd03000c104004c04040cc0c0301c40000000c00403400000030000f0007000c041c4c0f04c00d0000000c400000c1c0140c04003c44030cc400000007000c00c00044c01000400c0c0f0d000004d000cc01c001013400c034100c33010c00030c30000300c0040c000c00000401400d7000031c7050c00000c00d00000c0f730c0000000c01000cc51705cc00000000cc1f00c005000c04c001300004330001c003f000c00cd000000c0000100f7c000140000f000c000000030cc0c40040000000030f3c000001413f440c401000000f001000d4cc04000ccc40004333c4044000000100c031000034c1d0c00000c4000c0c4c004500c40c0000000;
rom_uints[759] = 8192'hc000000c0000000300000445030301000000530103c340010c000300c03000c3007dc0c150004000400000c00041004340000000044d5c40000001c0000000c000c0c0000000000001004d40c00004cc03c00cf003000ccc0c3100404000000114c4000c0f00c00001c300c00030c0001004040040000000c0403000c0c0040004000000400001c00000004003000040000c00000f0040000000c0400004000053004140700040000140030300c000000100000003400040000c000c00000100c0000cc000000040000000003000000000c3404000c00003000d00004000c10c0003000004000c01000f00400000c0f03000004000000000400040000000000040000000004000ccc0010000c04c0104dc000000400003004400004143000000c0c0010000004003070c03000c0001000000000f400000c0c0c44300c0000010040040000100000000c1400000c00004c0040005001000c14143c04000c000014400400000000c4000040000cc4140000140000000700030c0c040040340040343c030500300040000000c0c04c0000001000000000040c40c0cc03001300007c0000040c0010000000100c3004cc0f00004400101003000c0000040c040104c000001000000003001004400000001040000d00040c0c0000040c000000c000047cc4000000100000100040000c0cc0000c40c00000c00004000c0000100c0000cc10030000040000000004040c14400c043013c0001dcc07150000005c00000c100000300010000000000000040001040c0c0c1d000c000c0434100cd030040000300000c04410000c003c303c1000041c30040014300c0700343000004c00100000404c0000c4000cc00c0000000400000c4030030c0d044c000000000c000400340000040004d000c00c04001010cc350000073c00000004004c0c034000400400cc3f07000c040c410000000004000000003000000c003c000000000c00300000000000000c000000001000c500040c110000000003040c50000c00004000cc000c000c1000000000c00000041c003c000c0c000c0f000c0000000010000000003ccc30044c00040c4c000400000000c00000000000cc001000c0300c300c3404145100000000000c000070000c00040c1c0f00001c00003c00100030c003330000000400c000d400440030400ccc000c30000000001400000c0004000000043030000000000000001000000c000c00000000040000cc0030001c1040000401310c0000041400100000ccc4040400440004f0d4040c00d400c4300000000310000c040000100000000c00044000c00ccc0000000c000030000c40140000000cc4c0440c00000000c03070000440401400000c0410001cc00000000000440c0000000000070040000000000301000000c00cc04c000004044000000130;
rom_uints[760] = 8192'h443cc05000304c00004c000004d13104400010030304000004c0000000040400c010304540000cc004c00030c105c10303000d050400c0400001001044040000c005f130004c00c1000c4c05700c00010c00050040d100000c300c000dc4000004c053054c000c7003cc00000010030530c00c15000040400000cc00300c0404d0c30000330004f0430004310001c0c0010000000340000c401000004570cc00c0c00d01004c0fcc03c411000c0004400f000000033c35010070017030000f1040c00300c010007c00f00000000004040c0000d401445044300cc3000030400c4cc30030014010000cc00c0414040000041000107c030073400000000000005001400cc05131cd0103000400030cc00000013cd40300400cc50143c00010000351c03000c3000f00401d0000cc000040000f0000001000000401700f34010cf540000f01003c000500c0010f004f104cc00f0004f533c00000005c33c0001040400010003f40c0450043f01c04500c41c73000c3cc70101030cc500300c00304000340454445c04cd310003100c0c501000001400003400c0c0001003010000304010040c00500d00c00704001c130000041c0f0c3154000000370004c0503c10300010c010300400f0c000f500c0c03530100033c0000000130500c100000f300050c0000c004c0f01c4430000015053000100000cc000c01003004000fc3c1400000300cc000033043010000c30fc3c50c000d34cc00404f0403700004330444000cc00f003470050430414c1501000400400000413300c0000f0c000c43050040cc00330030100000340c03c1034004c1000000c100000c5d00c4000300053100cc0411c0114010003017300000c143c3c003d014403cccd04000100c0f440f13130110004007434530340340400c044c4cc000004740033f11ccc0013cc04000040c01400300430005c40501040040c443000404001d000330000dcc00d0c31000c3000000000040c001c40300000003401c03040000c40101000003010500000100fc00043101000f0c00000007100f04337000000300c0f00434000000101004100fc0330030004c000fc0004001040000c00340c00000010c50c3cc00d0003001433043030c1000003001000001000fd04330414fc0c000c000001c0ccf000500c30050033001f00f0000000000cc404010014041c010000003030100043000ff00c001000001000440007c01c301300010470d10071000000f05030c31004c30000f4004000400010c300040c5003444030004043340404131c104410fc030c01001040000030c030003c0000001003040040400000000000f10000300cc0f3330c000c30300c3cf434003010140c00005140040f303100100c000100001000043c0000010cc01401040000f000004300304041000410c000000000;
rom_uints[761] = 8192'hd44c4000ccc310000103100030003c4441c000300000c0000014c77300cd01400c30340004cc000000f000c0d030f10c00c4001c3c307c0d0c001c3c10440030101103400c000000c00001f11300007004000c04440cc01010304450c0ccc03000310040000000300510113000cf00000c0000cd00301000c00734c0d00300c011c4c1cc0c00001000147000000440070730003100c3c004c000c0101010c03130d0430500f00d0100000030100c300510c110000000030000040000d1d1004403c10040000000010c10004400000c000c55004330304110c3cf0004c000000031cc00f000cc00000c0030cd3000dcc0c0c00f5707040000010000044030010000010030000cc0013000cc30030003000040001cc003300cfd100000d00f0000040c3000c33300c4031cc0313c3050030003c0c0000410000030dd01c3c1000c1300000000ff000000313ccc400000000100003c37c400c100004000000041031301003c3c0400000034c001000003d000f040c34000c004c1cc010c7000c030f3104400c33030c01dcc04cc440c00c001003000000010400001c040c000100000430d0003304044000c3400000103dc0000040435010033040000001301d07031500030013040c330d1001c30000d303001000003014c3c103000c00000000000c40031f040010100410100c1011014c3000c000431000001104000040040cdc00c0c00c00d00003004010001cc010104300000310014000f0050c04f007000000ff0100cc000400010010010003400c300010f000c0c1000000001c100c00301c000000000003013c00c13404034340f000000c000010311000d30c140d00303d0c03111100100000000000100400003003350040000003010033000104070104010000000307500c000000100c000cc10700c4000000040cc0400404ccf04dc00030730711030c0cc45133030034500c3010c00700010030000c30000c0004c000000000000c003410044c00500330030f00000000010f03f00300000070400001003fc3c00cc000300005400044040000c004040000c0000000d734000010001f0c03f00f010400003100000030c1c00000040000104100100010544c010100cc000000c03000013000000c041300035c07010300030c00c01dc00cc704000300003001c00000300000030000c000000010000100704c03000c0333d3001c00000053c010001c00030000040000c001000100401401d1c400000050c5100013000400c00010003103000003043130000000300030c001010c004000000c0040c340340101004400100cc104c40010000cf00c0000000001303000040000010540003001f303c100c00c004374005f0000000000f04303000dc0030c5d00070d000001000001404341c00004030303003010004c10c1c730710dc00040004;
rom_uints[762] = 8192'hf0f000300000101044c00000300000c0400000c003fc00010050c4f00030000c00c51c00101c04000000c4000403c0003c040000000100c000000000cc00c000040000000000000000001c00f000400000c000001040c0310107c030000000c000340041c0001000000040033133040400f000500003000000440000c000000034400c300000000000c0000130000300300400000000000410c0000000100030310004100001330300000000c3d0c0000000fc000000000000100c3000040000c0431cc30000100000400040000000c1300c00540d1c3031cd00000000001000400000005400300000300004500c0d0c0000d00010300010000000d0c00c0000c0400010011000300003001df10c000004000400000400140041000030f00037001c1000500c004700000400101000cc00000c0400001c001004000000c000d30100300030c0f00030c7000000004000400400000000003010100004000000c0000c003c01000070000cc000004000000c0400000430c01d103040c03004c300000c0c10013101003000c000f100000c1730300c0000441007300000300cc0c3340c1000f00c001c000000000010c4000031010000000010c100f30004c01000043733004cc0c00010004c0000007000c10d00000000400100c43000010330c70000c147c0403000c0000004000c0030000403100c040000344000c00034300030040101544c300c10313400305040000c10c000500044c0000000000000f03100c1003400000c000000000000001010000000c000c0000400c00014000100c0000000100c400100310000c103000d04003054c0043100500000103000c430fc30100040004c000c0c0004301000004c000000cc140c0000004000c0cc50c00000f00c00300c043400013c007c003c0000c1cc101000000000000000c3c400000404c0d000005c000030c0000c1c1170003c000c00000030100000003101000c34043400000000000c000010000c40dc0000407000300400cc3003000000000000000000041000100000105040000c0030103030000c000004000040000001004000000000f00030c300400000000000000110c00110000c040000004c0100000c0c000043c030c0000001010000000100030cc0000001d0301000000034d0400010000001003000c0000d3000001c00000000000004305004f40000f030370305000040000410c700004031cc0000400c00003040000c5034c0000000300c007440f00030000400040030040c00040100c01000305c1c000000c000c113003c00040054030110500c000030f004003000c4100c000005110000050001000000101400000c00f0000040000000c010400100000030c0000d040007035000004000040000040c00000004000000005001070000c0004004040000010000000004;
rom_uints[763] = 8192'h374c000003300431c000000003000c0c314c000d0100000000440000c00d04101c41137130f0000000f400300100c30334040005d10c000d00300c0c10400010000000301010c01400000711300047c131300f100f0400000c5444400300310000314035005100c1c0007700300317000f71000310c0fc47303400d4000000000001043004340000000c00403004c0540c10400000030050100300040000c400c0c300010057300130113c1101040404000143000000031010c00000004c40000c4400c4400004001d10c0d40313303c00000704031004730f40001f00d7c0c0073010010c10c100003000c53c0100c040053c710101000c0000000d00040030011100000000c0c5000403004430004c40c50000034f40030dc00000c41f000003c000003d3d400100c000000cfc0f4c0c0f50d300000c00101000500f00001c1c0dc0040005000c4c033c0010010430153d000030d3043411000450300cc34c00100130f3f00c400c3104114110403000c004010403c00c001110070300330041c404003d1d400c0130c01040003000100003000000034c4043001c0c003000040003441300014300303f0c00010401c0400004304403004000704040100003d10000c00003300010100000cd00dc01f0000c010440103c0003300004c000000031c010000340c0000000d0300100c33030c00f3004f0001010000004334cd0051000030330140c0340000430041000f51c00030003d030053030010300410000cf4c00f03443400000d341700c0c7300403000030030300c304000340000004c04001c0c0000343c001043040c3030cc3007000040001040c10c0000014070000300cc0403100300003100d0000000000c7000003010000013013c0000c000034700000c0c00003c30330304d0ff00007c0000000c0040400003000000003001700300441c40300c00c030004000c1c300300d100c0003100000c01f001000c00000430000000400d0c0100f5003300004430100000070c030001000c0400004000d10c540000cc010001100314000400400c00013f3010001000040000300010010000f31404c30c0031d00300070c00040400c300004040c000010c003c0351400100700004130c0044c0c1435000000001430300001001c003c110c30000c131f003c33000000153c0300c00100f300d1d340d00450cc3400000001cc00040cc0c00000000403400050440034103c30003003c01110500000c0c000744c401001411300140000445c540303004040c0170c000040000c01030040c5000073c07c00c0100030001001001710071300405030300030300c0043000014000c00000000310713c00004c031fc70004400050000001010000037130cc005000000c0000010001000100540403000010000000000c0c04c4f0304c00c0c030100;
rom_uints[764] = 8192'h40c00001c1c00010300c304001001c04cd0300040cc17d000c03130000000c101d550f37100f000d0d0d000741403500c1073f033000c04001330c0113010003000c0343000c04000c00000000000104c530010c000f0000c0070431300d00000c0433004304c01304f0103300c0000f3010000003070c0300535d31c70007cc4070030000000010040c0005300300034300000400100c030c7c000040030013003000134001000d13000314013001fd0c0701000000c1c03c0400010c300c7c1f1300010041000004010001010d10001c10101d10000040003f0d04c000430000030004001000071104007100f0000c001d13004703000000130f03c00100430c01000700011c07003100011cd400034f0dc0000c0ccc04c4010fc000340004403d0000031c00311000011313174014101f00400754000000000c00c00000f011c3f10030370000000c0d3f301f0d00c1000000000f0710c00434c401100c0c00c30304071300441f154017037c00c300010300000401033f34003403011c34c0301d000401dd100c300001040cc10000003000000003400c0000030000000c00000005010dc0cd0c0703000001010c3500110101c0400c11000507503005c3410c0413001000c50c00000000c00c000c050d000100ccc00c000c07c400f1c00000000430343403344110704000f001000001117001c003310c0000110cc10d4000c1c3030105c004400100f0340d00000144000000c10704d007000c0001010000c70000070000010f040000001c0307070c00000c0c0f04c4405107c403c0cc031c3107000300050c00000d41001000000c000c0000000c13001003400c0700000300000cf04001000ccc030000000f0100100013cc00001c5c1404c7000345003100c3010034100300004003010f00475c000c10c1c70007000000074510f3400500050c03040c00000cc00000134c3400000431030c03000f0c43010101110031030400340000000c30040000010010030c07001f470dd0104001010700000000004f0300c4000103131c000c0c0cc40304000c000370f1f10f074130031100301f101d03003100300c41003003703100000c04300c00000001000fc000411d00013c0100070000c50d00000100c0001741070140040001c0cc00003013040f01043030010c0c00c5000c00f4004100030c0c400000c0040f00c00f040100030300010d0001400003d0c4000001c4070100ccc43dc400340001000dcc30cc0004070c00071c0000030d00000c53004401300c0000004033001cc3003c010c0d13010d00c0cd000c01000100000001000040070400000001c000010fc00c0c04031003f01000010c340403040cc001000c000cc40010050c0c00100000310034440013300d00c0744f3307000000c341100313c050010c03030114030700;
rom_uints[765] = 8192'h30000014f1100300000000dc00cd003030cf100000000004003000030141000000303dc400000000cc0c0000000c0000100000000000f003000c0030000000c4053330041000310000030c3000c0001c43000c0070c003110070700c00000c000c001000000040030000030073340404000014f030010000044000c003400030074000001004000000070004000f3001c000000d3004000004003304400003000c50000c3033000004001013301c003303c0000300030c00010040401c00000010100000003c1013003100004cf1010704c4300400010cc0c30000501000000000000001000c000f401f4410c000300000010000100c00c0c3c030040041cc1014000100010100000014c04010000c4040100030070000d30403300f00c0c000003000c00000003c000000000c400000003c00f00c00000c0030003f00003100000400c00fc0003003030c403000744c0440c404000030000c44000100000c010410d0300c1174f003013000104f0003400030c07400003000000000000005c004003000c5f00c3040010030010000000c3000000c030000000030c100303040030000001000000c30400000304003c0040330110000c51000430c4f03303c00000000400303003007000d0003003034400000043c01c00c10cc340003c0d300001fd00303003cdc400000003000f1f000000000003c30c4000000000043c00000c00000000000010010000c000340c03c0310000010300000000000040c10001c0000cc000500000000013030000017301000000340c00c0000005004000000013003000040000000c00010010000000c4030000000004101000000440c010000300000000100013000000400030040d000f0033cc40010000000000030010310000000005031000000450c0c40304101700c00341030003000003c0000001c0000004100030005030000130001c400005000000101000c01003030300034000010030000100f330010000133040010030003000c330f0410004007100c40000000041001000003000007c00300000003c543000300000010000030400004000010cc07000303000000d000000000010030010003340040300004404003030000000000000000000010000434030c000400000000400f10d000010000c330c400010100040000003310003004030030f10f00c01000040010100003010104100043103000310400100310400450000011000000003c31300000c00305400000050000000000001000000030040d3cc000010c0c0c0000010cc000000000000010030c0000001001000c0c0c0300300c0c004010000cd0100300000040000003000000030f3300030c0010004000010c04300000010000000c0301000300010300000500003030001004001f01300c0100000000010140344000000303100;
rom_uints[766] = 8192'hd030004c30000c010010000100000003c00044000c0040000c00c0003030000014c000c300d044000400cc0410103c3fc0400030041cc13340000000c00000103040c4d0001000440000000c004400000040404000d00000000000344c740000c1c0040c001c0c000005300c3130453000440c0010c01f000c400c0004c01c00140cf0000300001000103030c0c00000001000c0000000fc4000037003000cc44030c000d04400003c000c000c00cc0000f740000010400000001c400c00000c040410c00001700014401450304003000470145000c500400c30330000300050cc0004001fc0140000003000005000cc030c00001000013c00c01f4cc0000c000f100000000010300c7000c533c03010c0400014d073400cf000c3c0000000400c30100003c00510045400c03304030000001000000000000004f1c4040dc0d0704f00003c00d04000c000001050000000d0001005d000c0000000c01010307c001f00dc00c000c4c030045c3c1c30400d3000300c00101401c40cf40004300340147c0cc3d0034c00000000f00030000000c04040c4100100c0c0d0007c0c044450000403c000000300d0000c400004001001300cf0cc10dc00c0c47cc0c0034040c00000c01001500400040000f00f43c40040f0300f4005f0000000c000d01000400410304000310404030000c40010000004000cc000104000c0400c0010410000c00000001cc04400453cccc00000017173000100004c0c00040400404c307040f0000000000c00c000000f003003d00000c0f400144f00c0c0000c003300004d0000c000000d03c30003cc00000000701330f0d040001c30003131000440000000d3c00000300010001c100400040000103434040004143043000000c701001040000104c3100010000030000004f03c0c4c00c04000f03c01400000003000441001303c70d00000c000003400c0c40c040000140c4044c04000401004400000000000c3030000cc00c0c00c0000c7c00030000031030cc11000700400000040504c000310c00000145044004000f01c00005000040000c003c000000c4040000c041c00c0f00034100c00001300300cc04000000000c000030c0001340000004070000030c04cc0003c00000040030c100fc000000040344044c000040f00c0c0000000300c410d0c3c0000c334000134100015d4f00010000003040040c00400040000000000004cc003c000000cf4d01000007440d00440c030c000400fc004000000000000d040cfc010000c1ccc00300c3000d0cc0040300000f0cc0000070000c0c000004000400d00000100400000000010c000300000300304500037c0c4301011010500c00dc001000000c00000d00cc410300c70300004400004000c00000f000d00100000c0000000000310c0000001001000004400000;
rom_uints[767] = 8192'h1c000000c000001100cf00f41000d30100000030400000c014000030033130c0c010c000100040c0f000c104c07cc31750304003003040335c3000100301100170000000030000c00010c00140f000041030070c0103c0d010c050301000000010c0c00000c40c0110100000000001300300053000400000c0d3401300000001045000c04000300400000000c0000f03c3000100403cc0530c00001d0c5000004c01d000c0f0c00000005410700040000300100001331000c001005000100040103000100004000003c0100040d440000110040010c0004c000000003c000101000000010000100000004000c01c004370371004100000040130130000013000043000407000c000000001d0050043103000100030c000d01010cc5cc300000130c0000300c01000003041004001003170105040030040f000000001101030030000d0c01010004cc03050d001c0c0005dc1f043350cd030030401003c00c000100040300510010040d0004030005000d01004030f000070d0011031307000301c0c3043003030004004c01040303034c01000000000000c000001c0400030001cc0100301000000f5003000f4107310c007d0004040700000cc0070103c0001100000c131000030f010007000000431143000c400c0000010030110c0c004c31043f0000013d003c03000c0f4000f4c040370f0f00410c0400040474014cc13000010300010000000d1c00c130000400030f0711010000030140301101003c030c0c034400000c0001050c000f3001c0c00300040044d005000010100041cc01004000331300000c030100cf03005c01400004003d00010300400c3c03010dc040130113044d0cc0001c311004501730470c3cc004f01d005c300107c00003010110c3000c4d030d3d0d0c00cc4300000c30010c0f00100105000c000000c00c01c10003c0340400000d0131044c0f010d0c004301c00f3c010140c031000000c000000000004114030000c1010d300c00000d0dc000c0010001074300c0cc00030700000c0343033500400004000c0003cc00000003000103000c0c0000105000000f0c003f0c000000000340003c0c04700c004010010d140101013ccd3c0400c003010c40000d04030400000333cc1105400c00414c0c5003030d000f00004003030400330c00f1003000c1330010c00704040034001004c004030401c0000303c300300c4300000000000dc00c000340000004441000000400010153001c0c03300003001f00010303000c00000c0000c00c0300000100f000004000101010070c0031005c001000000000000000000d000001303301710000030404000100c1000000d00c05000d0401c040c000430d00c70c340c1541011301c1000c41000c0d000047000500000c03044f350c0000c0030f000330300000330c001;
rom_uints[768] = 8192'h50000100500004130030c00044004404400000c04000100000100000f0103000000c0440f000c4010000c0400c001007405004040010001050000c00c000043000500330000000c00c70030000004140f010000030c000440300c0005400000040453000000cc00455400400011000000000050000cfc000110000341000005000300043dc00cc4cc0c000010000000c00cc00030004c300d0c01000440000f000400003c00000100000004ff0003040347040000cc445404000ccc050c000004040f00000500070000034c000f0c00300c000400010030010000040300c000100400000c000c030400c0100100050cc5070c0000000004000003c000001c00c01c04300cc3041001400000000000000f001c0c0c05040000040cc04d040000004c0004000c040c004000000404010000051d0c0c0d0d000c05553100440c0000040f0000cc000c0c0005cc0000cc03040d001040041c54000340014000000440000001f354000c00000300050444040000000c034100000c05000000000000000f0004000000000c00050cc04c0000000003000000001400000c0404c00504cc0044400000050cc0000004014fc00005000c0c05050000030c0000000407000500140004c033000454004000000004000300040dc10f0400050044030000000003c10000141410cc10000010000100000c0010c0000c01030100000000430000300c0504004404010c0000c500000c000300500304030000f04c04010c010f0c04010051040c0400030000000010005004000c0000010400010c04000403310400010000010005100c0c040c0004007d04c0340c040d000700010500540500c00440050c45c00000c051014001cc0000001000100000070010000001000300303c0404000014cd01070007c000030f050004010c0405000414000c000101f0001cc000044c0c0403c00003030703000c330400cc00100000000f00000f0000000000010000040c0400f003550f0300100410503000033300000101000c00010000003c0400c304000004340300004403010c000000000c00300004000030c400040cf00004304c00410f003c5003c0040401030100000040000f0007c000100100000040005000003000070c0d00005c000f000c0400430040cc004f0c40000c0404030403c40c030c00450053400c000cc00001001c0013050cc0000400c00010140c0c01fc00000000c000040c0f000c00004400040ccc0c00000d0500000403000c000554cc000c04c000040c01000300504000000c0404000c000c00050004013c00040c0c0000cc0400c0000001410cf0000004400300000000504000c013000c0f0d000040000c0c00f0540003000351000c0c0c0c43c0000703101004000403000401043f050400c455000d0c000001000c0cc0000001000000c0;
rom_uints[769] = 8192'h1000000033fc401c300000cc00030040c0400010000c0000004000000001500040104000303000300c0000007040c0f000100310000003703c1c00000010c030004430000000040000000c0400000c3fdc004000f00040000003103000fc00c0031000d0300000007000001000c0040000000050000035100c000000000000304000000000c000000000001010000000000030000c003043f00000000c0300003000700004fc0c1000f00f000010005040cf0000000c3000034001000010000c3cc000c00000300104500d0c0040000040507000030004310050004c00c000400530000001300000500000301000140010000c3c4c0000f010000040004000300031c00000014c3000f0300cc1000000c0f001000030c003c15000c0130cf0100000000054401010f0303c004043c00030100451001030f004040010c001404700d0703030c00000c0111041c013c0c000c00140000440d00050103000c0003000400017c000000410c030000300003c0000c0104000000000c0330000000000cc00f003000000400000000030c003431000003000001000000c00c00000341c1f40cf40000043340000c00000000c000000000f000000400130f00003000000000000003410010044100004000000104c3c04141431c4c00003000c003300400cc000101000000000c000400c00030c300034001c0040f0c00030004030f700001000000c000040004040000010003000030000100004003001100030030010000033c0c0c000300007d0d45000004003305000c30030300000f00000005040c40004000000003000c300000070004000f0000003004000c0100000100000000100000010000400003400f000010100000100003000003000c000001000030030cc3010400000040400700d0000c00000100400c00000000030500c0030100040cf0c300000c10000ccc000c00030d0000030030030000c70104000000400001000000000000040000045000000c00000040003500c10000133000c0105d030000000007000111c400001000310001100004030000000010f040300c400100000003010000000c33000003004c0100c000000c000000030c0140014c130500000000000500000000041500100c00001000011440c3010000400000040c04000470010000000300000100000703010000003051010000010001000050004100000c0105000304040511000001000400000004001001000000cc0c0500000110000307010000010105000003310c01004014000030011000044100000103000000000c0f0d0001cf00000004300000000000400c3000400040000000004c0c0cc01c00000001003400c0f00c0001000000010001000000140fc0c000000c04070540000040000003c00d0003100001000c0000005011000c0c04000001000d01;
rom_uints[770] = 8192'hd0100100c00c1000c000030000000340030000100000c0c0070040000001001001300000c00d000040001300003000000040004c0004000041000000c3d0030c00000040000030033c0000130040300040500000000010000400007003fc00001501104000c41c00c000100000000000c03011440000100000303000f0001000003000010400000100003044040000100011000000100004004000000000300000100c300030000030700003000000000000c07000c0040007040000000001d010000000300c0040301070000300c3001010000003f300000044000f000c00000c3100000003007000c73000400030001000000040000000000010000c000c000030f000030000300034000000ff0000cf0040c10000000040030000000000000040000030c10f00c0c010013040110000041000300c000030c0c0003300000400407000400000c310004000000c3c00130005043000c50000400100000000300110c000c0000007770000000000001cc03000103f400c004000031413030040000000300044010000030000000000400100c000000c00400000300000014030c030001100700000d00010000341040000c400044100f0000010010030003000000010000070d0003000000004000c300d40403f0000d0040c00c5c0010000c010c3000300000000011040003300c00000130000000000c040c000cf7c00c000004000073041d000010100c000000444500c00400000011000000010000031004000000000000000100040004000010010400c0000103000c00040c0404000000400c3000004000c300c00311000030cc0003000000000300000c300513000044300004000000cc1000000100310c04000000000c0000004000c00000030304000c000000000c0000030000040c05c001030100000c110000000c000300c00000c0000300030000000414000d0000000000f00400000c330010000c03010000000000000000c00000010010000000f00000074033000303c1000304004000000303c0030000000cc000000000000d1001001300000000010000000007000404000000001c000144c00000000c40000040010013000000040000000700d00001c000041c0045000000c407c000000000000004000c000004000000000300000000c000c000003400000001005c00c0040000000404003300030c33000031000c00cc1003030000000000031400000100030300000000100004004100430000c430000001300c000300030310c0000c000c0040000c000000400000040001703154000000000000070c0001000005000000000103000001000c0000040000340410040c0000010c3004000000c00000000c00000000000000000000000000000c07000001000400c000040000000040000400000403041000030104000;
rom_uints[771] = 8192'hc00000034000000004030c00000004410400000000030000c00500c00000001000740034700000010000000010000f010100400004000f0441000c0000000000003000030000000000000000000c50000100033c3003000000000c001010300cc000c11100300130310c0000030100300000d00043000100000053c0400004000000000000000400cc00010000000000000300000303000000000040000000004300000000000cc0000000003000130070410000000000000000003300c04c1000010000004000040000100010030300004000000100c013001000040000001000000003010000003000d30103d000c000000003000000000000000000000000000004000003000000000c0000000c110300100010000101004000300003c30040030030c0000030000305000000000300400000000300010003000500004030c0400501000000010044000fc100010004004000000505000010300030010003000000310000c0000070c0000047000303000003000000000000c0000100c0101000000040030300003100430000100000001000000340700c300000030041f070300000c00000000000000c000c00000000000040000000000001000101100000040040000331000000000001000044001000003000010040030014100003010000000030001000400300000000000300000300000000000000030c40000000001101000c0000010000400403000000c005c0000000f00400000340000010c000000070f100300000c00044000300003040000000000300330410000001010000c00030004c000100c300000000000000440303400f0c000004040400d03004400000c100c00300000403c000100303004000300f7040c0000000010000000040004000000330001103000000000c01300000000c0300000005100000000300000000cc00303000001000440000c0010000007000000000004400030300000310000d040030003100000300000000c00000c001001c01040300000000013010000c00034000000040c00000030000000040c0000300400000000000010c00000c4400040000114c000103003001001000000000000100000000010000c000000003000000050300001040000000000000000000000c0c3154003301004100c00000350c0000403010c0004003010000000010000f00cc0000000000000003c000000100030001100030000100010030000000003040000c04000003000403d00000c0000000005500c000000000d14003030301000100300047000c00400000000030c0000000001010010300000100010030c000000300013000100001000040000000000000000003c0400400010000001000400000c000d010000000000c00000000c000004500000030000100c0000000010001c100004000000000c0;
rom_uints[772] = 8192'h100304033041003c0003050000000c0000000f0c04c0000035c030514c4000000103051040000004000f1300034f3c41100104030c00c000000001400c000003041d0001040c0000003040000c34000000030c0f00000f00045c4404000cc00705cd30330304001d03cc0500000d14000c000033300c0700000c0c014340000007000000000000000c00000000034000400400003001004000000104400414000400040dc734040c00000005000000043cd00001000c500c00004c000f0000040004c00000cc00040000000000010c00030000000700c000c00130030005cc00000000cf0000004001044004000100400c100c04100f0c0c00040000000004004c000c044c040000000c04040000cc000000330c0300000f00040400030000000400000c0004004c050300040300030404000c010400004c0c000000040c03c00400000500400c000004c00003000c0100030000cd000000034d0c001000000c40010400040cc050000c0c07000c10000f000c0f40040c00c0000401000400c3c400000c0c0303c13c000c00000000000c00000003c00000000c0004004004000750000010040c0007001000004100030403030703c3040d03c410000000cf00c00040000703f00f00c0041001000104400c00003c00c000100c00000f1f03c000110004c30f0c0f03000c4003000c0c000c13000000000000000410034c0c00000c03c00001cc40000d000d00c4030030030000000c00033043030100101000014403c3000c000401440000000f000f040000000003c007030430c0040c000000100000040430040000300404010000041004cf0c000c0300000400030101040c040f000c000c01000c4300010003000d0c4001030c01000704000300c00003000c03400000c1000c0c4c440d00004cc4000c0004c0d00300000000000cc307cd00000c434000030c00041c041c00040c00000000000400040c00000c0300c00400000000000c00003300000103000000000000c30f00000d0450070c3004000100000c0403001700440307004003c00c0c040003000c000004030c0000010103000404040f13400000000c0c04000703000000000304071404007c01030401400004000004c0030300030c0000030c0c030c040c0c0010cc0403100040010d00040003030304000004050c3103000cc30000040030000c0000000000030730044400000000004c0c43000001000700070c30030c0110c0040c000d400007004000c00004c00000000f041000040100001c00000c030c0c001c0c4c0300040c0400cc0c000504440001040004030004c400410000000c0c00000c00004000000c000433310c0100c0c40300100300000c000003000000070001040fc000000d0f000c00f0000d03003c030100000030000f000003cd0000400cc40000400;
rom_uints[773] = 8192'h100c40c0400004005010000c01300410000fc01cc00000c0040045443c0004040ccc0100000400100010005c470004c0c430c0c01030040000100000c004100c3c00004c0c003000cd004000000c04c40c0400340000044004101c000000000c0cc4100400403100d00030000400000000c00400044000304c004004c0005010c03110300040301c00401c00044400000c000000c0100000100004fc300c000c00000c04f04c0000000030400000007f003000000300c4000070000010000ccc00000000040010100044cc000000041404000000000c3400141004fc00105050000010000000040040000030cc304cc104704400000c30040c3400000c000000000c744000000c3400004430000010d0000000c0c4300430043000001000c040000401400000045000041000000000c0c010003000000000c004000c4000c004040c0c000000c450107410000c0c0000100010000c44040030d40030c00004050000000400c030c0000000030404007c0000000010003c5010000430000cd00cc000400c0c0cc000c0400cc01c040004001c0000c0000c0040c000c1004c3040300cd030000010c00c00045c00000000000c000054301000041c000030cc0004040cf00c0c10100c000000000030003c0400000c0000000000c010100410000c3030040410004cc40414000410d030101c100c10001040400000000000000034100c00c0000c00001400000030100c30300400000cc04004034304c410044c04000010000040000c000004000400104cc000005000c01ccc00000001000c000f0c004c0410c00c700000c0c0000000000000033c30000c103c0c3c00d0c0d0000074000000000c34004c040040404c1c0035c000000004000034c0d00c0c0400011000004300010c30000ccc4040000c0040004000000400c00000145000cf300000300004400cf000d4000c3c04001000d0fcd010000c0411300cc013043c1040f0c000340000000000d0c00000004c1031c000cc1cf000000010044000c00c00f000003000001c000414000c040c400140100c000400000010cc001000300000000c000040d000000004000005400000000c0010c01c0000000c00043ccc400000401000000d100040000100000410040000104000c1000c0000c450c43000000c3c100000014000011010c0000000c000c3003c0c00003000c004001c0c00000cd040000004401004400400005000000007004000c030000c0000003c3000c000000c00140000000400c040704c340c1000370004d410700000040000cc103c3c300c40c000000400140000c00c00000c0000343000007003000c0400040000000c00140c00001c00c00000c0000000000400047c0c3010000030d0000c00000010c000040030c0c01001c000003c0000000410cc30404c000004000;
rom_uints[774] = 8192'h10000c0300000101010000303cc0c000000d04100400c0030001041140011100000000470d0d000304100004000003c04004001000000003000c03001700410000000010000c0300000000300000101c00303c101d01001c00347030000ff30400ccc00147000400c3400000000c141000000004333f0054000000c000c001000101000000100101000010000100001003300003000c01000010000000313400330300103000c034000000000400001c0004001000000c4300dd00003f003300000c0104000000100103010c3300000f000104000000003000001341015030cc000c0000010001000011003f41c30000101c011c0000000000000001001000003f000001cc0003c0000c100054100003007f0000c3c40c0000040003400f00040010330000000003003003000101511c0034103c100300000070110531030f000000000004030700050400000c000003001c303cc10400040001f13300000330003700301140c00c73300c043701000101001500c0010030041ccc3000403c0001041c0110000005334340300c000031000000000000cd00c4c00c44303010103301d10003000c00000000c0c010000000000000000d10004404003000000110011d1101001c03400040c00330013005cc00000000004f031001001500000000000c070303000131044000400041000010000050030401033304000144f000030c050c141030000000c00c4100000303000001c400017315001051000c000c03050300030001001000000301c30040010100010100110f03000105030000007034040400154001000000000c0043000c431000003330110011300530003031100304c10015100040c0030f1000001000010300003303c01100003c000300000000000311010010003310c03013000304404173111003007000c010400000c510003000001000030000c0003cc400104300000001050300000cf3010403003004000c030000000010000000010001330000010033043f000003c1013101000c4001004c040001003000d0000d0c3000331d00c0030c100000000300030c00300000000000000300010000300f0011030c03003c01031000c000041031331d41010f0f000c011000f00040c1c00003100000d0010c034f00000000010f040400013044000037000701000cc0000000400001f44000000f040014041d00003c000000003033030c0001c10011000700317730c00100cd005103071d00d0001300c3330d00000004000c3000000c0000000c0000000c03300000d11c1004300000300003051c14000433003c0000c00c004000000c050000030110440300100c040410001104000710c440070000400400000404040000040401c31c00c10000001f044f0000410c001100730d100c1041001f34c005000000001011041000010000;
rom_uints[775] = 8192'hc000041f000000404003000000400000000000c000c0000000000041005000004c00000440000dc0c0c0c04040c01000000000c00000c00000000000000000000400400440c0c000000000000400c00010000c40000000440f000c0000000000000000100000400000000003404100000003c50400000007cc0000cd00000041400000400000000040000cc0000010000000000000000333500000003c0400c0c000000000c00004c0000000400410000000000000004000000000304000400c00000000034040000000c0000010c000015000000010040c00004040c0030000400000000140000130030040c0c000000f30100000000000c00000c00001404007000040000100000050c0c4c000000c00001000c00010001000030040c0c000000000400000c0400000c000004000000000000000000000404100400000000001000003f000001000004000c000c0c00c4043c100000c00000c40410100000c40c00d000000d040c00000004c0100040003c4000300c00300400000000000c00000004004000400000000000000304000c0000000000c0c40440000000100004c400000000000000000c000010000300000c0c00000d0000d000000c100c004440000c0030000000c0001c0000030400000c000430dc0c300000000c1c0c0000cc0000c30040000d0d000000000040000c0000000000000c0400ccc00000000401000000001c0c00400d000004000000000c000403000d000400cc000000000014000c000000000003000d0004000000cc00000030400c0c000000000c0400000c000440c00000000000000c00400000c000000000000c1000000f000000c0c0000040000030000030000010000430000c40000000c000050000000400000000000040003000401d000404000003000000000010cc10000000000000001c0c00044d00000300000000000c040c40010c0000000c0400040c007c0000041c0c000000000000000000003c0014003000040cc3004000003f0c00040000000000000000000000cc0ccc000000c00400400004c00000000c000c0c00c01000000c04cc0cc0c0000c0500004000000405d00c00000000000000040000000030001c01300000000c0000040000000004004000000000400004000100030000c1000000040004000c00c000300400001040000000000c0c0040043c0000000000000000c00000c0000000000000c400004c000cc000044c100c000c0000000400140400040c0000c0000c0044000c001010c0c000000c000000c0000000400000000c0c000300000000000c00011000000c005400000c000000000000000100c000400c0c0c000c3304000c4030000c30001400000004300047004000000c30000000000000000c0000100034000004004000000c0400c0cd00040c000400004000;
rom_uints[776] = 8192'hcc0400401c000000000c3010000c0000107410004010000c001440000010c3304c0040100400000000001cd0040000000cc03000000000100400000010fd400f0000004000300c4c003f0004103040101c7c300c1000000000c0c0001000d11000100000001100000410000040401000cc1300000034001104000003544000047000c000400000c030001010000000000070000cc0430000300c0000d000040c43c03c00400004303000040007c03000303030001030403300cc0c0c44340000003000001000000100110010c01d10d00000000040130c7007c0440000003410003000000000300133000010703050041c00400000cc300000000c300000030033101000430000000030000cc000100c100004031c0030cc7c10050000c000c00000040000000000001c00c000000c03300c003000440c0c0010000000000d0000100000000000001030c010000c00101500d4dc004c0c5040140030010030f01014003010300c0c00040030000014003030000c3040c00000403054d0400031c0000000101000400010c030001c1000004c000070000034103000004130000010000010c00304003010001000300000041cd0c0000c00005004003040000400404010040301001400c0f00000000000cc40d000000400111004000c00c40300000470040030d014543c004d00000c441400c03c440000c0000000010013100000300c00c400043c34000c000cc00010100000000010100300001004150d0000c00040000c0003000000003f0c3400c030000010fcc0cc0000000000011000000c000c0dfc00fc000000041014040400004000100030303000000301000037107010400010500030000c000030500010300004000c3030100000007c0010001000000300c00040040013f00cd730030c00001000d0100000c00000cc000c404c300000007003ccc04c0d0010005c00c03c4010001000040070000c300034000c00001000100c000000300000000000cc00300c04403001cc00c000c000104100d0c00000f01000003000001c00c0001000c00000303000335030100540cc000030000010001030f053001c04000c00001400fcd4c100c00300000000100000330400000000000000004c000000c00c00000400100c0070f0110004003403000c00003000743100f0000000d300700000000c0030c070000304100400003d44703c001100400000d300cc10c000000c33004010c0443000347404001000010010000c0c0030c03d0030004000000c000040d0000c0cf40030540000005fd40400000304400000000c1000d000000000c0000000c010000010400704010030cc000c1c00001000cc0004001000000010400c00c003041c00cc000c00c034c0000000000300000c0010040400430000000000c0000000c04000c03000;
rom_uints[777] = 8192'h330000300014c0331004000000401000100000300000c010003000000440000000004c00005000000004000001100000303000000c1000303000100000300700000c101000003000000000000c004000c430000013404030c0000410301c0c00000003c00000100000d0150c0000100000103030107c003000000c000011c0003c1004000004301000d00000000013000001000000004000000000301000340c00000000010004c0005000c73030000400005400003040110000000000003c000000000000000000000103f400140000000001301040000000003030c300000000100000000000100c1000c0100c0000000070000000000000000000fc00001000000000100000040000001000003000000c00404c3c04001c300cc00051103030500000003000c01c001c00000000040c30001000000000d0001410103000001000000c40c3c00040000010c03000301c3f005d0050003400c03710101100000000001430000030d134000c000040130000100030000c00700000000000100003001010000000300000000001000c340000003000303c0010000000300c00500010000010f30000000000300000004c300400313000003cc0010000000040303c0030000c0000330000100000103000c00000000c10010300000000000c04700000c000000000403000003700030000100c0000003030500010100034000040c0103000000040000004000000101010000000300300c4003000400431100130010000000004300000003030300000000010300000000c3030300030000000003000303001300040000000411000000c001000003000103030c0000000000100004c0c1000000033300c005010005010300400011000000010d0c0003c0c0000000c00003000000400003000100004001030000040000400004000001000d0007c001000300000000000000c0000100000310000000c00040c00033300001000000031000000c00040000000001430300000000000003330030000100030300030000010300c003300301000000000300000000000000040030400000c100000f00000003c000031000000101000100c000000000000300c001000000100001010340010c040001000000c0000c0100000000000300000000010100041500000000f1000100c003000c030111004110000410000003010101c000030000030300030100000000000000000014c400c00300000114c3510000000000000000001010010c3000000003f30044100001010000030c0101041000c0000301000400040003c00043040c4003000000040303000003014c400000c0000000000003330000100000c3010100000001000143030000470000000000000330c0030000040003000c33000000c0031c00000000000000000000000f31010104c00000000c0;
rom_uints[778] = 8192'hc000000000001000000000000100010400000000000004000c000c0140004000c40001010dc0000000c00100000000000040c00000004040c0000000c0000005000c4000040001000000c1000000400c0040010f000c0000c00000000004000003000005000000100004000011004100010100000000014004c003000003000000c000c3000000c00100000c00000040000001000400030000000000000300c00040400300000c000d0000000000040400c00000000000400300000000000001000000000000000000cc0300040100400000000403000500c100000004c000000000000000cc000100000400000000000001004000000001000001000000000400c00100004c000001c00000000001000300000001000000c000040443030c000c03000000c000400004400000000004cc000000000000040100000000000000c0000c000104c00100004001310400000000000c03070003000004000000000000000000000000000c00010f00000000010000c0c4c000000000104c00004000004f00000000040500000400000013400000c0030001c0000c000d0100c0f00040c30000000000000000000c00c0000c40000c000000000000000000040300004000040000050c000400000000040c000000000000014401000000c040040000000000400000000000030040400000c000000400000101000000000cc40000c3400000000000040004000003004c000c0c00010001c0000100c300100c0003040100000001000000000000000000000070c000c100004104040000c0000003c003070cc000000000000004c0004000000c0000100400000003c10100c00c00000000000300c000000000000000000000000000000300000300c00003000c00c000400000000000000300000f00010c00010000cc00000300000000000000010000000c00000000000000c00000c004c00000c3000000100000c0000045000cc040004000000000000000010000000000000500c300000000000030000100010cc00c0003300300c00000c0000300000000000140000000000000000cc100000000000040000000c00000400100040000400030044000000000000303c0c00f0000000000003000300430000000000000040307000100400000400000010000074c000000c0000000004c000300c4c000c00000730100000000000001070300c000000010000000c0000004c0000000010001013003000005410000000c0001010c000440c000000c0300000000c00000c0030003000c0004c0000000000000000000000003000000000044040100004000004001c0000000000000000000c030c04000000000430000404000040000000c0000000000000001040f0c000000004400000000000000000000000c000000310000000000430c000000400000004;
rom_uints[779] = 8192'hc0000000000000000000010000f00c000c000c0104d0000003000400040000000003040040000c030000034001000000000000c100051000004004000000000001400000000400400000040000c0004400014c33000c00c000c30000040d00000001004000000000070000030000000c00000c40040011000001c000040000004000000000010040000000000000004000000000000c3010000004430000000110000000001010000c00000000000000000000000000c300000c13000000010000000c00003c0000000404c000400000c044040c00000000000000c00000000c000c000000000000c000d000c00000401000000000030040000000040000330404000000400000040001000c0000000c04044c0100000cf0400000d30c0d100d500001000000000000010f00000c00000000000000000000004000c000000c000000fc400000000000030f0000040000000000010001010014000000000004000c1d0043000040000c000c00040000000004400000c0000400c0000000000005030000000000040100000000cc300c000000000000000c30cc000400c00004c44001000000000000000d0005000000000000d400000000050c0003000003000040c3040003000000403000c00c001004c0000000000001030000003c4000400001000c00c03000000000440700000c5000040000000304011000000000c0011c0f000000000d0000000001c000000000000c04000cc00400000c000000400c4d00000000400070000700040000000000040000000300004010000c00000c0000c004000c000000cc0c000c00000000000000000000000000000000c00000000000c00400000401004000030400100301000040000000000000000300c000000c000000000000c00c00000400004000000000000000c0000c340000300000400c00004c00000301010000010000000c00c000c0000c000300003000000000c000000000c0000000000000000000000000000c0000034000040cc3c000100001000030000000000000000000000c000000000100000c000004010400000000000000cc00cc00000440000c0003000000000000000440000004100000030000040040000c100000000000000cc00400000c0000000c000c44000000000003000004cc0000001100000010030040000000000000c00cc0000001c0000000cc000000010c000000000c00000400c00c000000000c00000c40000c0001000000000010010c00000000000000000300c00000c00000cc0c00000000001c00007000040101000c4400000000100044c0030030000001000000000c0040000000010000440d00000c000000000c0000000000000000000004000000004100000000040013000000000000300003c000000000004000000004000004050c00000000000;
rom_uints[780] = 8192'h1001000004d00c3000011010fc00330000003001000000014003f1040300004030f000000004001000030000014003400010000333000c00040c00004000c00f313400000000000330054c050034050000c4040c04040000f000000c040031000431c0070010c440d0c001c300c10c3001d00401304c0d1000c00300010430300030030000010000004013000d000c00030000040d0100f0040000030000000f1300000111c0040c041100100dc00000d03003004cc00400000c05300000040000140300310000c00f0000c300000000c1000004000cc00101400c000c00000000030000000400fc0000cfc1001500c70405c1400000c030c30030003000000100000005cc00c001040044c000034c40341300003404340000100070c01000000004003000c030100070000000030010000034000000430c000d4340300f4400cc00001130004000033000000000000030c01c43000100000004030c3c30dc310c130000050030104d303c03300001c7040400c00000050c0f30004d30040f0050044030c000053c0000300c433000000400100400000c0401010f04100ccc301003000000100c1405d000d30c4000000334054000cc10051c4c100431000004000c000000300000c0104070c00c0c0004005003cf0110000030114000051400c0c001001cf04441000000100f013304070c000c0c0000000400101c313000010030000043340100c40300100c00034001c4c0001000c400c00000403000040c0000c00005100c0d0404c0000004010300013000010000c00000f0041f730000c000c410000000c40000004001000000100000003000000000030c4000001444000400300004040c333c000130c3d0100105000cc0c300cc001000c1004d007004010044c3010104010fc0000741054c0400004f0300004300004004000cc00001344330500c000c0010f0000000010d30000c44000c400005010cd0303c00000d7000000000300004003000000000040c0c7100007344004001000040000000400f34000000300100f0c0c100043f0331c01000000100013000034430000003000f10044000400000c0040001000004003c0000010100100c010c0000440c000000000300d010040000000c300000010c000004040341000c0414140000c030040c000010001110000030004000000000000cfcccf037030000003440110000cc0c4000055000000c007001000000000004000403001000000ccf04c0c0c0103010000300c41410300003000c000000000f070c73103033000c4400033000340301c00f000c00003000000000040040070100000003030070050304003004010400000030000c0dc40003c00f0ccc5000000c300300010400300414003713000000004000003300c4000033100140000440100010007cc00400000004c;
rom_uints[781] = 8192'h10000000000040000cc00c0c00130013c030014341045000010d000c05300000000d07c34d000000010014cf040003011410000030100430100c0000f0000c03003ccc00000040d00000000000001300103404003c0130005f050c0000cc100000040401000004000143c000010737000030030c0f0101000cc03000c40d0000c4c031100000000d000000004004410100010000000040043030700c0c011030000010010400043c030000400100000000330700000005300d00010001c00000004300000003000014c00010140001040330c0000c3c00330c33c00003400000c03000040f0000030400400001dc0c11c50411001f3000000003000000000130000000f1300cc340033003030c0004000001037f01030003c3c0000005000000000000000100c00004040000000c010400000001150033000030100fc1000000000000303000300000040100400003300d403c0300c0001000040000000003000400001001000dc0000c0c00d404170000000310dc01104c03000c0000000004030140c1001000000001000040003700c00c100000000000010411000000010101100c0303410c00000cc00000d031000c40040c0c0001031033000003003040330c0001000010040cc40007030000111000300c00014001014000000c311130000403411c0300c000000d10000d0000000003010400000007000031d000000050070003001100001003030000050c0f0400141100340000033c00000103c413001c00d00cc01c0000000103000031000f3500040c30000001000000000011c000070000c010000010c00c0000003011010410c0010001000000001000070340401f0411d0c0001003004f30c0000700100000000c00000051c0000d0c00010c03030010040000030003404003030000004c0000033000f00301000dc100000300000001004330000000000403000d00000c300c033000104000001403100030c00301c0100001010000000010000000000000710030000004000000040c1c0010000004100c0000430c0c00c04000030d00100f000000000005c00000000000100300033100003030000030003000041c10000001100330100c00130c30000100c000000304170000040307010000000fc300000405000400d0f10c070003010300cc01033030000000000300000000000500041470c0c1d0050004c401500030000005000400d000030400c00c1004c00300100010001440d00100c5c3100000004410000c0c041300000010010001115001100000000100010004c0c00100100000001100c0430003000400000100010000001003d103010100040404014c004f310f010c3300000070000000000401d0000000100c0000000000300030000311000000400dc101330000110400004000000c00003000003c00c01000040;
rom_uints[782] = 8192'h440100000430000100000c00cc00001000040100030301000c03400000000000041040000cf0000c01000c0c000004334f44c10004c101c0000c01034dc30000000000c00400010000030000000000c0110403000d430f040003c0300430030cc000cd31400c00000043cc00400d40cc10c00001400440400003400010330000050fc1000004441043000000004040004f00000004000000c00f0103730303000c3000000000c4040c00000c40000100c01c0000004730400100c0030100000c0100000000003000000005000000c0c00300000000000730c3010003c10005000430cc04001000000c000c300000040000f31c000000000343000410000000103000040001c00c000034330c45101c000c000d040030c040cd00440c0f30004c0104000000000c30000100c0000d000000000000c010040003000034000c004000000430c70004000c3035c00000004c4d400000001307010403c13000110003000404100040c01010000c03000000c0010000010000f0000133f00c000000003c40c0035c00000cc0c4410c00010cd1000043000000c0c1cc010500030000014ccf100c0000000003140000010c000c00000000010000431001c0000c013001c10c0401400000000005f000c0c00f1007c000000000000000c03c050c03c000030010000004c0c00004054003400c00000031c000000000070040000033cc04000c404c0103000c0100000000010043010417000000f0050000100c3004c00010fc4003010000000003400c0c030100043cc00100cc7400ccc41015000c0010c04010c0000c04cf45c140c0004000304d0c0700000000c103c000000000fc000c40044f43100000000070000000c30340004101404330001400030300c00cc4c001400300040d040043f40104000341c0c3570000103d0400404c01010000001013c00000000400000fc400000700410cc400000c000500c00c000c4040000000003000000003040000030004c00000070700000003043f00c0000404c0000300000000c100c30c0401000000c00000000c00414000d000000d00000040c000400000000fc00ccc00014400c0c0000d040c0003c3004cccc0d0c1030f04030c0140000700c44000000000c00007c00000000103000c000c440003000dcc0cc10c0c000300003040000c040d400410400c00c00c04340403c404c004001000000c0c10100100040f0c003000500734040000300000c040000000000000410c03100c10d70000c00f4c00000000130110000300030013000c0c0f030c1000000cc101cc400000000000f000000000004000c00000100000010440000300000c000000000cc04040400100000000500000030c0100c310000c0030c300400100001040000400104c003000000000030404000000000001c003100c40000000001;
rom_uints[783] = 8192'h300000cfd0c40003000c050000c00010000000000d3000030c00003005400000c00c40030000000031000000010001500040000c0007d00000007170434c001cc004c01c01000000003004400c0100405c10137301001140304f00c333c7001c303f7000000000cf0c43cc00004701001300400003104345c3c57300d000070330000cc300000007d303004000003c00000010000100000000704c100010010c4d0001701104400001c40004040330141040c00100d40c00000133d30c0010000c00c00000c100004430034040704000c100400c00030307c040403300300000c0400c00100004404001740030000030c000000040c30040c1050c4000031c3c0c0405413005400300300040000c0700350010300d3000c14003d00000c40000440000031000000000000005030c00017cc403400c0c0100100437004130054301000003100307000003c3104c0c101000000014004075000434501110030000000303c10000050054d00301c30400040700110310c1000311043000071000170c700000030040114000330003030000000301000010103f000340000300400000300000710c0000000031070100cc0010000413100300c1000c00000040045511030f000d0f40404c000040011400400004001033d00004010c0040010300000040050000030303003c00004000030001000011400fd00400033100410d00701c005c0341c0031050000c70041c101004d000431c3000040100001c014140300400001f0143040030040c11000000c33dc000000110c041c4c04000000010403000401001c000340003c00d00300c00114403300304005c04cf100cc0030c0100000174004000000001c3c0004000301f000c7f351000040cc7c000003003c100000c000400c00c410300000301010c1c40c300400100000f400c00004001c103000311431000400004c0331037040f0f01341f030c701040000c00100d00f040d005000c000000100000430100000000100030003f000053003c30000000000c0001300c300000c00350014010000000000dc000000c0511000c0010000340010000c0c0c03100000033030300c00c10c430000000c10430003c0003000111700010c00c050001c4000c000310030003d43f1044030103f000c043010001004005d0000000000000410cc0140000000d003100c00405474000000c304f000c1005030000010070000000c30033000003430001430173000c053030000004304037004001110040004000400000c000050c41304000c3dc0530100f00010c004300c100050000500c0010c0010d710001001c7003040000000000c71040004003c303c0103030300300d104014000750c0000000304004304400100431fd00c0001000c000c3000cd000f40004003000000010000cfc4050100000000000;
rom_uints[784] = 8192'h4000300000c04c00040000f0c00004c040c000c0005140000004c0000000c000f0000c50c4c0000050cc001030000004c010c00030005c40c000004c00c00400c05114c000f044004000c04000c30000c000c000c0000430000010300040c000040c7cf400f004c000003040040000005000004000c400000000c00000f0000cc0100000000000c400f0003c40404005004000000030000140f030000c4000c1fc4000044000f00400004010000000000040c0c000400c500000040050c04000000000c010040cfc10c000c0f004cc000c4000300000c0c000004000404000000400000000c3000000100c3000c05440c40010304cf0500040400150c000040000c004000c00f003003000c0000000040c101034c00c5000000030f0400c00dc0000c000c40000000c400040000000c40040c00c0000303030401010000030001c004000003d0000c00c04d00000000040c40414003004000c404c400050f00000000000000c0000500030400c00c040000000001c00000c004c04000400c4005040f044d00000c030700000004c010000000ccc00000000c0c0000000c0c40004f0c00c00c400400000c0000c0050040000c0c0fcc0c4c0000000000c0050004040c00000c01050c010700c4c000040000030000c4000c004d00000000010f0c00100000000c010ccc00000000000c4000cfc440004003000000004d041000040c000c00cc0005000f0c0000004c000404000000000000000040c0cc030c00040040c00000004f0000400cccc0000c00000c000404040c04144c0cc000000d00010000000530030101004cc000000000000c000c410000ccc5000000040004c00000004c01030c000c004c41000c00000fc000004c0c030d430c000c000cc00cc4c4c4000000c140100007c4000c00c0c0040c040300c4000f00000000cf000c044f000c00130004c4003400005c040c010c000000000004000c0c0c0000c00400cc00000000434001000404000000000c40000c030001c400044c3000000c40000c0000000000000c000c00050c040c000053034f000003000007010030000004cc04000000c50c000300001c0000044000000000c4000c010000f0c00c4c0f00000000004000000100c00000000001c0000003404105004c0f0c00cf1f0c400f0c0c01040000000701000004000000c310c0c1000c0fc401400000c0050c030005040400000cc0c000010103410041401c4000c00504074c00c00400c50c0300030000000001450000cc00004000004000c10000c1000fc50000004cc00100c4c040000001c304030400c0004400000003cdcc004c00c0004000000000004cc0000c0f454f000cc0004c000100000001000d00010000030300010001004f04040c000001000f000000c001050000c00cc000000300040005000300000000;
rom_uints[785] = 8192'h1000003000000000103030d3001050f1007040000070000000c0303000301000303000000000003000003000f0105000c01000100000c110000000000130c0c04000c0000000101030c00000c00033101030c1103000d000100010c01010007000103000c00000704000c000c0c050700011c0001000000030c000d030303030d00140000000000000001000c000300000c0001000c0000000000070c000300030004000c040500000103000300000000000d00030000000d01000000000401000001040400000c00031300000000000f0100000c001f0003000700040000000005010003000d030000000d04300300030000000304070d010000010c010400070000000000000001000003130000000c0100030100010100030403100700000000000c0304010000010c010000000c000100000d0000030c0000030d00030301000000030000000001010f000303000c04040c010011030c0000050000000100070d000000000400000c00000500010c00010104000001000f01030001010d0103050100030300030c000000000d00040d00000c050d01070100050300030505000c00000105000100030c0d00010f0d0c0c0001010000030110000300030f0107000101070000000d05070000000100030701040000000303010403040003000f01000100000300000010000c010303000f000000030401000c0501001103000400010000030c00000000030300050100010000010504030004030000030c0d000100030003010c00000004000000050c000c0000001000000c1d0304010101030400000d00000c00040c0f140000000301000f010103030000000001030d0301030100010030001d00030530010130030400030c000301040001000c010c01011c01030103030100000c0c0f05000100000007000c0c01050000000000010100010d00000100000003040f00000d0f000500010f000c0003050007010f00000d000000000000011103000700000307010c0000010300040101000004000d040d030005010400000000000003000101010000000100040c010c00030003030000030f000315000d07000100000000000000001100031c00000f00000000040400050403010300000f0000030d030005010103000703050100000400010003030100000001040c0c03040000000c0c00000101050000010f0c0d00000c03030000003c03010003030400070301000d0c00000501000000030007000703000100000310000100000c03030c0f0000070300030c0c03010c300003000000030c0000000001000103000303000f000c0d00030700030300040c010104000305010c030701000001000404000004000003030c00040001000000000f040000010003000d0400000f040c01000c0c00000300030f0000030103000000;
rom_uints[786] = 8192'hc00100000030100030f04010111004130000330100f0c300004003300171000043303050d040c04030000000030031f0000030400001700003300000f3031000c13001113310c3c000000000000041c0103503401044014030000430007100c34011001731000000400004000100c410000031d000f0450001fc10300113f0000344014030f0000000400000000010c000000013003000000034104000c0000051011c000040f5c111100000003003000150141000034300001000003040f130c011100000010c301000000030134044430135301440d400c3314030c11c31104040100010100c000030103d00000000313c304301c1005000010100000000f0c101d30f313141c00010313001000041340d5050004004100304000c3c40c0004030700000700310c04000003000c044c001d374503000c0c000430031000400f003f13540c3d000330070300000d003f010f00000450074f13040c070000110c13100f0000010703001000031000333c100374003030310c05013300033040043c310f0f1105100014111105003c0c33c00000100000100405d000000003004dc00000100c050c0010003413040010030c010301130f401104030003000471000400030000c104000cf443000c4000000c00040d40010010100004001304030000010004000100040700040d03000c003317030010401f11003300031341030f00400710000000000010000c10041c7f0c04001004403004103300310004040c040d100c00530004000d00303303000d03500c0010c14c010c0300001100d7140000400704300010030000000f10013c47013000030007040300010d000001300000000f730001331c010c00301030c000003000030331000304c0031d0c000c0c070c0c04000d000d100d1dc304030310533307030347500c0140000c1c04031133050000000c0c04107170400c330440100010033703000000c03000000f101400010c000c0013c0400000000031010050111004030c1d3403cc03000040003001040310400011000000400c000005040004111d3304000500040c13000000f0c1031d030001000c0c001c0700010300000700010030100000001515000c05040c000fc4030044001305040410013c001d33d40c00030404050c30004f043010c33100030f00000ccc100f0714451737100c030100173043000401000f150014cc010003000c1c00003133300c1017104040000c5440070030031013c037000c000003000000700030100c300000040000103300304304340c40003303000f040100f5000441f0040005010c000c4011d4003d00004030440000000033000004010c00044000110010013000040340000040040c1c00503000001c0d000003053000340000f311400c04000c34300000010431400c000010c303030030000;
rom_uints[787] = 8192'h400000000c0cc11f00040c10040cdc0df0c00c05c1440100000c04c004c000000700045ccfc035014340041f010c0d3044013304007400f000c000404004000c054c01050c004c73000cc000c04cc10c41000c30f4044004000050f004c303100f301c014c004c0004cc4400030c50000030344c00010c0c404c00000c0000c00143100070f00f0005f0013c000100c00000001000040300c004cc41cf000c1000c44c00017f7c000004010404000000c4dddfc00710c0c401c0010330040001434000d0000c11c007440c0040040d05fcf1304101cc1040003401374700000010c000000040000000040073d34c0c0000350df13cc400000c0c01030c0040c3c00cf01d4cc0004010000c3c03c3044005040010053c00001cc0030000000c010130000004cc1c0000140cc000000c3000500040c0c4fc0cf00030c14004c04070010c0040c0c00c3001d7c0004004004c0140000d401010440000000300400000c00300c40c1000004fc033100000030c10c07040c004404f1443000f4cc0010c44303033300c00414000c000005303c000c0300000f000040404300010c04001300000cc0003000453100401c414f04000010f40000c031104000000400401040c001400f0404000000001cc0000d00c530cf0000011400c1000034050000c100c50c0000cc3040d4ff140004c0c000c0d044c04400004c11cc000540000004cc000401000c0c0cd0040003301d00c4443d00c40040401c004f0001c703010010400004c004cfcc000700000c00cc0c300040c00d3400000c01040400303100c4c1004000c000003000033043000c04c44400010c0333104001c03000403100050034c4c430f40300100c400c5f100044000000c000c01cc40d01c004003000c00007000000c000304cc3c07304c304d0470ccc5000050000c0000cc00c0010450c403100000c4343000c0143f10010000044cc1040304c000404000000000040dc0000000f100f01404004f03000000c4040311c3004000c0c00000c0300cd0003345f007004c00c000000330c000000001c10cc0000ccc4000070d04005044401c4753504441000c4401c1cf04001000100000044cc010000040004f00cc00300040c00c0cd00000c0041c00300000c0fc400000000d100c473000104c1dfcc00000010443044f33700304f000000114000c070c1c304c00c33404040701100010d4700000500c00c440000f0c00dc0143000000f4400df005c0030041001c11c000400c43c130000c000000013001c0c744104c0001f003000cc0c0400c304dd0c0410cc74400000c0100300070010c0d107c000000c000000c0000000000c0c340104c4d100040fc004d100f004014c000030f003100c0c010c400100f1400c00034040c00cc00c00c00004004300404c0400c0c000000510c0007300;
rom_uints[788] = 8192'h70c000000c43c100d0c0c0443c4400d0100f0c010301c010c03fd000000005000000d07104130000c1c000414310410700010100cc0fc0300004c0c0c530c11043010c0040c03030000000440400000035f4000103700c30000371c400010000c00413c0d04000005c0101010010dc0000307001d330003100000000c400030040cdff00004000c000430000070100070504c0f000000cc00011000010000c0040040c34d00d400700c0333004f3c01400000340000400c0050300c100000040d0fcc040000113014113001037c0000000c31c00000cc0c3030045dcf4440001030040000030130000400000c00c0c0c000071c05ccf00000f0c400034010043170000dc001300f100c00f000150c000040dc0005330100101050473011c00000005c000400004000f004004030c00004000030f300dcc0000007c13c0400000cc401303d00431c073c4435c0330400040c400d007150034cd00f0050ccc31c34013c10000c00070cc300330104c1000c0c4c13443440003000000000003c300f444c0410003c0003434c100300000005c00037400007040030310700cc0730004d000000030c0330070334c4070c1c10400000005000030300030c00001c034c03500003000004000c00c000d003034c0040440000cd33000c10040c13470403000010d0310c001313400d40000030334004310f000c00040c510100d40000cd441c041030000034047c3c0d00000000400cc40010c0001000010033300c11000411ccd004330030000c13045c0001047c33000c01045300030400c3003333c4114004c5f700013c3f04000300cc0000001d0100050014c3103404301001004c40d4001400d1000000400003003070000000300c1c740400c30000304100000031401400043001c03f0400000004001c0c0c040400400c50013100cdc1c00cc300143c040c000c0070c004c00000031d300c000400000001000cc35444c034000c04000030000c1c0000030c0030530c0000c3310c0300c050434134300000c0f00c0c14400000c014304040070000000000c00c00340010041300000004000310c40c00003c0c0c003010400000000140043000c004000c40113c040c000cc310c0000c010c003400c0010c000f003c003c0cc40101c07d100d0cc40500000004400000004040004000110000030c040714cf30d41000000040300000c0c44c0000f01004c00c1030144000100cc303f04370f040000005d4c000f0110000000ccc10100000013c10100040540000cc00f7044c0c0000000044040c00000000034300000000034003441400f030c11c0cf034130003000000c0f0000704501003333404000d04cf00110400000300003c00030130004cc40773000c10430430540c1000030000000010001c00040003040030000433000c4001c4000404001;
rom_uints[789] = 8192'h474000000000c4c0011000043000114040000000c0f00000100c000001c4040c1030157d00110000c050000c00001010030310d100000001c00000004340004000c050104000304110001000d300040000f0c0d11300044d00401c0100000433c0000030000000101000000003c33014c000003300f00141000c041144140000000500030c4000c30001001000300c00000000000000033000000000c03003100c000300c010030003c400000000c00400c00010003010c00014000001003000001c0000000000007001000000c11044001040c0000030c0000000c000c300701411c0000100c100001c0030c110003d04000000000000104010c000100000500000440010401000011000d00343004053c0c0c510c050f3c000000c30033030030003001010c00010040000040000c010030000000000000000000030431000c1000cc4110c000010c00011400040000c14300401003000f0c0c0f00000400c03c4300301000040000011313440cc1c0300c0104c000000c014d0f01000104050000000c0000000400000011143300c000004d0000001401010c010f10001000c1000c400c000030040100000150000034000c100f0004340000c010700000c30100440ff100000013000003700c0c03c000000400041000003005030003350c01cc04000000030d0c03003c4000c00000400c00000304000c000c0c00000300300f04000000000004040f100c000000001300000c1000000107000dc0001000300010040f53011000014001cc0113d4014300040400000005cc000fc0000300c000005013000030070535000404000000cc0010c1000000303c0000000c0c030c01030400130000000015000001031100010043050401100504000c000330001700f40000010304040c01300401014003000110cd0000001000000fd00c40100fc00030c00000440000340030100000400000000100400c003030044000100010474c000000000000700100000104000040300f04000c0f3100f14000130010c0000c030004003c00044000030010000005115001000000010000c3f0c000030004300000f00f31000c01000100040000000001000000000305100c010010450040000300400c00040c000c50011000101003c5000400000000001c0c000c0100400c00003000000c400d04c0001c0007c0330f310310400c01030c1030310005c3070400000c0010000007000c70040101541030000004040005040037c30003041003c004000c0c3040100004041101000c4034f040011401400044000001c0d000c00000cf3000040005000c000003c1400030000000000c0000010c0430040103300000000043010500000000040c000c0c0c3000410c3054000000000c0000000701c000000005000000000000c0103c001004040d041100000000000;
rom_uints[790] = 8192'h10c000001000004000c00000004c30000010100000c310000040000000c0400000f000000000001000000010010c000003000003000003100000000000000000000c0030000000130003000c00030000c5100000010001001040301000004000003000c10000004000cfc00030133000000040000f11d500400000500100f00103c1c0000000000100000001000007010000000000000000003000000000f00000103000c040000000000000c01041000003c00000040000001000c0c10010400000000000000000005000c000cc0040003c1040c001000000001033c000030000000000054000004030030030000000c000100000c000000000000000000030c1c000001040030000001003f00000101000054c400100ccc040000001000040004000000c300400010001c000010000703000100003000000000001c1000000000000c010001000301000001110001003000100003103300000001000000000010000303000c1003000400000003000001c000c4100c003001000c05040000430000c01c00000001000c00010000030000100000001100300000000000010000030003c3c000000011000000010c00000000003010c0000411c0100001000400000433000430010400000000000000000000010030403c000f00043c0c10000c0000070000003c335003000000011000001100000000000000000000000001cc030c0100000c00000400001000000030000300f000010c000003010000000040000c00000000040000000004000007000d00010000014100300000000000030000001400050000033104000700001150003000000004030000000000000c070d000000c300031000000003000c0000310100000030010403010304000000000140010100000400030c0001000001f00000110000000000000100000400000000000c0c0c00c00c0000000c000c0300000c00000700003000040100100400000000404000000c003c00000400330000000300000c0100010100000331000400030000000000003000000004000010005300000c000400000000c0000c001010000001033c07001350003001000f000000000c03030c000004000400010000035000000004301000044100000000010000700c00100100000c0000031400010004003003000001000000040001000000130000340000000403000030000000040d0000030004000400000000000400000c00000000030fc00010000000000010000000000000070000000c00031c0333100000010c3300000100040000c1000000040000000c070d00110010300003000013000c00000730000003000300f400000000c00000033c0003300000340007c0f000000000010cf0110000030001000000100054000010000000000000f0000c030000030030000000000000000000;
rom_uints[791] = 8192'hc043000000000400000100000c0401000000000000000c0000000c0001000400000400133400040c00010013000000000000030043000c00030400040400c00003000101000000000000000d00000c04030010030700000c03330301000d000000000004340000030040c301000c04c000010c040110000100000000000004010005000000000000010500c0001001040400004c000301003005000000004c0303030300030303004000000000000000300d30c000000004043503000c040300000004000000310010030000c0000000010703000000000c0000040401c0004000d0030003030000000100300100000101040c00000300000000000003000000000000000c00000c00c0000c0000000040030001000010000000000000000001030100000400014000000000000c03000000444c000040000000c101110000c003000000c000000c000300000400000c0031000014003f0004000003000100000100100c0003000300030c0000000401030400070c00000300100f0c00000100104004000000000003000000000cc0000000000300030000000c04000000000000100000010400030040000001000000030300cc0c040400030003c7000001000d0140010000040f05140000000000000100040c0003010300030000030c0003000c0000000300000000c0340101000000000c0300000c00c00000000000003c000007000c0400000030011000f14100c00c3000000000000400000003010c00000000000011000400003100040004010304000000000300033000ccc10001300c00000c0c0f0400030f000c00030000000003001000000300cc000000000301040000000001000000000440030005000000000101010301400140003004030f0c0c00100000010100000cc4000c000000c00c000003000c000304300100000c00030040033c0104c00000030700000c0407010c000000010400c0c30000000c10000000000001000100000303000000000000003000000003000c000000040000000000000000000003400000000000000001010000000005000000030d00000400cc00000000340000054000000100d00c0f00000000030030000300004010030100000c03000300030000000401030100000000000000000300c103000403000000000000000000100000050031000400030004cf01050030000c000c0f0000004040030f000c00040000100000010000000100030000000c000001030300030700030000000004000000c00c010000000000030000000100000003000000040cc10c00000c0300000000030000000001000400000000050d000000000000010001030000040001004c030f00000d00030000000004000000010400000000000c4000400300000003110000000d00000000010001070005000c0100000003;
rom_uints[792] = 8192'h400000004000000040000030000033001340133000c030003030305104113000001000004000000043003000004d000000c300001003000000000001003000c00001000000000000000033000014000010c000070000400000c00100c0003300c40030004000000000000000c3000003300000000300003c50f0c0000400000d007000000000500000000000000010000000000000000000000000c1d0000100c0100001001000000433003540003100c0000000030000c00000103000100000000003300000000000003000004300000101100400c000c00c00000c00000000000000c0000010000000400043000041430000000000004c0010c000100041000000001010030040100007003000000000c3000000000300c000030004000000130000c0000300003000013000003000c00040001003001000c000003000003004001100c0300010000300000000000000001000000c03103001c0000000000010000041000000d100000000000000000c003000000000007300300000300030034000700000000000000000000040100000000000c0000440000000300000014001000000430300cc0000000011000000004400c0000c30000c0000000000301010000100300000000000c4000000c041430000000000000000004000010c000000000010300030300000000000000000000000000c000000000000000d4300000c0000000000c0010034000300040000000100003000000000003000400000001001000400400000000000000000034040000000000000410000000000000011c04000c0000000030000030100f30000100000000000c030000330004100000000000100000030000c4040010000000000401040000000000130000000000000d00000000030000030c10c00300000f400000000301000030000000000400c000043005001303000000301000140004130000030000000000000c0c00000000000000000304000000030000000000000000011000c40f004434030004440100030000000c040003010101000000040000000000000000000000013000000000040000033001105000000400000030f3000000000000000000110010000000301000030000c04001000000010000000c0310000031c00004000400004000450000000000030000000000000000010000001000000004000000000c00010034000d00000000000110400010000000000400000000130010f000000000d00000030001003000004400000004d004011c30000c000c4300000300000011300000434007010c004c00000300001000000000000000c003000040000000000c000000000003000000000000f401003000000c044100000000000c0c00140d0004400c010304c03000c001100000300c00000c03000100000100000000000000000;
rom_uints[793] = 8192'h5f4030400000cc00cc007000cc4c0c4300044000c0c044000070c0c04c05c0cc0005300c00c40000000c000c000004074004430000110c503c0000040100003004400000030000704000013000c0d1004000304c0070000040d00c00400401300c000000000030000c030000030cc00c040034400c0700140074000000003100c4c04100500c00c5043000000000f0c40070000c00005000000104740401f0044000440000d04400410400004c00000000fc01400000000d0c0030000c300400410300fc000400c00c400004700f40104004004000000100030300c0c00cc01000cc000000c40000000c00c5fd40003cc1510c00004000404c01d0c040000000440010ccc0c00004007040040140000c000504114f400030c0d000004c040d00c00000000300cc0000c00c0004c040d03dc0000400004000c1004c00040c010c005010c0044c0000c003004c34030443c401c40470d00000c510c700c00004c000c014034040c443c13000cc00400c0c04000c0c4f001004000cc0c4400000304c3c7f40000000000400c00043c0007004000004000433000c004040000043044c7001c1c0000040000000004000000004405411303007c00d00030400000504f34000fc0000103700071d00c1c00000c03000043000000704cc000c01c4c00000000c0c0040c00000f0000c000f00043d00c400c01303300030000c00000004100007430300000dc0c4c3d000cc0c000c00c001000070044300000c00044000150001c010400043000040004001000004401c00000c0440c00cc034404054c3001000300f0c140401cc70300000000340c00000400000000400004000c4400f44d70c0000c000534000400c301000c1100300000000430ccc4130000000c03030154104c50010cc401403000c401030d0c40433007300cc00003000dcc1530cd00400043000700c7003000c5000000c1f0400c7c001000cc000c540040000004c10040400000044440c00000040400300c01c0cc4034004000100f4000c000043004f000001040000c0000304400030c000c00c4c0c0c0000000410403003005330041c5400c4c0c1c000403000c0304000c000000c0004c00c00040400c43014010000100040010004f00c0000304000c1001500300000c010004c300004c000c4c0c0c00040040c00000c4401cdc40c0c00c1c14c00c030cc400000c4074c400c30c1040000c4c7c00c40c00c1400010054003004f04c40c3000010005f004cc004043000cc004040501504000000030c04030000d4003c03c300c10c00004040000f0c00c17c01400000000000f000f4000c4f000001c1c01000c0040c0000000c00000000c04c003c0000c00400c0f00f000004400400001f00c0c03044004cf00c04030074140040c40310000040cc0c000030c4d4c000c03c40000000;
rom_uints[794] = 8192'h300100010c00043c433104400c10705000004000703100403010c40c1037300000303111000100030100300c03317d10130c03005004c10c00300031c01000300043000000341c0000300043000101c300c04c33c70015303500f1014dc00003c31d101401300030c000001001131501100d1400005404000330154043ff000710fc40300c00000000000413c3003d003c003000410c3031003000010c3300010d0300331407c000000004d001004101dc000d00300d30c0c3c043ffc041000004100c00030f0050040041f0004005001174171430c300f3101103000c00003400000100c30000001c00011001041400000f05c00c0100014d40c00c410000013c011003003733000001d045103103013007d033c10003003730ff0101011003043400040007053cc011301000100000110001c110cd0030000c03430114c0cf10005000013c001000700cc3704100d31000003c4000104000370010000004004344dfc37000c303c00c30000c000000040c0033100100ccc17300301001001d303003c0c100100100040005010100000000300000c500000000c0004030100030c0001054713c03300000d015003031001000c0cc3001ff440400103c540104401411cc10001504101f01541300005c303051000310400031000000701d700000041010001001c30000150010010c100003000c30300cc10000033000403104000000003100c000000410d0c0000c00cc1f500303c10005000430cd0f33100310005c44dc0c3cc00cd5030000000001f10c00c100000000310c000300f00f000400041c0003000f31000100cc700701400300304c100010031d00134000cc0547130017010401c0007403000030000c30110000cf0004130330c00f40340c307cc010d03301c4017500c0340c04c30d103d0300300c43030003c5000000004504cc00c3f5d03500c040c140c001304001300f0335cc0000040050010c00003045014000000004050c04050403f031014014001335001301000103f10c0301000003004110007004003000000100111010df0500303300313d05013030c00010000d0500c000001300c005000c107430000301004100000003c034000000030710004004403003143d040c10000c0cc04010310100000454411031c3cc440004401300000500007005cd00f3411000044d10150301031500d303003003030c050d035300c100001303cc0c43000305310050cd40f3c00010000cc401340104f4f407040301c300750c000d030f1704c000030c0f0330010000300c300003c00c0510100100003c003101d035f000000400c4430000100010c30000000fc3100005c10130115103000031000000001f00304403100301341070000c44c030c5c3000000003cc00040440300c00c13000d00000300070010f3f003100fc01100;
rom_uints[795] = 8192'h410050000100000000000000d0040300300000100110000004c030007031c0000103c11004400050c300010c00f0305000000001307001004000010010c00030000040400000034000003303f000300000100c4040d070c1d0c00000c000003000c0d00141003010400f0003000c0000cf000004001041c000f0001003000030c150430000000100004000c00004c03000400010000000003000000c003000005cc040030003c03c410000000030cf00010300000000037300000040401000c11003f0c00003c0040050000010004000003030004000000000304c000140000011334011d313000000004cf0403000c00004f010033000400001010000000000c000700040c00000004040cc3400c000100000d300000000f3d000c03000000005003000f1300030001130c0f3004c0101c3100000303003310000310f00000cf1f10030000140001000004000100000c0001050100c010cc035005000000000c03030303103c00c30c03540000110c000000030d4c4000001401003000330c100105001300040001dc00000400100110000100cc000000300000041c00030004c40003003f000003010c003044c000000000010c0140000c110d3004003c000004000301030001000f04000030003005000000101c1000000c0000c0030000050003000404000700c00c0030000005000000103000000004130000c0300000100ccc0000000000403011100c00000003070004100540001c0c501031000004c00130cf10c000c0003034110d00030f03043000010030040000c0000d000c1000000000c31c01c0300300c000030030010d041000010300100f00000300000c010c00000c530c00c030000004034c1004000003003004010700c40c31000c000003310c0000030c000000003004040c100c04000003000d00340c000c0400004c0304041000000300530c130014000f014c301300000444300103030500000000030104000003000314000c100c010010001000000033c00c000f3000045c33000000001050030400000401003000040f000c00003300000000000433000000100400c301300c1d0000010400130c30c004011007000003010c0f0f110000073004000403000c0000130030000c3400000c301c400300040c4300040000000c4330000000410030103c4333400000011d01330c0c0504000000000000010c0400000030000c000c0f000000110433001310010000f0100000c0000f043110000400301c00000c03000c0331001013100c0400050013030000003000f300000700010c0000011301003100010000003d000001140000004000100400000c0c00431104130c05301304010c1c1410000c04000004011000cf00001000000f00300c0100001003013c00d13c00000100000c0000000c001c0c000004030c00000f;
rom_uints[796] = 8192'hd04000010010073410130d107030044003c40000c1140134000c0c00100707000003033d13000000070000000300cc10403033030000c00f0033000053000c11000000000100100030003040f303c407d043000000c3100030300f5301f31dc1001330c433000003100003000300071000404c3c00330303003c04cd031303000c04f00c000000030300001300011000044c0030000030307003304040431d000003000004030f3000fc3100311c0003000107c0000101547c030103114c010074fc00c001130c330000c11343010040c100c3c310c000c1cc0c01030c0500000c00000000f3c30000300140433000001433d043c03c010030000040031000001c030000000003004000f00300010d01004300c33c31c733c037c0c000140101c0530100030c001c111030c0f3c1010700000000d11c000000000030001000000301c0d001410500030000c100400041030003040333300c0fc0c44403004000400033300f01c5310c4f00001c0170c330404f10000010100011c11003013c01f30c0030131c0c304000100101310030350000400000030131d10000100003030113011033031300003d31c001043400101d000410340340000030000130c3000033000000c0003c0f30c00c07c0101100d0434000c010130010340103c0d04c3000041000010031000f0c0354000010030404001c000100c13000c300011c310f300333303000003030047710000000cc0101c0070041003300135001031300340300c00010031303011d0030333033c0fd1000003d0030000001103c0031cf0d000c10003100c0c73d00c1000d0103100334003000330370010010000030004303c03007000010003303031dc54000000c00c000040113040301000403003000f43100000000101130cc4010010f03007c1c00000100000003334033cc033010010300004000100cc0c0c11000040030100100000000300c0c00c3100c03f0c0000400000001403f000001403300c040100110333100330174701c00c0f00300000c005cc100000000010303100041c00000d7001ffc0303100000f0001d4c7300010f000000c10300000300030300331103c000000d01003f00000000001313c300c730c04fc0047c0000000003040c03d00000734c3c0700030c003103770007330c0000c00c011300c03300111400010050030130100000030000f103013100001000010004f400000137003310c00303f1c00000000c140001104045cc0004347033401005c43c0010300000040110c04100300310130010010300000333000301000010400c01c00cc1001103000000001100130007000000000300010004c10c303103c000cc4d11004000030030c0000000000000000001041000103041000040010c0f00410033001003037dc0c1000f00c0001030300373010040;
rom_uints[797] = 8192'h11004000310533000003000100003310c00000003301000f00000000f10c00310000000000030000000000c0000500000400030000000f0400000000003000410000400000c0000030c01000010f001c000003310c11000000000011000433000000001030000010000003c00340030103030000030000011003010100c000c000000300000144000001c00003000030000103300c00000c00310c00000001040010000000100000004000700500000000000000000c30000001300004000000400000000000c0404f330cc1040100c0000040c04001000130000134000c00450000c00000c00314f0400030000000030000000000000c0000000000000001703400004100070c0000000100004400030000330300300000001300003300000c00040000000000300010033031000000000001001f00000000001000500100003f0005010043000000000000003000f000400c0005000037500100030000010f3100001000000000001000001000000004000037f140100300000f005033c000000000000000003003c100003000030001000401001300000000001000000000000100434000034400030000000000010000000000400000c0000300004000000030053100000301001003c00000000104031001000010000300000013c004f000000010400300000001030000000000000f0000010000000000d00004030033040700700000100000000003044000003000430001000000000300001103000300d00000010c00000000010003000031000300100001000010001000000500030c00055000030300400000000000013300000cc000000400000000f0000051c00000000c030000010301300003001c10c0300100000000000100000005000000000003301001c4000c0003403c000c00000000000103010000430330300300c00000003001400130140c30010f00000300730000011c0000000000030400000000000007000010040000003f0300010000c00000031103000000010000000040000000030f030000000000000000000030000010000c35000003000004030300003001000300000c03000500000700000000004040400103000004000000001000000000000001000000000000350303000000000000014001003030000400030000000500000000000000030040c0f0000330000d004000000000000c400004001031000000f000000000040003000000030301000003f403000300c01000004003100110040c000000340001003000d00010000303110c0003000300000300c3000040000001000000000c010c3f00000000030000000000000003304300030301000000000c0c0000000004000100000100310000000330040000000000100311c031000000000c0050000000000031010000000000301001;
rom_uints[798] = 8192'h50000001400330004001030d0310404c07000c30440000000405c0000400700001c135c010c0010003c030343440c044c0001c300000c00400c0c10300cc04400010103010c340000010740c00c10f330000330f4700001cf15400000d300000cc31d30100001c000015001c000300c03f00c0c0410001000d0010cc4340004101440000cfcd1004000c0c44000001c03001440001c030000530040003040010c51000c30103c010310d000305cc00430c10000000010770cd00c30340304033ccc050300051003c04000040001001c0c0c3dd00044011000c04c10003c10541d04330cd30340300100c350705000cc01543cc050cc0070000113c000400000005c00441051031440cd1dcc107300044c00c3140000500407040110004c0033500010000100034c400010c00007011d030304404330000430c00007d4710c000000111007330400100400440303000004c1030470003c10c30014004004c00400c0c0d1001340100000000004400100c000000004344000c4551440000700cf033c34003c40000001d010c00000103c40000403100cd00c011cf00304400100013401d030300010c000100c0d1000034c03000007000017000dc000030c0c344dd0305010400f100371000000004700c14400000cd71000c730000103004fc000003f0003301300040dd0100004447103000700f000050000f1040d0031000c03003010004443007043030cdd01400400041001040030041c0c0f043001005cccfff0101010103000003034300c044001c4304c1c0034004104141001000740003040030010300044103100cc0110cc000001100000010c0300043c00004030cc0030c0404007000730d405300000504007003f3474400001d473100040d00013030300000000701c1cc0c70000c13753d3000010000300003400001003070c000433400040040c3cc0004c3001000c10040c043040014330300700000400301040000140004c1cc0700c00c010f0c00d041000301040143004003c4003c4010000000000000c70000040311c043000000d01f3000000c0c0403010140030330001000010000cd3c0c000400100031000143c113000340000000003100341c30f00000000010070030040100004003310cc70113cc30300010c1d104004730c34343cd0000300000c0dc10c4c100011000000103c34143c043000103000f040000433300000001c00000040003cd001410c10103003010000000c0007303010300dc1d00030007d000030013001005001005001c0000040f0047004000000000000d003530053c4000043000c301c700010047330001c043440100c145000111050d0077d0d000d0c0c0504403d00301003003000030cdc0000100100c00450c034400304040440030000000070400c0400c0300030000000000c340040004;
rom_uints[799] = 8192'h300c00000c5510100000cc00000044004003300c000010005c500c10047100000000fc400000001040000c1000c0003c04001400330033030000000000c0001c0000000c000c000000300c3400000034340300003040c43c143cd000d4007c00041130000000300010c40c00141014400c00c400500000000000131010301c1c001c0c003000000000000000100004000000fc00001010c004340001303000c3c00300040c004000301000000000100040f000000c0c5400103c404c003000001c004c0c001414401340000f1030cc0000c00000140c30004cc00430c0000000440000014c5004004030c410d030140404301c0000000000000000f0040000c0ccc440d054000010c010030c100030100c0000300c0030000100000c000044c00440000004040000000000104000333070000400300400003400103f0cc400000c101000c0010030c40004300c000c3c04001033004040330000000000cccc1014001c7440003c3030100104000c140001000c003c0000003c000c00000c00030f100030000030c03000000c00c00d000c00c01000cc0000c004000000300400c00000104400100000404010344100c0300c000c30003050000004d40074303c30001001040c30c0040000000000401400c000300001300070000c303070f04000401c0c000070003000003010301000040010000c30c00000040044330c0f7744d0f01c01301000000c00d07117000c0c300401000000c04c04003f1cd30004c0440c0030c014000cd03cf0001004003000003c44c0040cc07c300300041c00000c0000003c30004000040cc00005010c301400000073300c00000c00101c04040400410000100c10041000000404000c300000101300100030103404540c00310000001c004c303110145003f004003c04500000104c0000100015c004000031d000f0403074cc3c0c00700030fd0030347040cc101403001030c000000c0010040c000000040c0c0000304030400014c000400c00c0cc04000407000000000000003040c030004000004003100300ccd0c50000700000300cf13030000000007c003cff0c3131000c040000000100cc0340f0f03c000c141430c13c0000c0c400001400301030010400000004000400340030c40050000c5404001c400c00000000c030003000040004d0004c0c00c03404030300c400400100010c300001000010cc0f007c01c00c0c4cc0443c3030c0c0400c3000d3c0000000007ddc3040f0000c001000340010c0040005013003301000000000c000500c14000c00040c10010040100cc40c0c0030000000000044100f00c044004010000000003000d0cd303c3cc4040000100c7010000000040c40104c00300c0c00103c4130c104000000300c0000003000300044043030c00000000004c0440100d000400400;
rom_uints[800] = 8192'h1001100c101000010440000300003100300c00043c00301000000c000c513300000000f3000440000034000c000c0cc0000f0000100000000300003003000010000003040010001400000f0c3000c700000c0cc1000f043000030c43000c000c01000d0040000c4400d04000403d0101303000c4000000300000003c70510400030011000000001000043000000000400330000000000000cc000c0000040000001c44000000300000000011300000c000cd040000000400001000fd374403000000004000000400c0000000000000100000100c0010000404000304c0c0010040400000000303000001001f0014330000143f00000000003000301c0c000003cd140001141700000031110c0c0300000c30000430300103000c000110000c010c00f30000000c00000003100104370030010c0f00000000030c000c04000000003cd000010fc00044400d10000c070c000010047100000d0000000c700040030400000100d000040400c00300400c0140004000c4300c0c000c001000003400000000300300443000c0300010c000cc000000cc00000000000440070000000000150010000c041300340c0c00435010cf34000003000c14300c3f40011030f410c0000003300c30040d05000001033004043000030100300400010000000c03030c0100c00c40c1103014431031000000000c03043033000c0000000c0c000003003010100310cc00030001000300000cd0000000000c00503003403c15100000000400c01400300000c00c0c000d40000011005030041000100000c1001013000000004103000400c00314000004000000cc140c0cf4000100010d050000c0000c001030700c3000004040000000014c00310710000c100111c30000030000100000000c0000c0000400000300cc3000400001000f1cc0000c010000004001303014471003f3440003000c3c00c033514c0400000010fc00000cc000340000001000000000004004000c0f000400000000713300130000fc00004c001c4040140000000f000000000f33000001000100c0510f00030000140cc00004c40d000c00c000301c003040000000000000000010000000003003700000000000104403cc00001100730c3cc0000300000000000400000000001030000400033c4c3040c4013300000c14030c040c004000070c000000011d044c30010000340cc333000000000000000030300c000c0d00034c1010000034300c0000003100000c040c010000010003007f030050003000031d1100c00000500050000100400040000cc0010000c0c000000300000000103000040c0d0f001000010000003000f03004000c03000300d5040c001000010000000013cc01040004c004110010f0d010003c000000033047100c400000013100c0000030000040307000003100000000;
rom_uints[801] = 8192'hcc000000010c0000004004001000000000400000000cd0000000000000000000000030c000000000000400000440d0000c0000000400003400000000cc00c400000000000c00000c00000000c0000000cc7d040004c00000c000c0c000014cc000040000100000000cc0040004c40400000000040000000000c440000044000000400100000c0000000c0000000000000000000000000444cc0c0004100000000000000000400400000040000000004000fc000000000c00000000100cc00004000000c30000000040040c400c0000000000503000d00c0000000400003000000004000000000000000000050000c30400c00004001000000000000000000000000c0c040c440000000000c3000400000000000000000000d0040034000c000000000000cc0000000000000004040404000040440000000000000000000c00000000010c00c0000000004000000000000440004000040000030101000000400c004c4100000004040c00000c000c040c000000ccc0300c0000f000500000000030000c000c000000000c00000400444104000040000000000030000000000c00014000001000000c000000c00c0c10000000000000003c04000d0330000000000c34c0000c040003004100004c004cc0400c000000000040c0000000040c0c04c0000c040000040000001c044000000000000000c000000c30000000cf000000c000000c0000000c000400400000cc00000000000300000000000004c0c00010000000100010000000000c000000010000000000000400040c00000000000400300000000400c4000000030000011000000000000540000c00000400c4004000d00c0c000000000000004000004c0000440c0c0001030c4003700000000000c0000000000000000000440000cc000c0340040000c330c100000cc000040404000c0000000000c00000004010030c000000000c000c0c000300d050004000000004401000000000c0c010000c00000c1000004c00000000000000c000c04000000000040000000000004000003000401040c4344c04700c0000001c000000000000c01cc404000000c00000000003000005000c000000000c040000400c000000103000000400040000010000040c300000400340000400001001043000000704040040000c0000000014000070000000c0000c00000100000000000004400030c0c0001000c0000040040000c0000400000c400500040000100000000c03000000100000000000000000000014c0040400010c00100400000000000000330000000c00000000070c00000000000004000010000cc0000c1c000000000400030c00c000c0000003000000c0c00000000400000000000c0000cc000c0000000000000c000c340000c0400c04000000300c000000030000c4040000000000c00000;
rom_uints[802] = 8192'h700040004030110000000c301400003310003c0000050000000430c000c4100000000040f310031000000040100000040000000c0310000000000000400000000003000030001000000c0c0c00001100cc10041000c00000c0040c000c100070040040d0000d0010004010303010013030040140000c10000041c030c430000003100000000000000c00000070000010000000c00000001c0000000000000c000004100004100c0000000000400030000c30c00000000c000000000031c04c30400034340000d0000000001000440000000c0c000000c0c031300000703000c1100000001400100000c000000000000100040c00000000000000103000000041c0000030001c40000c40044000f00400001000003010c00000000000041000000030000030000000000010003c30041000000044000c000c10340000d4000000c03c0c1104307c0400000030004010001000100004144430c0005000000000d000000000f0000007c0f00030000140c000040400300000f000701050f03000071c001000f00400000000001000c0403c1000400000007070001c00040c3c000000c300c000c0c0000030c00041005030400030003000007300000010004cc00d00c000c050c000000000000300000034000000000000d40031001000c0040030000001044030c03030d400000c0000cf000c403030100c40500000003010003000000030000040004000000310300c003004000cc00050000000000000000300140010c0003000000000c000000000c00c003c00441000000000001c3004073010000000c40010001000000004040040001000000450000000010000304c1430c000000cc400040000400cf000000d0010403000400000000c031000400c000000105000c03030f000000000300000301004003c100000100041c00c000110000400000004f00030305303300300000c00c0301000c07c0cd000c470400c0c003000101000000100f070000000000030000430003000001400c00c000000000000000004c000d0000c0c10cc1000000000001d100000000c0400404030c00404400040001300001c100c000c00300000004000000400100010c0f000c0f0000040c00010c0c000000050041000001000000000500c710c70c00cc00c00010000c00c30000c000003010401c010003000000041000070010030c0c00030501001300004f000300c0000003000000c3003c030407000c0003040040000040440144c100400000000301034c00430c1c014c010000001c0000330000000000000000000c004c004004000000000c0000400031010044000300000c010000410000000007030c000c300c0000040000000c1000000000000000c100040100000304030400c301430300000503010040cf004400030340000d000000000041000000;
rom_uints[803] = 8192'hfc10000000050000405044f0f00000043030c4043010d0c00070400000000c0c040000143370c00c4000c0103004d040401c0000104004cc30000010003004300010f430040000300000031c00100010000001f033300000301070100000341c00cc100c000000ccf0040010300100001000001040400010074031f04c40000c00435c0000c00000043c04000010131000400000000cc044c000100040700400f0d3000c00f3303000001000f40005c4301030300000354c30c0c001003010c1300030c0c000040c0030444c000000c4043000303c0000340000c0000000000010400c000000000000c0041040c31c74c10c10c0037010000040001030300300dc00303030000400c0704c0400000000441c1c00000104040c003000011000c0f000c00030001c3030c0040cc034000c00013000f0001000301c003441c0000c10f0544010f4000370000c30000000000030103030c0400010000000400c100000004000500033330c100400003003104000000fc030040000000050033470004354c0000f000030d11000c3f0340300103c30041000003c300000cd00c0100034407030c1040000000000fcc0fc410010000003000004000003d0303010c0c31000403000301004007c000c103000c1040410003d4000100000300c0410c40330003c000000305003000004004004f0c040040000d00004c010c00000d0000000c00010c4400010c40000101000c00000000400000cc01c000c4c10f007000cc00000c0344104300000303c303000000c400400103c000000cc301000330110000c0030000000000040003000c00140cc00c01c0c00000c00143030301040c41c00300c4c40013010703070000000004c300404004030f0300030c054003310300c000030c030040410c001300c10040014000c031c0010000000040000c30010100400c0041070c0d4047c300000500050301004001054003445c01c000f0010300040000000dc0c3000d01010101000c0001030000011d0c04c00c000404000003010c0340010c03440304030003030c3c334f03c00000010c0170470d00c001010d40000040000000004001004100c0030040000000030d030500c00340c1030004003100c30fc11300000440c000000054000dc0003045004fc00f00030003c00001000100000c000c000003000c03c0c0c00c070340c3030003010d0f0003040001cc000104040003000304400404000003f001010c03000340c00c030003403000000c0000c00043c0c300400c0f30c30003c0000300d0030004040103cd0c0cc30000010c00000f030000c0014003030000c04000030000000000000004030c0f0000030c01400001c70000c30001040004004d0043010001444000010300400301c04004c1000003d0000001030f400c00c000c305c00fc00c4301;
rom_uints[804] = 8192'h103d00000000404c000343030003300700111000140000000005000010d0000001410071310000503000c00000500c04d00034040003ccf3103010c0000300030000000c0003000000131303001100031703df0c0001010f00034000c0f10400c0c3450400004001140000700d0100000000010c03001500cd03cfc0400000000f10c130c00000050000050400c00005000003000000c01001100107003140001000000000300000000300003033c00000300000c3cc5000000000434503400000053300107100114000c0000000000010001000414000000dc03101cc000343700000cc000000000000cc4101003511114000000310000000004004010000c00001400001400300f30cc000000000003f0003330410104007033310110003001103000040000100d000134041000100040000d10000000310000000c000000003010003c00c00c4030000030400c3c0014c00530000c00010133c030003c30103000050030013300371100041c300000030000c04001000007cc000000300c00330000100000000c001003c0000031c00301000001000300000c1000c3005d03040001030013000000300010117000000030070330011430000330000c5c04000010030050c0400000000000003300403000000307400110000000003000c00030400010000d00410c0010000004100500300300300400c33314c11000000c003000000000100010003003101000003f0301151000000100304033000300400c30c000011c04000000010030000431043510000031100005100300000504100c5c330500c00000430400100000004c104030d0340010100000100300007040001400311000101003300403000000c530f03010010403000000c000401003000c31304000000000010c3403103100000c30000000011430034110000001400030040c00040000000130000300000004000330300035000700010000000004310030300c10001114404c0c0000dcf30003010c0c4000000000003000100030001004000cd0001400030035300cc030001310140403d00000000111000400300c103c000030000f01300100040000003033040014001000030300c07004105010001000040000300000c110010000100000004c0d100114030c0310c00300040010343300c0010004000c00003c000000330000010010001c10710000103c0300030300010300000100003031300001004100c0001d010c00c000000d070000010404c0c00000054000c30000000151c010053004403000030000100000c001000c300c50000c0ff30d30010004001c5000103531000003d0001000000101000001053c073c041000000303000030004000000000000004100c317c010c0400030c40000030000010010430030004000f0030040400500c40100001000000000;
rom_uints[805] = 8192'h300000000f0043000c310300000000110c00000501003000000d100401030c00000d01001c100000101001000004070c04c00c01110107c0000010cc0f00000000040c000304003d0000011f0000031300100004c03c030000cc00000101040000c004000c00170005000100031000000010000000000000031c00300f0400000c000c0000300300001003000501003400000000000c000000010005040000c33410000003000030000101000c34033100030c0004010d0000000005700000000f000300000c0000000005330f0c000000003000400000040000300c04000c044c100c000f0000000c00040000f3010c0c0000010300000c000c00140c00000400000f100000050fc00300d035000003cc0c0400010000035300000000cc00000f0f00000400000d000005000000001f00030c103400030000003d0000000c010000000300004003000300004c00330000000d0c0300000304053550000300c00005010000010c0003001c00000000100000000000000000010514000000000104030004003000000300000401001031000004000000000f04000030003000000f031000030000000c0c030003010000030c0000040103013c03c0000001c301030000140d01000c01000000000104000400000c00004003040040000400330c000c001c010c04000444004c00000003010c01040c013405030304000000000003013f000404010003000310103f300401000c000000000c000c0300c5030003030000000000030000003c0c0000000c00000000001400004000030400000f0c00000ff01100000100000c0003070500000f00100000030011030004140501070000000c0c00004c10430c1000030c00003000c004003f00007004000d0c000001003100000000000004000c4100010400000000c00000000000000010000c10c00300000c0300040400010004430400000300000401000500000c0000400000000001000004101000000000040404000c01030c0300040000000000040103030000000000000c000000000000000000000c04000c0000001000c004c00c030000000c0c00000000000400000c000104000003000005000000c00000030003000c3001001003003000300c040c03000000111000070005030000030000000000000007c00000000000040300040000000c300333040f4300000c000c0004000f3000030c0f000c010000000c000c000c044f003d0300c00f0030000400010000000703000000010000030c0400000000000100401011000c30000000000c000000c00103000c007004010c0000000dc003030c000004000000450001000010000104430f04000c03000000000f00330c000100000000000030000000010304040500010000000f0c0330000d000c10000f000000000700140c0000030000000;
rom_uints[806] = 8192'h404000171541000300501000c0004d1d5c530030100707004014c00070103c0014c14c4430500c4134004c4f10133040c300017000004340c1040043000013000030410000000441400c1041c014f0500c10503c500404040443040300f4000130f0c100d0c0003070404000c00c1134041000041411c0c00000030c0c40300dd030040044000404005000010004c3c0000000100000001300c310030f00f040030cc0000030c0000100c001031050d0d0f03000005540014100500045031014710431f0400000d300100010404050005000100030001400044c01c00033c0c0104000004d0d3000400533000000004f1334404401000047004030ff00f0005053c47034c3cd0c030100400f34d000030fd1f10cc0000000c0f00c03470f43cdc4301000003000cc00003001013c150330f013100700400c0040f0511300000040003014050c0405001347f000540400000050c15c40c3c3c000c10d0001c1400fd150003400f00cf001001300c0430c004030000040c071004017c00000140c0c54000770c5040cd0c0c0073030d05050c000400001100004040430c000440c305c30f4033400c10f0003300340000301f0c3110dc01fcc1010011000001cc0000004f000000dc00d00304c31c0400110001310143503033330300cc0130311003cf4f0005033540017d1c0d05c10107040dc4000005c54400000037cc30313303d5000f010c0003d1410100030000040c1ffc431030034c01000514153501310301000000004400004303150004000004c3004407100010f3c30d0000041c03030c0c004000000cfc003001013000000cd030300003c010c00077531004c035c010333c40000404d044000401500334041c000030c4000f40f00c30044cc1400c100001100000003c031313010700c01c050300303400000cc0010dc105400f3444401c005c01003301403c003331154000d0130103331400110cc001c5003000001c00000040440300030000000304034c00cc343c000c4034f071300035c4001000301f30f1030030cc003001000c40cf470000030041004004c0150c01f0003004c10c500f10000030040300140047003c0544013c000f400d00130f040030001034c4f00343050f10000c450740c1d0c100c53300dc310c3410cf1511701d0c100747000001d40c0301001000040c0cc0fc370030000c0000cc0c00050c03c30fc000000d01c004c0d00414400c44040010000430401300c03c4004500003f00c01000f00000004cc33cf7300054310033c0c00001100c000103000310044030f30040c04c000001f0044003c0005571000003f004000400007c51000404007cfdc0305c343300003c100013d030330000000000c000d010c3400410c00040000311c054501d007c0000000000f1c00100f00004d1437000400033cf0;
rom_uints[807] = 8192'hc00000fd400000010000000050c000100000cc0400c00014c00004c301000000c13f0300004c000d00030c000f0ccd03005d0001000000000c000000000011000003c04000700000043c0040040500400000c0030000100033cc00413030000f004001001c00cc005000000f000403c03c4000300c14003000404011c0000c1441c00000300000000003c4030000000c00000034c0c10000000400003040013cf700c0003000000000303010001d0000000100000c100001f004dc0030c0000330c003400c010400c041000034000100000001011000c0400304000144003c110003140013014403000100c11000000030000001000030001404000000000000000c11dc1004d0400033000c0000000c0051cc000040cc400100c0110734c00000003030000c0c1014400c003000003300000330c000000011004c0003030300101100c0c000100000c01c0000004340041030500000000041000000400c0010010410f00430c3300015f00c0c10000003300c10000300c001310000c000f0400d003330000031000040003000141000c0c0400040000cf004c0c0000c10403000000000cc0000030030c0100000300000003c000001c00c0f0000000000400400c3030000304004040040100003054000000c000c70000c00001cc000c000303743004c3404c00004000143d00050000d300000000100030000f00000050000ccc00700c0000300410500c0c0cc000000040400c0040c00105cfc003d0c00000303400d000c000000000000000100c53100303030000004c0007000c000000400000c03000004010c0c10c000040004c0100010003001000030330000030c000000d00400040c3040100c00d00030c000d001c0c001c004000cc40000c0000040003000c0000000000041301003cd00fcc00dc0000000c1000010000000f004c0300f000f03004000040100044ccc30c1000000c40c4c0c003304001001030100000000c04030010000001000001010c0000410000c300430c0fc3000cc40000c00f0004330000001cc00000000c040f070000d0000c10c3c000f0110003400304030cc7c4400000003000010000c000300003000043c030c40000f0010c000000000000010000400010000c0000050c001000100c01305400010d00030404000000400000c000f000c010050403c01c0000000c0000f340000c00040cc003cc04003c0004c444001001400c5000000000000001c4003100000041c010000044434000000100000001100005044cc050000c00000000d0300c000001c00004c30000cf0033c033040400010003000010c00c00000001000030000000004040c04000c000003004003fcc030300004030304000000130c4145c00c00001034000000050c00001100f0040030170000000000030000540c00300000000030;
rom_uints[808] = 8192'h3040300033300405300500300000433100030003334300300303101040051100305000441c1000010000003000030100c050001131100330011001d0c3011030000000000000000000001000d000401000004330c0010333101c00f005d00030011000033030c033300010003001040010c00001001010100330004001310000104000300c030000d0000300c000440013000030003010000000000100103c1030030000000103100110000d03300000104000000000010000000104301030011c010030000300014000000000000030010000100300030000001110c0000000014003304000403000100010003100300303000031c0030000000000c00001c0030000000503c00301c10c01001000000c304140f0004000000000c03340403c0000000000000030003000040000d0430000037c4330100100004111c030000c5c001030c000c000000473000000030000134010100000010004001110410000310100c0103010010310f0005004100010000003300003000033033c100300300030000c10000003c000003030310030c001000000001030030000035003130030000010700003d003000000005100330000434030101000c003000300f01010301000100300301040c0400001000000c0100000000c40301000000000c03011033070303415130001310000c1033c0000000010f00300f003000003c0530f3c0000000c011f00300100040010c030000300300400133000410f103000c3300100031000710000000000d0001000010301c10010000010000040300000000000300030004001000f043000300000301003301340107013000030400000314000c3001030000040330100100300011703000000c0103000004301003000130030000131101000017030d011c01001f01d0013f0000300300000d000010001c000000300d30001050100303000130000300010c0000330100030300001c0000000400000000000000000000340110003000130540100330013034300000300000300011003411c031000000003030003005300000000c30000d33c030000000003030030333000010100c10030f731311400031000c34030000000000010c00003001000c7310000400000100000000041050104030000001303310000013501030400130000000300310f000010013000333c014140703430007400301c001010cc3d003030300705011000000000d030300410000110000000000100300300000000130000003003100010300000000130000003300000000000000013010000113000030013400000000000300000000130300c30033011053000001031400000000c410c4000100130000300303100000000000000000030c0300030130330300000005030031110411010000040000110001000003030000c10003000000;
rom_uints[809] = 8192'h403000310703d000010710000344000010100000000030000111007340c03105c141c000403103000000c10000170143000430010005fc00c00100f005000013c0530c000000100000030010000070d310c0c71713000400f403400070c41040700345000000703031430d4c00004c0700cc0000c1001010f4400004431001d100013003300d000000040010000430c0003000010f000f000441c040cf403000014000710010100033001000300300131041000c0d0301030003030000001004d003101001000001040100c0114c7003000c3033004c0303c00000030c4010440000f100040000000000c00c100144c0c31030005000000330000000010740300004000010000000000141cc00c1070c0000401000003000d00040c03013000300d00010000c0c000033005000d4700c103c10c3000c00031c0c50c00043000710444000d3d0070000305000000000c70003141141701f000735313000010100303c0040301013000003305005c300c000001000110000c50104010007000403d13000fc030c01d001013430000713430000110000c000040000000000004004031000000400c000151300014000300c01c30474d000c0100001000000c0003404c31001c001100401700c030000d3400000000c0000010040000173000f004301d3313cd41010000d31c041dc00000010d1137c01004000003001000d0c10370000d0140000331001100130300c10110c1310301d4031000c010c003041040300010003113400000004c010040000cc440001333010100301000010000003103c000010000d40000c10000d34000031043100000040405c10c04411000f013103100c000d04003301030000100104d1001000035c10000034100004114c30000004100d0000310c004700000f03000005001000000c000d4400000000001c00d44004100f07cc0033005c000544f03000007000040c043001101000000c0000003000000001007c000d3000003000030110030000d00010000f5cd0c40004c000000d341000100010040000f31c00410100404003d00000010131c01111050000000100040c000001000040004000313010004000c01000000100310404000c700004c10130511104010000073030001304301001000004040100001004130004010000430400040300400c00410c3100710004300f00c01001001c0000101000c0740030011300030cc3c041000050401000cc00300050d0031301010c00110470010000034000300c001c0400017d704100740000030c0030c73100c00c01041c3dfcc0033cc00003004341010001014000c0010300001100001140c10c00044004110f43004d33c001441100000c0304000fc000703000400c0400050000003004000001c005c010000cc1100c400003c010070707031001000000000;
rom_uints[810] = 8192'hf0000033c5704c703003f300040000000c0c45c054c000000cd1000470f0000c0133c1013030c00d0030040000dd30000f1c44fc305704010040000000c000c4d00d43cc470c013000033010043403147030010cd3500003300000300070001d430044c000c0000001c000000c4040001c00000c0d0c5c0000404c0c41c04f10c4d0000000000c4030300000100c300040000004c0000443003330314001f3f104c0040c00303030c000000c40113c035000c0035c005cc030f1005c0400000c030f001003000000c010c4000004003000c404035c0000ccc0044050400040007000400d0004c0000045043f54000c3c301030300000c004c4000c000000cd00000c0000440033143000013d000000051000000000f34013000c013014f043000010001c1010304000040000cdd000c0cc00c1014c000134f01cc00301d307d000000ccd53400fcc0000c0f030701ccd43c03133400f4140000340000c10c01300000010004010034c34000000f001000c000000c00700004300000c0cc305f0cd00c41c3cc010f030030ff0c003c00000f1000000f3cccd000c0110c000000130004040014010000cc400c140017cc0cc100c30003000c00c1c0c13011103040030010d000001c0c410040003004770c0300c00003410003300cc00d000c04441104f0f0000000cc400330c0000c40030c0d1040004c0c010000130c0d0c04040000cc03300400030004000400030040300f00010000c30005000c000330400054000cc000c3040104073c040000000c011100040c3d004c0c000400c7013d44003cc03110030470cc000c000400c00040000c300004000c000110400dc0070c00301c4d0c41000003c00d0004004c0c0c0000143c0344430000000c0400cc0c300c100100070310010405cc741c100031c000c130f5010cc040100c07c00d3c0c1000000010404cc3000c0c4c00c10c1001000000c000004001000c0000c00034130c0010c00100000c000000010004000000c0003c0d0c041c0010d4dc0300c0401c00010c040c03c0031400000000cc4300c3cd0000000000030f000c00040c0c00cd0010030f03000000c400000c3c01030030000005cc0c0000c01330040443040400f00c4c10c000051303cd04101c0c400000001c000c0004400c1004300c0c000d070dc31000004cc3c000007014403000040105000000400ccc00c040314cc000033c070c0c540014c000430f00c01c0140300300cc4404300c000043000c00c000100414cc410110041100041130c0400c0c0405001703cc001f00310000033144040303000000000f005c0701d500010000003000034f41040c1004000100001434c4c0040d00000c700cc50000000004000c44001c00c30c040400004ccc01cc04c30000c0000100030000c0040040001000000400300040;
rom_uints[811] = 8192'h304400003000030f030000cc0300000010cc30000007030000c0440030334100000010000000000003001000cd00001030010000c01000cc301100103000c00000c00403000000303000030cc0401001031050f3000000010111331c00cc404000440000000400d030c0510000c0510300000110c400000101040003000110005dd30300734000c0010000001000001000000000000000003010c0c01d000004c0000000000011000000c000c33c000f0003c00000010030f100000003500001013400c3001044c0000000030030c0c003001000c0c0404000000000000300000300000010010000c101000c3300000043004000003300000100010000000001000000130051030003100411c300000000cc0051310440c003110000000000c000400000070000c000500004cc430140000f003040030340100000005100300300303040cc30330050000f0300010100004c00c10350c03000c003510000110401ccc0004003105100000131430010c30000c00010c100004140d0000000070030000000401cc1000033000013000104000001000000410004000c00300000000003031030fc000000000003001003000041310f1051404500000510000341010000410003c0000101c00000c0000000314000000100400004000000010300c000c3c0130010c03300501040000000017000100000c0003000c0010000000030ff01d0000010c0d3004100d3004430100000c0004000000000000130d00040030100f0030045000000003300c0c00c000013003000c010000330000000000000000000010000100040300040c101000000003040c3c01000d03300004400c000030000c0414440f0000000c00c040100000130c00303310000074040034000c000d10301010101400300c3c03c0003400010f0011000401000c040001100c00003000000040000400000304303c034300143300000c0310010000000000100c0000f10000000000100000000004440000003000000000c000034000c00000000470040c0fc0040040000000103400300c00c00d300010000cc0000000440000001f0fc0000003057130010c3000300c0d040c3000c40000010014000000c0440000100000c0001c300004000c0f000c00000430c00c310000000017001c110c010cfc0040000c030000014c001000040c0c300110333004c4010000001c00000300300c030310000131100c050000044030000c001011003c0010000330101c4f0000030000040333301000000c00710000003c003c4c00001000c01c000010000000374000000030030404000101040004011c070004003003000000000000000101000c040370003000000c0c0c001000000330030004000000007000000000011000001000051010000d001004103334000c00c4040004003c00001000000;
rom_uints[812] = 8192'h30000400401000c3000003000400000010100001000d7000003c0001300cc0000040d10000100000000c000c0d014300000000010010c13001c000000000010000c073000000010000003dc0c00000003f07044c00c00000c3300c0000c00344c300004dc04c4c010c0000000400c40c4300c530000001c000470030c1d30000c000300033000000000000001001030000000000004033000000010c100000473001400000c0f000400001000c43134005001000000040c0c0c00037c0c000c40400170000010cc00000004000c000400100ccc1c103c0c04300c0dd3400010000c00c0010400000c0070c7c054c31004130000d070000040000500304000003400000c00cc44040c014330104000403330743000031000013c0d040c00000f001cf400000cd01014000004010001100c50000010000000c00050004100001c044010c1005004000cc00d43040c00000040000c00c0000cc001000dc1007030000400c110030503f30301c0c0404d0ccc000010000001430c1401c0c0000040103f0000140c010004c7c0c04c00101100000100c00000054c00000f0040000c50f530030f0000c0400400030c00c000c0540000f0011d03740c37000400c400cccc00c0000000c400110c00c430000410340300400c000403300cc001c403f0300000000c413c300c3d001c10cd100000300400c30000c504400000070034c4d00cc00001c000000014000c00500c0001140040cc0c401400c10d000c000040c30c0004004000000000004f4001010040107700c000c47300074034030040c14000000001c0000001070000000703cc10004000703100003005000c0404334f170100000000cd10003c000c0000c00c00300c030007001d30c13000c001300400050d010400000f041003001c00cc00c44c170c0014100c00c50c10000c004004030004011000010017300d10000430cd00f0c000c000130000f504c000c004400000000000401c0000004000c004045030004300000010040000c30000400003004c00c440044404401030c007404400000c001c0100000000430030000300130004004404000001000133040000740000010000001d0404cf04c034404000071c0001f3010400000000000000c00000f0353410040c00300030401100013100000c0404c00040000410001300c000314c1400c04c0000003c0c0040040400000103c001000c05000000403d0000000100010041030c003c010000173040f00f00030000000fc400033004001300c3000c0000d0700c000d10f44000c00c10d00d00000000113400030000004c00100004400c54000000000c000000403d40000040007140cc0000104c40040c000000070040003000c40c040c30040004143000100000040c000c4c0c0011000d34040030000001c0070c10c00c101000c0;
rom_uints[813] = 8192'h100000000001400010000040c00000440000000c0001000000013001c040c0000044000040c000004000003000c0100000000400c30000c00000000400030c0c0000004000000104000000470000f00c401c0403707000c0c0000040c300000001c4c014000000100d001000c0d000000300c0000c040400000000c0030c00000300040000c30c000000000000c001000004000000000000400034000c500c3c0000000004cc40100000c0004000030000000100000400404403000010700000c5034300000074400cc0c40c0043c3c000c00000005c000c00d400010c44040300c00000c04000000144000d411000300430030300c00400c000000c0000003f0040400003000c000000c0f0400340c0004000000000c0440404003c510000040000c000007000000004000000c40000c04000000000c00c40c100010040f00000cd00400000000000c001c0040000000400c00034000c00500000c40400000cc000400310c0003040000003c003c0000c000000c000000000c3000400000003000403700000030000000003c00303000000000000000004ccc004000f0c00c040404000000041400000000cc00001000c0000004000000c44040440054430d4400000100330c4340303c00310400000f30040000010c000000000440c0040c00005440000300c040040150c00100c00c0010000c400c04040400001400340c000400001300030cc40000300c0000100c0004004400c00003000f0c00000000000014040c3000000000040034700000000c0000400013d0000cc0000c000c40000100400400010000000300000000001c40000c0c00c04000c0040401000000c44400000000000d0004000c00000000000c40c014000c000410c4000000000000001104005000cd00104c05000000004104003000471c0d003010000700000000000443040000000c0004c00cc00000400040300000000004000045c0000c000c4000070c0000400000000c3000000000303cc0c03c300cc400300c0cd10300040040004000000c040c400d00f0000c000c0c440043000c30100040c303cc000000c000004004034400c40000000000c0000c0000000c0004010004f00014c0004300000000041c00c03040c000000000010c4300cf40c0440340103004043000040404300001000005000400300030000c007001cc000000000300000000000000c005004000040000040000000000000c010c00c000000040003c0c400c0c00040c000000c00000000000f0000c440c00400c00c000000000000004000000cc0c40000000030130010c470000404000000034400000c0000c00003000040400013000040000000110cc0c0c30004000040004003000004407400400000000000c4000404c00444400c0700000043000040040014004040400000004000000;
rom_uints[814] = 8192'hc001040000c000000000003c0000000011014000fc000300000c500001010000000000c00044000001c100100d0104c40c03000000400c00000000000d0000000000010000000cc3300003f001004fc403c03001c00f03000300c100000c0f430403c1c3000010c43003000010014cc0011000400040010d0000004000000030701010000000004400c0000340000000000000000000310dc0010c000c004030070100000330014000040d03300100400003f0000000430003c0f001000300000c00000000000111040000000c11500000030004000000031010001000cc000000110000400070000000403dc0300f430c0004c00700000000000407c01000000001c0470000000300000013000000000001710003000000000c010030013000000340000000003030030000030030000400c0000c010000f0037304040c00000000010004470000f3000030030000000000044100540f4041000300000100301044010000000300404000007000000000c004003fc30100000301400c000043c0c30110003030c0c10100c0030000000000000000000f000100c003000000000000073040000100000040f00300003000000c30f0001400003141000000010030c401030010d010004100000400f0000000000000000cc40003000000000400000c000000000040040400010010000013003d3004300003c3d00400030000c00003c01c4f104300000030010c000400000040100003c1030000000003c0003004cc0100110c00c00000300000000044030000000304c000003014310000000000000030040c000003410c00030c400003c1014000000300140054c10001011001100010cc500000300041010400c0500000c30000cf030003c1010010010000000003000000000003000f004f000c0001c0030010c3000000001000410014000140c0300300c053000341c3011403c00000000003000000c400010cfc00c0303001300010000003030000000000000000007001000000c04c004001003000010300000070000000000001000500000330033f300041004100c000000100310003010000300000100c00000000400030000000000000c400010000010c00001001000000477000c004004000c0004401000d0c0000100003000c0000003c0000010000000003300000c0000001000000030000010107401d4043030000330030c1000001c030000c000000000f034000040301000000c3330303004000000030000400500000000000000100004010000000000000000000300300000f00004000013003310040cc10300c000003000f01013030c0000000001c000033c300000000035000000110000000000004000000034c010040000330c0c04c0400000000000000000c004000400000030010100c30000004000400101c041004030000;
rom_uints[815] = 8192'h4530000001004100c000c10300040100c0c000c3010000c001c31000003301c00cc01cf040400000010101000101c0c000f00100c0f1c300400103014000000000c74f70030141c000010dc0c003c10040c3430013c0003000c04f0307c00d00030103030100c3104d03c0030000044000c3cc000cc3c31000c10cc000400043c001c0c0000000400303000140c00303000000000000c7c13030c00c400100c0010000040300c000030100400003d3c0014017400100f131c3400103400000c3cc004330000443c0010103f000330c0300c3c0004110030100c003c13740004007000003c000c00101000dc10c0c03403004d04003c00000000001000000000300030101410001c143440c014010c00030c0000003c00040c0c00000c0410001c400c000030001004040d000c003c0430000100c3130c300030040c3f140430103410071407303c30000c000000000003300000303c10330c1c153030000c3000003c003000303c30d0c0003c1c0003000030001c3c04143004101000333000301c340c1014300000303000000c00110000310c14000000300c403000143c7010f41000d0000401300c0c010001100000000040d00300001410003010000c30dc000000003c0030000f3000140010100014103c00cc303c001314003c1c440d000014040001300f00304c3114dc00103c0c00000000301c000030000010140c0004100c0c00101c14c0000010040010103000301c30140000003c400000300040f45c0310000001001004003000103d00005400000c0c3c04130000030000d00c000000003c0c00000c0130003c30050000040000003000311c000000303f14030410303c300f0400000011340004c0010c300c0010001500000010300c010c000c0c3c010c40103000040014000300dc34c00c00005c1c305c0f100d001000310000f03010f300000c3ccc700c14003c030000000c010c10103c30000000103000003010003400000000040000003c000000104c003c0c14343c340d00f0003c0000000c00000c000c0400001000300000303404010c0c0010d4300c0c14003c10000030003c000c400010003030100c10400000001300000c040000003000000000100ccc0014304c103000033000000c340c3c000c0034310c33013cd00001001000000000001cc131144c3c0000003c0400004700000c00743c00303c0000101c443c3300004c0010000c303c0030300c00d00003100000340f00d0043c00100c3c3c00040c70000040004300000004111004100010301c1430030c0000300f30040000c01300000c1000000400003c1114340004000000100030300003300000c00cc3340d303c00040c111000030c0000100c00c01000000013010c0440100c004c00100c00330000c0000f003300000000cc010034001030000c3010;
rom_uints[816] = 8192'h30700001004c004017030103030003041c0001004c000000000001030141c70000053cc0410000c0000400c0000000000000000044000d00000300000300000000000041c001003000000d0d000040000103300404030334074300030000100000140000000000310c01110300141000c0103010000c011317170c410113300003010c300004300d000100c413101030c0030400003400000100f0c0000400c3000030000c305441040000000001400000000c3000030000110300c10c0001000004400000000000001044010010c0cf44030300014d03f00c07c00001011400001c00000003000000440100000100000000340031c300000000003030000000000030010500c00003000100c0003100c00341030103070005000030000001010001c10005000001c00340100000c0000400000c03014100030f0050c0c400030003c0d1000310003033000130000000030000030000101100003700c001470700000110000500040730000c0104c05000c00000030000310300400000000000000001000500000000000001010010c0000300c30000030003040cc000000104110000011c0000040300010c03311070000000030c070330000cc700c010440c0001004400000041040f500013000c00000000000703c10300010c03003000c000cf0040c30c31034000440000000400030040cc0000004000000700450301100100030dd30000c043c3000c00cc010010010d0010000cc041000000004141010000c0000417003c410001000f00004c3000030000000001c300c000040000000300003030000300303100040010014c0c030000000000330c1300401400030300100010040310000303000c00c300013103300001000340010100010003400001330f000400c0030100000010050c00c30f000101340004004110004305400033030d001010d3050007033df000010030030504d00000003000000c00000000000030c000000044000000330001000000430000103c0000c000010040710c00f00004000100000404000001000400010001000d0000000300c0030000d30c000001000010c004c1000310010000100330010000000000000300400c00004101401c30c0000000030031000000c100010013cf07000100010001100000c30000000c0cc1000300000000c030300010004c0d000300701000c00c05000004c4000d0000000700000003cf00c3030000047d00010103104c01040000c300000033044d30400000040030100000f00001c0030000000110000003030000c3400000045040c1c104c000003000000400001000107000040000011015010000001000004340310035000d0110010001100010000dcc000400000cc0000101011000004c10000001000004000033001400101030030100000043330000000c00004000;
rom_uints[817] = 8192'h300310001000010430000c0c110000003c03010033000d34000000000330411c0003c43011100003000c30300300301000000c00030300f0000000004100000010013110030000000c003100030030c40000130f000010000c000c0000300731030140c000000330000301300400370400031001040310010031033100300010d3000000003301110000000400300004070c00000000000000073c0004401c0010f0003001030c01030c00001c0c000d0400050300000f000100000d0303000003000010030040303010000300000110044000011000070000033100000301304001003000000000303000040003003df001000000000000300000000000000c0003000010300100001c10300005000c041c0300031007c0007500400404330100713000010030003300000000001003010000030000030004030f000d1301010300000004000c00400030000300000c0003c000044031400101000c1004000c30100000010f04000030030d300003300010000033000003001010000100030003031030340d0301000000101000100d00000403000004130000014c03010f0004170005300101000c0c03c10044000d030c10040007040310010010000004003101010403000000300005000000004131000003cf03030301000001050c00010100003000c3040014401d0c040004000500030000100c00030000030000000f040030c004000030300c0300c0310000301303400003000c0000300cd300c700003030000300000700041d030000000100c10100001d000010f003000000000340011c0303000000344d000300cc0001101001411010000010031000030f1c30c0100031300130030c0000001c000170040c000c0004000004010f404530001000410003000000300301c3100113300100171000330300000000f003031005034100040003300300010c170704c0040c13f010000003010103000f000000030c30000510050000c100000000000c00000011300c1101000000000000013700000300000100300c0000400c0531000000030407040000000000000c0c00000000300001311f0003001000003f003f001007000f3010000014103100110f1030071c3d00030100001005003000000c03000c01041500000000040000d31d040010010000001001000300310140000000000010103000c70001543130000c0c1013010c034013130030000030033100010000000c03000030000103000000003110000001000000040000000001010131301300005c140001300000030303301000000001043c10070f0c000000000000c7000f00001c00030100000400000300000100000d0303c03400010000103000000000040000440030000f0033040030c00100000033100c001407c0000000300310000041000010004031073400000004;
rom_uints[818] = 8192'h13000003100001303000010011430073000130000000000304000000000013000030d00570000000010000000001301130000c04030000000010303000000000003033000000050000030c00010c0100040110331000300100000001cc000001700c0000000470030c3000310cd0003000000004000000003050010000000fc00300000100000000000000000011050100000000030c000c000000f03f1500010000c0311043003007000003300130030f10000000100000c00c00100130001300000000040000030301000003003030000000000c1403010003000c003000000000110000000000000df04030030100000030300001307100004000000000f000003d0130310000001000000003000000311340000400040004000c00003000030000000000300000000300000004400c0000c0000000100300010000000000000100031103000003050000011300d103030001007041300101d00000040000300000000100003c30000100000000000300130300000100100c0c00003004c00001013300000000000003000103053000000000000000000330001000000103314c0c1300300100000000050c000000000c00000001001000000000000c00010030001030013003c000100000300031100100100010000030001c010031300000003003000030001001030000000000011001001000000010300100000700300000000000030000300000000000000000000103103001c00400030c1c0000300530001500000000000c070f000003000040010041040000001400000030000000401000000c0030000003c100000001c030000c000003033010010100c00030030000310000001010030000000000300000040100400033000100300000300000c0c100003000353031000000013c00000000000000000001000000000304000300030004000031033300c300010000300000000000000000010004100001000000000000c1003f100000000000400c0001010f00000000000c3000003000000000000301000000c000000030000000030130003300000000000000030000000300040300010100040100000c00c0000000303003000000030c3000000100c000000003000304010000000000c000004c0c00030030000100000003100005300300000000040001000004100f1103030030310c00003c0340000430303000000000000300000133000000000030c300010300000f00005000000000000010300000400000103430000330000031100301c0034000000730300000000300000c1000d000030001000004010000300001f013110000000f0c0000000000010003000000000040003d00000000000c3000400000000400300113310c3030030040300003000f0000cc3300030000000000030000000d0001000040004030000;
rom_uints[819] = 8192'h103100000000100430010000100031000d0130030c00303000053c003c10340000000143000100311004005f00000000300003100001000c000000f030040030000003310c140000000000301000300000010430300013101000031000000010cc00030f3c000000000c300c0c300300000000030111fc140001003300000000000d0100001c0001000c00101400011000010000000c003130001000f004300c300c3000000c1404001c0000c01400000003003000001030000300101c000000000101030c003c1000340035000031003c00300030100403000f301100000c00000c00040c001400000c00040004331c00001c1c300d00300030043000300000000100300c000400031030000000300030c00c50103c31000007001031003c37000c3000000010330030000130033010040400300000001000000c30010010000c0000010030030c0104003c1004001030400000003c07041305000c100000000c0010001040000007d050003000311c00340c0313c00000000000000000cc003df001000f00003074003000000000000000001010000030000000cc0000100c400100003310140010400010043000100000000107101c00000c1005001004300400000c000400000011330010000014c50004001110004c0010300000c000001013301300301031c0ccc000103000003c0010000700000c00c4000c00000031010004000000000c0030001000030300c00c0430730000400040103000000000300000000c0c31100000c30000100130000c00003c300300013c0014000c10d000300704000004000033033c010030000000043030000c00000c00040010000c0400003000003000c00000000000003000000300003f30010c05000404000300003400303003300000100fd300303c00c11334000c034c00001000000170140c0003000010001030303c010d0000003004000000c0000030100000000c01000000000c0005000c000c3000003410100000003c000000001003001000030d1031c4000c013c0c00040004303030000d0000300c0300000000000400400030030cc00c00c001040000110000000043000011001c0030400000000f00050c00010050cc000004030004003c1000000030000c040c054000300004300401110010000004000000000001001400073c10330000001304003f343000040100040c4031101003300000000400140030000000000000000000040c030c10003c300001003404030400007003111000000400003300001500030000000c1c100cd03000300d00040030c0001303000c0000303430004110303000000001330000000d003000001c000000733c003000000030003000300000001030100300300c00000c0004030c00000000440400001000f030100c3003d000101700c070c03000000c00;
rom_uints[820] = 8192'hcc0000000c03000300000000030040c00000004100040000434000c000c0000000000c000c00000000000c00000df000000000440cc0c400000000000000000000003000000c0000000c0c4000d0c04010c0c0c30000c000000f000000000000c00000050000010040d040440004c000000010000c050000c000c0000c000000310c400003000000f000004000f4000440c04000c00010000000000000030100c0010000c4c0300c0000c00000000c0000100000000003400000c0304000000410400000000c000000400000003011003000c0000000000c4000001f0000050cc00010c000000c003300d4300c0000ccc04000c00000000000000c0000000cc04c00300c00c0cc00d0c0010c404000030000000000c0104040000003c000030030c00040000000c000110c40003004034000000040c00000c00000000000000c0400000040000000030000c0000000300400000004444010400c0000004000000c0040004040c000d000003000c0c00c000000d3c004414000cc40c0003001c10300000300000000d04000c100040300000d0c00000000000c040004000000433033000000004004000cc10030100000c00000001000c040040000040004f030c4034000000041c0040000100000000000c0000000c7000000c400004000c100000404000031030003c104040000cc30000cc00c000000c000040c00000000ccc007430c0010000305c50001c000cc00404000c0000000010000c0000000000003c000000040c00000000000000000010540400030100c0ccc400000000c43000400cc40000000400000000cc00000c44400c10000010c000c00000400000cc04440400c0c00040040c4030000000c000000000003000040004c004000100c0c04004000000000c0400c00000c047000000c000040000400000000c00000003400f001400000000000000c0000300304004c0c03000040000440000c7c0000c000004000004000044000cc00000340c0050c0c4c050c3040c0000030000400c00004000000104000000c0000d00000c0000004040c40000000000c00000140400000044000400cc000400000004000010c300000004300400000100000400010d0000000c0004300cc000000003c0000cc000000f010005400000c010cc040c44004000c400000400000cc0c0500000000c1c400010000300000000050003cc000005000c000000000330047000100410010000000c000040000c00c47000000000100cc0040c0040000004c0000000c001c140000050000400c000000c0000c0040000000000000d0000000004000000000404000000003400000c000000001003c004000c100004000000c400000cc400040c00300c10300000c000000c44000c000004040c04003000044000000c0000000000400003c0040c000000000;
rom_uints[821] = 8192'h40000300401100010000c4c14c0000510000404003c0000040c0004000400000d1c34000d0c0010000000040010d07000041004000070100c000000000000001041000000000400000c04c0003c000010003400c3003034100430000dc0f00404040000001041000c01400c00301c3000000c000c1c40000004001014c300c000040030000000000000011030041300000004000c0404000010040c040041c0144000003c0001000004000330000000040d0000000004040000000000000000040c000000010c000400100130104c00001c0c0000000c000c100004000030100000300031000400c40034040cf004003c04030000000c04000c4c000000000c0000c004004c4400000000000000040c0300000cdc000c0c0c00f0141c0400001010000400000400003f010c0c300c0000100030040000000000000d300000000000100030000000100c00000010000c001c0000000030c40410001000000000100c100d00c03004040c300034040410141400003000000034000c00000c0004540c00010030003400100000000c110000100030003c003030003000c04c0411000030340c001040040030040d100010000000000000000c04300000033030000000000c00040130043400000c1001000040000440040000000430001000000404000430dcc0140c0c0000100410040f0c00000400000000001000300000043000000c30000004400d30000100001000300c000400c431030050040034411400000400300d040c00000f000000d01c001c0c0000040c00000100000000300c0410040c0000c0000004000c003340300000000000100c0c00c400004100c004300d0034c43004c0000c0000300c130400000c0c000000000c10040cd00000003c101000000000040000000004000000000c0000301404d400100410cc000000dcf4004f000011001030003001100d0400dc000010300c003cc0000c100400003000000d000000000c04000c04300000000000000c003001000c00003fc444004d00c0000300010000c00004100400003000001c34000c00000400000c10300430000c0034004105030000000010040c000000000000040c0400301000303100400c0000000c010c000410000000000000000c1d00300404000d043c10001c0c000c0c4c0000d040003c000c040c000000c040000000000000100c000030400000040430300c001c1003000000000c0000001c000c40000100cc00000400040c040470000000c0001c0000101004003400001c000000000000300400000000000004000c04040000300c0000000000040034001000000100040400000030c0040c0f04000c00007100000430041400c00000001000000030000c04001100000000000000040400000c10000c00000440300c000004000c003004003400040004;
rom_uints[822] = 8192'h30003000000000c30000000010033000000000070010300000001003040110000110401000300004000001170034000001000103000003400000000300000030070340700c300c00000c000110001000c01003400033000100101100001c00030c0303503101034403001010000c030400350000013005100d0033000030000010000301001000000400000cc0d001000400000000300040430001040c00000f4310700000150c3c3c1c0007000000c007000000000004010c000003010000101c000300000000000f3c00000003405331034153430000100c000c10c0f00f0c0c00030000000000031301000f1410000104000000000000000100d00000003030c30c01c0103300000000000000000003000000041350070500000400000100c4130000033000000000001300030c0004000003000000010003000000040033000c0c010033000410034000c000140403303003341000100011000c0f00100c00c10001000f0101000004103100130004030000050000311c3c0000000c000314131000000c05000310030340001100400100001001000410000413030000003f01400310000000040004000c000300100010110d1001000310c03001004000d3100000000c0300010000070c1000000c000101031cf3000303000c0000003100030300000010100010041003d00f340004d0400300004437130000300f0f0304100010101c1314000f0400003000001000c00000033000040000101000000003104c13010000300030303000000000003d30000011440c00440003000100c40000140001004000000000300000000000010003000000101f045030000040000100000c03001404000000000004100501001444000300033054000000000000c100c100000003000143110003370000110330001000031000f10401c00100040103300c0001100007000100000003000043100103001003400300010003000000000c0000000004000000103c100000000351314c00000404041030130000310003000700000030010000000000000c0c00030000000000100030004004000003000100000000100000033070c0100100c000000000110004000000c0c0010d303000010c01c00500010c030003300000000d0400400cc0110013350411100170400114000700000d000c3f77001000040400c003000000000d000013040000000007030000011100c00031100100000073100c0134130400c000000000000000004103c00c00000110000100010c000071000131c500001c1c0001000003000010001010c0100000001401000c00000c00470c0000d000100c0000100410015114010000c303030010000030d00c04000000030100010011001f000d030031000000000000010101c0401c0c00c0030400000000011100004000100000300;
rom_uints[823] = 8192'h34300000000c05347403000c00000030003f030c00040000003330c0400440300c0cf0143d7c0000000000000c0000f00c040000300300003c1430030c0000000000400c0000000000000c0700001c0030c030531f031cd10004400030d0001001710000040c30000c033c000c000003010000040000001c40000004103303000c4000003001000c00000000f434c040004c00f00000000304000007530100000c3100014410330500000034001400300000cc4c0000004c043000103c400403c0000c3000003d00103c00c03c000010030030d0000c0000c0cc14c004310000003c3000000c00000000113040c000144c0010003400000c00000004004000333c3c0c03cc340c000400004c50041000000c003f0003031003c0300115400404c01000000c0000004c040cc4cc001c000c143c0010010030003000000000c00c030004040400410013000000f000100000010c00330d040400c0041c0c100f4c040010000c30011040000010000c000340405f403f100001c000c00400000f0003f53000400f000003140003c0c4030005003f00000010000c300010044c0ccc003c40040410003100c00410001c00000000000007000c0c3010110000001000c40410345050001c0c440700040000011030001c0c0000c040740440030010000c005001003f0004000000000003004f0000304c440300044000cc0c000040ff001c3cc00003000400040f00100c0c0000300010c4000c10430f100fc3073cc040105dc0000c003c000050040c00000304333c000004c0c000c00c000100c0031010000c10c0000030c403c0000c00040040010030001c00000410000004300d3c0c130013000010100000430000000000001c500034000f00007c000400000000000400100010f0000400c03130030000300c0c07040000000403000000c00000000c040c03300cc0040110001c0c44c000000400c000000100cc0c000030000400740c0000404000030000003000000c0000f000f000000c00d070c00450030100000013d01000000030c0001500000c000350003c0000003010000d00070c5000000030000d3040300300003c00c00003300000c1030c005d050300c00c4c03100000c44c4c300c700000340c403000000cf0100403340000003c000cc03c04030c4d40c4000104004070000c000000c0440000010000100400000c00c00c003470003c0c0000c400003004000000040c4c0010030700140000c00400040f040401c00000f0000100007001d0000400000400303040040c0454104000000010c41400103040310c3010c0c07040030000040003000c340313000000000000040010100cc440041014f5701400000f040400000000001c000003010013033c04001f00040000c0000cf000000703000d0c040040c0c1030444000000004c00;
rom_uints[824] = 8192'h100000030d10000c140304004c11030000040100400000c001f0c0001404400000c0700000007000d000005c0004c03100c040c0007400000c04c0d000c000fcc4c00c000000c00004cf0300040001004001500c303400344010c0043000c44007111010000000100410041003001030c03c04740000003f0c34304000c0c031504400c100000030000000004004344044004000000340500000000cc034c34500000c007000f00403400000c00300c0c014d0000070d00410000dc3300000c440004430030000031000000030500000c03000104f00000430c04005d400400cc0004000000010c01004c110f400c400051040400000003c001000300040c030101034c0300000d040043000f0300000043300c5400000044000c0000c10000400300000cc0cc0c07004c3000c001011300c1000000000c00c100303101000d0c004c040f000003030c01000300101000cc00c74433447000004003c0000c000000000d00100701004cc00f0c000100c0100037c1500c0040310c0000c003170700000c00030000000004030000c100000300004043000303001f700000000c10cd400111007400000c04000d0040030000430043000000004300001400cf03000c0f000100040031010001000003040c00000340f00100030100c0000100030014004100000c17504107c00300003100500000000300011043401004413cc100f3030010404010013000000010c04040001011000d010713c00400404004001400150c4340c30000c0143000010f3000000047000500c10d0033700033000001c0000003040c0001003c400003000010003030050000004c00001d0030f0100c00c44c51c10003003000000040000100d4c0001d1c00110d0000003103404f3014000c40003030000000340105104104030c040c45040000c3000004c000cdc000030001104cc000014300044d010704000300c00103c003001c00000000000074000100405043c0000c0003000300030ff01c371ccc001100c0001103c00c0033001400400c40430107004000043c4740c434000c00330030007c0c000010000000004000c5000000c1c00000f30700f00000040000001000003c00000d040000044f00000100010f401410cc0043000140040101031140000000050c03c1000d000df403000cc30300000300444004017cd10100c1400000000000100c0004c0d10040c00400c400010704fc40100000000c0004001000000c0133000001335c110c00340dc30000000c0d013c4c10000000c004000c0000100c1403404000000004000010000f0c1443003300000000000f00141d010c400000011110000300030f0030d40004000f0d010000c1100400400000400000000c000030c0070001000d47000300f3f000000100000400000300c04d0003010400010000c0;
rom_uints[825] = 8192'hdc0000c0001014300c000c03c0000140014400c10c0030040c04000000f0400004143400100400300c4000037004d000350c0000c40100011440c070314000301000c10300000000000000cc0000300040311f00400001c3004000c000c033cc00c0000d0000004304f155c030007d50f000400d3003004403c0000c30100000404000000cc0000100007047440070c00000c000000f0004c401f000001000000004300000410001c0300000cc000003c0cc0310000004d0400000003000004040030000000044150050c01000003d43c03c1470d0347c000013004400000000300010047d400004001000c1c0330000001014c30000000400100003400000c00000c000000044c034001030004000000010304040cf00c000000040c0010ccc400030000000c000000041c030000044000c00000410d00000cc00010000c400dc30d4c000000400004400c40000000c40030030f074307000000001001004010001300001f03000113c57000410005100cc4140047000c00cc340c40100000030334500d0c000c000c500c000005030000003000000000c0030007004c01400c0341300000403540000cc030c00f40007400cc000100003003003000cc43031000c0000c04c00304034000c454000305c0c0010cc00300400c3c0004cc0c404c000104c100d0cc04040cc7305700013c00000d00c40000400000300c31000051c0034340040d400041001300c10000030c0000000000010303c115c5000001000030000000c10700000fcc00000c04010c0d0c0003304d014d00040cc00f0143c1040700c00100001d000c00011004031441c00100040404000c00010003003c04400cc41000104000400443004004000304000c0c40004c0000000040430c00300000c004043000c00f040001c4000014331000000d001000431005c10c010003cc0f300004000030340d01000141c0400c0300100040413000044000000000c301300100001c0301000400040c0030130c01001000c040010f03000103000d0003c00c044c0000004000000c000cc300040c30003000300103700100000004400d0c040401000300001000000c1c00310400000044c10403044010440400034010310c000101000000000000100040001000000000cc0001001d04051407010f4001000000010000044004000410030c0c041001c003000330c0000003040fc00000c00000000f00040100000000010cc4000001cc0000043000cc03440000000000c30004000033000d00000c10c44f017003c0000001400d5c01030000004000000400004433c00000300000100000c40f01c0000000101030073404c0c0003cc1003007000c00100c00030004100c10000000000000003c10000000447cc0004000100004004c00041007041c001000c3000404c000403000040000000;
rom_uints[826] = 8192'hc301000003314001c00000000300000300400103011000c003c04003300001000110003150400010000000300001000033403030000ccc00004003410000000001010043000003c0000001c000030010001000013cf0c010001040c00030000001704700000000100000000000000300040000000001400000030100000330430005000003000410000041c0000400305000000000100330000000000000011100104000300100000700001c040301100c0100000300010040100103c30400004073000000030003300000400c003111c000000000c03000000100040300000000000003300000000310000fc4003304030f0100d00001030000010000000003001300010031011c1000004143000330040013c0331301000101000000c300000040000030c0c03003d03500000343d000400301d50000000303cf43d1014003030370f003010000c00000000300000000400000010030140001c10040c4000000000303000313c500c004c371004fc000437003c3013c04030010010000004c00c1100d1007c00000100303c00000000000130010000300400c0303c103000101101000034100c0000071000301050000417000010013030000c100110000010141400000030000033030001000000001000300030333100001000334c3010000011033c14303d00004cc30c01300000303030000000000010000000100000030010000c3000010311300100100c001030300000000030ff00000000300c0400000001000d000000101010c00101003000000000040000010000000000303c30000400300c0000003f033000004000c0001400000000000130300f43140030140000103000003000000300300004000400000c00001000001000000030001000401030001000300070100000101004003100000000001000073000131400000040005100c00003001301f00503040300001004040c300c00003011000000003c00301000000000c0000000000300003000300033000430000130030c0400003000c010dc07000010300000000031143300301033030000000011000c030000304000000110003514040430000d00c01000303010000000c0f0f000400040040c1000007c0030001103100400003c0000003054010004000033103004300401401010001000000010401004340d1001c00000000000001c1330300000000400000030000030000000010000000030103030113351303000030000000c0004301000103100001000050c0040000c300430011000001001300c4c14300c000004300000000000c000001000000000040000340000070000110003000034300004000c3c00000c00dc0010000300d0000000000c1000000011100000041100300c00000000f01000003000f00130000000000000c0000000300000001030003000;
rom_uints[827] = 8192'h1310000c1010300007000430c000f100c0301104330c0c30103010005003000000004c3dd0c0003000000c3030303000003000003000000c0010100030000000000015303010001000000104d000401100040004040000031d00c4003040040000103c00000030c000340000001d430c111040001304044000000d043000000031000000143000d4040004000000105040000000000000433c00003000000030f00d3000033100d000004000f100000400000000000404c0000000c0d70000003110000cc00c057c00000000000033003c0440100000000c0000040310001c0030c0000c0004000000000014c010340000101330000000000000000000000400400000c410501103d010000000500000740000003c004400300000000c700c3004110004c0000000000c001c3c0000001000000000100000c0000c04403010040c0c10143f003000003c301004303030c300303040303010100030100001000000047054c00c0005300030100010400000000c0030c0030c0010031c0004000030c1000010c04000003000330c300434000030000000100c0110c400003400001404f01100300c0001000cd03000f400330d30410410105030001000004000100000004c0031000100fc4000c00000003010040413004000000c0000503c30000c00000000101030c70000040000003c47040000100000000000000010300f30100034103000000004330040001000300070004f0000300c000400100000003030000c000400100001041000f0000030041040000c300400000c0001500010003040000c3030cc300c0000003cc0300c4030fc100001000000030000c0000c301000001070c00333000030340000d100100004000000003003100003000c0030104100000000011033431404000030c407c00010433010000000000530051000f0033040c500c00000003410301010000000000004000033000033f00c0000001030440010000000000000c004100000000030100004000030000400001700300000c00070010110101001000110010000004030000300003000000030700030300c00000000000030040000000000047003000130c0f30001c00040400010d0c000000001440c1000000000000000000103304000c0340430400004000530f41430c00000000030000c101040003000c03001000c0000000000000000000000100c3c00000004703000000400001010c0150010c030001000300c00003334040c000000000c000430000070003450100000030c3c100000300c0004f00000000c00000c700d04010300000000000c0014000003000c0003000000040130c000101010113000301000001c0000303d100005000000000000330f501c0000000000000000004004005300570c0000001000c0c0000700f000305c0d0c3000000;
rom_uints[828] = 8192'hc4000c0000044311000340000101c00c4001c00000000300005044000003000310111010400c000003400000010d30fc0700300003000411000000000300370030030404000003000300003f3100000400000000c000c010041011300070c01000004100030000003003310300300c000730000007010033000140f000010d0031000300000c0000000000000000000c00030310000000003301001033001c000030103103000004003000100300030000410001000003cc0f000003c00003000304030111000000041000000030150700001030000001c0303000013000000401000103c0c00000000000001030004310000133000000001300010c000000004000001000300000013303000000001000f00001003d0103c1000001330d00100130140000100340005300040100c03411000110001000003010000003000400000c30330010000001000100010000001c01c00010000411300030004000010001004030010015010000103301c0000030003000010d034030131104300000014400f00c00400001010003403500001d0000000003003300010000f00110000100000000c300430c00100100103100330000000030303000010000000033000c300100103001003c000031000330000133000f0000010104004003d0000f00310000004330004103043c30000003010030000105000003030030000010000114000033030d000000110000003004110000000000001000c440010450350f1141100003001000004d0100030010030000000301000310000000010101300000c00000013110000030000000000007100f03000004010d40003000010000030010030000133100000043004000000000000c0004030310f00045010100000000d03001030000c00003104300300301033000000111003103c00031c00040000001001000041003030030010c11010c000c3000000000c303003f100000000000301040010000001010030c000000000c000000100300000c030000000000070000000000c03701001403010001313000130134044040300100030003000000000010000003100000003c000f0000013303033011040010000100000000004111001074000003441011100133010000033000c44001000010000000031001310d300030103100033000c00cc0000004c00404000300030f0000c10101030100c0110410104304000003413330000000070315003004030033041000000103c300000000000000000101133300c001010040400030300013440000007000030030103300040040001433033000130000403000400401000001000000000003010c10303305001000130001304010c01000000000000000000000c03030140731c0000000000011000010330c0031300010000000003011000d013c10000401010000;
rom_uints[829] = 8192'h1d003000001000010d31c03c30c0000000000c0007100000430000001300001c0000000c000c30700c00310d3010100003033000000003000110000304c1003010101000000000000c400010300033013000100401c04000010f01031000c0030c300000c411001400010004050cd41013034400c000400d1000033d040404c03000500030001040044700100000000000070f00030110400000001f41000310371c011100030d001c01003001c00000030000000003c0304330000410d0000031103100c33013003cc1000f373000130310d0000000000100010303c000000c140300300003410310010004013f3003110301000001000000000000030010003730040cc41130cc4000010330004000000000c13403030f0c004004c3c00003000340040044130010000c00001300310c00030c3130031000330010300401007000113300010000007f003000007c0440141300304fc03ff00000004f100300001000000003f300007d00000100100030000000d313030004031040001100000403000c001310ccc104133000000000000010c70c00300003300001d0031100c01003000c30103cc0000000030700c11003411300c3040000000cc00000730c000c003400000c0000030107000000000310000000003003300c33d000c13103010401c004004001300c1530003c340000100c000000030330103c010030c00000100d344f000700d003040343100000301003000d330fc400130101037cd005000010000001010003000103d100040c000411000003040000003000000000300030030310300003001010000c1000000100000000040113041df31330010c0100c1030030040c3000000000d103300101c1010000000300331000130cf000000000000003010010010130000000013c3000040c0000003100000030d00000000cf000003010301000d300043c000c0f000d037c0f300000000303000040030000040301c30330041c00000501074000c0330c0000331401034300000000cc0000000003000014170400030100000700103000001003041000c0011010100f0000000330000c000031030000000000c00c000000003353101000000c000dc37000100003000100030000000300304000c10030d01c0300110c000040300c100000000300040003001100003000003c050504000001000c0000000010000010031000004d30300371031000000000100010311010110000300107000c5471100000330300030401100004300013700311040000303100004030000000000000000000c017100100000001000c3001013001000100000000000df000037110030100030000074c000d0f30000303300015030cd03c004000000001000000000c03000003430300000d30cc01000000000c00413034003d000000000;
rom_uints[830] = 8192'hc054c000c010300000000007040001404c4c0000030c0400000000c10140000000400400137000000410000400034c03c0030c000000301400004000000000040003100000003c30000c0043000000030400000c3000000c001400000030003000040c0003100400c700000010c100c010000c000004100000403c011100000cc34007001330000100000000f00000000000040000000300400c01003030001000040000c300100000303003000000000000000000000c0c001000000000003000010003010100100400001f0004030000000d000000000c00700000000000000000003030000000010000000fc0010000d000f0c3000101001000400000001100100004011040030030000001103400470005110f3400030001000003c0010000003000000000030031cc1c3000000001040400000300000400010c0004100040d00c1000040000100000d40130300000400400300c340001031314000010000c003d001400304330000c0033d50010000040100003100004100000c000000700440c0f43000004000000000030100000000030000301000010c00000500000000c00000c0400000040000000100000000000005000100300000100000c000000000100000400000f00c0004000000030000004004504000000000030000000000005400cf10000003000c101c0044010004004000000000000001c0030000cc03003000000004000440101000000000000000110004004003034000000100000000000000001c00400000000003000430000000000000000104001000033000030700100030030033030013400303503000000004000c70c00003000030500000c00001010010000010000cc10c00d03040000001001000010400000400000013300000000000300000cfc30041c0404010000030400300010000d300d70001000010000030300304004544300104000000030000000100000030000000000003400300000101c00000000000000000004070c00300000100c3c00c100003300003c010000040004001000040000003100010400000000c04010c0000000003000010000000400000c04100300000130000c00341000040030000000c000041100000030004000c000d301330004000c0c30000000400000c000000003000d5c304000001300300c3000005000000004000d0300c000400100000030303010040034000c30000c00000300000c0004100000000000000410f00000100000001d000d30000440001000014000000000000000300400000f0001000000000000001000103000033000000000d00001d00430c00000000c0000040000303000000c0c303003041c000004c71000400c0d000c004100000c001000330040300400000000017040000c010c30010000000400000004000300000010411000c0000;
rom_uints[831] = 8192'h307000000000000000000000000400500000300000c0d01014000c0000040010cc0010447010000000440000003c300c0010433000000000300004004000c000100c000000004c3000d00c0c00304c003010000034300400000004100000011000000000110000111300100400000000c0000c000400003000000c04100c300c4400100010000004000004000410000000000c4704000030300ccc4050003c000030000000000c0014f430c010300000000040400c003000000000000c010000000000000000000000041414000c0000303000c40000001004100000100000100c30700000001040103000041314100010004c0000004000000000040c0000f000001330001000100430000003000030101001cc3400cc040c040000f00000000c00000000100c000000103004c01010400030000400c0000004001030001030c044000cc00030000c0000300c003030c0010040c01c1c00000000c0000cd04010c0103000001c0000000000343c30c030100010dc1c001000300010300300001000000000001c000000344400000000001c00300000040c400010300f0400003000100000c030000c3000300000103c000014000c00000030040c4c3c3000100c00c00030001050001000000000000010c000000070000c301000c0300c0000000004000010110400000004001000000c00401c700000000040100c3030000110040034401010000400100000000010003404d030d00c0c10000004000010100010000cc0000c30000030004000001004000000500100cc10040c30000c00000000040010cc00005400001000001030000004100c00000c104034301030000c403000103000c00000001000100c0010100000101c00003004000000000c300000001c041c00003c003c50000c04000c00003c30000040040000000400001c3000401c045400d0cc000040d00410103014003410c010300c0c000c101000cc00001000d00000040c30003400c000400100000cf000d03003500c00000000001404000400004c0000130014001c005c00c00000000c041030003000000000000000003030004000000431000000c000140400c00c31100000000c000c00000004300c0000000400400000001000041010003030001030040c30303010003000400404000c0000000c100d000000001440100000010000000050000c00003030041c000000003c30010c1010d0140c0c0000101034000004043c001c401c70100000000000003000000c0004d0100010003410100c00000030c40010101c000000100000040000001000000000d010000000300040110000001c7000001000343000000c0000c0000000043c0000000000000000000c100c4030000000110c001c0000c0d034000010f000003430003000301000f00000300000c000;
rom_uints[832] = 8192'h7441400001300001d000044000450010c41500000070c000001df0c103000000000f0cc00c0000c44c100c3100400c45df00000005c040c0030004000000000000400cc0cc0041c0000030cf4040000040004030400003003003f301004010440104153340c00f40003474003045c0000000050040000c70400000c00000111013c50001030f000f0000003400c0c053100000300f00000005d01f0fc00003003040000040004cc000c000001cc00c4000440000003cc1010070000f00c000031c1400c0001c40c1004c010000c303f014d01500000000c3031533c100400031cc400001c0c000000440030100705000403f430c40500000300040030000000000c1c0400c000040000504000000c4004150c503740540400000030005d040133000000c000c0000c00000c04f1303034000c004c30050c00000015400f400c4400001300cc04000c0c4004003c040100440000503303500100cc00000c0c0403003c10f3ff043f00440c00004101000400001c0300500000530013cc310c04cf5410c3340c0c0340500000fc31c0d0c00000003000070044000c00c430cc04003d010450000d000004000014000d000c0c0cc34304303100003f00000c34045c03000000000434100550004c000c00040c0000000140330014000014040cf0070003c00000100403130c00071000001004003c1c10340040c0f003f7010043c0003cc004400c00c00c40341d07c00004c001001c11003cc000f044710040000000c1000050ccf0040174040c0c001004400404000c00004c04c00c1400040c0c0400140103000040003030000cf000500000cc0000cc0044c00141110d4543000500005c3c50370300c0c0c00d410cf414f3c40000c134040cc0540400c003004540000c00005433f10400f4c047fc003c000401cc044000c31000530034003f00000c0c0040cc3003003030070003070100c010c0070404000103f00400003000043c100000000c00000000500ccc00cf0f005130f0c10c00c0c0f4c30100c40000000d0001f74000001500c040005400ccf000343000330040510403040cc0300500334d05300c00100c00cc57043400000000fc000504030c01310400001c00c0000440305530040301040c0d1500104430301104070004500d00140f00300304c50c003f0000030c11cc0c10440c0c130710043c0c00103400fcc0300c000003100c010000c1401c000400c000c0070f10000c0c0c00f00c00040c34013fc5c33c00000c50f3040000c00cf3cf40040000403404000c0030fc30c00c05355044340c0c300c0040100004043045007c00003000000410530c003000104c0307103f003c40f0005014cc00c400100cd4040410300c3c0000501c41c0000300070000c00003c10101414c40f300045c0000c00431304cf10134500300000c;
rom_uints[833] = 8192'hc3000001cf00041c040f3fc00704000340030d000d04000003d0011531c10000007403c37f000000c1000c03031f01dc40014c403cc43fc0030300000000030400401001c001000c000f01c00004c0c001013000113100000340000040033f04c13f00010f01000c7c5d00007041001040c4d50000c30144c3c00400001000cc400001004100000044000001000f000104300c003000003001000003044c00300c7300001f010f0013c000010100c0c31f00030030c00403000c100100013cd130003000000300110100003004300101050414010315000471500030700013031300040cd30300000340440400000735c700c4c3040040000030c341000003c103f33f0303c7f33010000f3c11c000000d03d00c301100ff0000313d0100010c00000030040000000f173031003c00c1000c41000c010000040d0c10501305410114000ccc0000033c140310000000304030101c3c03c000c5173c0010cf47000ccf0f4503000114033f431701114f030c3c00c0000000000cc3000c0c30000f00030500c4000030c3003040003cf4030010000300450c000000410133400100c70003174410030004100c011d05013c1410c001400c000000001001000300c3300000100100030c4410004001030004300001c0501030040dc300030c000d003030f0013000c3301c03000f0d0000d300715c0dc1c333030000303103cc0004007101000000100000140333000014000044c00d030c00c050c400003000c400000f1f0041000300004131000005c003ff4100000000100043cf400000007100310c0000000100000c710130540503010003030001000041440f0450000100c00310000d011004c103040f010000333dc10c000304030040330000001033000c0000c100000150c10010000005003f014401000044003c000f01000300410cc010311f00034101710405d7130000ddc0000f0c0f07f040c504300000104c003d000400000030070311000100500033000400001c000d043cd130400510140040000104040004040010000d000300001500000f001404000f3c0000170c040030000f00043000000d00004c004d1003033004c00400000f000003000c0c3003400003000100cdd51030c0040000030400137101010c040411d4000403014030c533f314000300000c0000004007000300c140400030004d000430001045400003300c1c3100001f07110305c400c300c03c000c001001503c030055014310053003100070000001c1c0101000430c03010313700010150000000301050c0000430c00004c00003300c31c0400c00101004043030c0000c041010000030100000c51030c000d540300000c0c03c3010d0000000411f00000c30000430703010000430300c401000304010c0000044103100000c00001700303c3334d04410000;
rom_uints[834] = 8192'h30c00000041cc3005cd0c0d00040104f70040430000d114c50c1f00300041110f000104c300701447c0000500000f0030000703303014011040000701000033000c0cf000c113c0000c301000c040c03000d00004733017000df00043c30301c040010000c101001300000113c100000030300c0304014007c04c00073130ccc1cd104ccc00000000c000100000c04140000100010000030100010c15c00c10010400300d01c34000303c0000c000000330c000041007010c000400f40c00000140c0003000c0c0000005000100c0c000000030010ccc0ccf70c1004f0004c100100014c44000000c00030cff30030043cc0001500007040000c01d74c0030100c00071304ccc74030f43c0300000400c0c00c00550000f310700004010400140300000040000cc001300007f00c103c00103300130000740304c05040cc1c003310300143000170c30cd4000054000c430000000440000f000dcc100040c14dc00d0530d3c04000103044f00f10030033401ccc300100143030f0000000101cd0000c00000005077400dc1cc030010000c0000101000000cc0430404034044c0330004d0f0c03000c00001030104007713500010400003300f04c000000f7000000041010c0144c4c000070000030400400374003400c00041004000031033000004000c100301000c033100404400cf0371c5c004000cf0000c0141011c30c5400d30c000000c070010c007100d410f0044410001c01000044000007d10100030f100c370304000303070c0010004000000c1040000400400430004003c0437001000501d000100f0004000c117c000c0c0001d04c0c170f03000d0c000001100014440c04c041104c343030000c07140000d0071451c30fc0000000d00c040400414001000c0000c000010d000000c3c030470003040030400030044100304014440001c0fc00000304034dc03014144004300d000400011000304100c0300001c000000001430000cf30d300000013307cf0c100003c300047c7000040f400000440000000000134c4031000100010d00d10000c0000144d00cd00d010434c0341001fc0104030c13c01c300001d04334413130000000304001f01d00003300014040c40c005000c01000c0c00000000300c1c50c01000000004c00fcc00030040000130440d0c0300030075310010710000c0007330c0000040000000c00400400cc0033030000130140030040004403400c003d305040000430d00d01000000c41000000040130350543500030c0c00014100000c30314440c0400c0000403c0040040dc00003c53c1001000001c044043001400030014003000c003030f04540041041c0000f0c37410003040c40000c00010000000c7c31cf05000140c300070000c3f0100004c1073000331400000000030300c4013710c010000;
rom_uints[835] = 8192'hc5000000033000403c043300040c0310440044340000000004014100105cf3c1000c043f0070001003c000c0130033c0310c0c00114000700441000c0c304c04430cc300000010300000000003005000c0013004f10d000103033c4d400400314030430101c0300570f10c007103430cccc0d0c0035300100004c004000300c41c030000003c0000010c00011100005731030000001000570040100140c030030300d40040007300c0401000114000140c004043000040d00071000c3001000000d0000000004f04017c00033c1c3400000000050040100000f0000041dc000310070311dc0000c0330c00d301371d0114410d0100000005000004000000000050000034000f0003000040c000300000d0005c5030404301300300000030c303000c00000cc0000003041f103140004100000cc0c0000400c0100c003500dcc030c0044400fc5300010040c3000013001f43d10c4040000100101030700300c0005000c000005000c00043030011003d00cc00c00000003303f0400073013f030003f100c0100c13000505003c3000df130000c001000303705034030003110103ccc000c0f400100000c00701c31c017000000f0c041305c000c040001340000f0530030330007107140330000011004010030c013040000003410cc0d314c7300037d3000030c0c00c44000000c040cc00003030537d431c0f40003570c07000c3010fc30040430000071400f1033000c00000300100c0400000333047010d10030c3033f11033000c00010310c431003c040030c303004f43c4d304001001010300003000c3000043c0040cc00001010170030440430001c03004c310003c300000c7013001000003043300400003c00070cc040373130300c00000d404400344300030000033010000300000c00fc001330100dc3041000001c04003c000d71f0c000100cc0500d010300300f3c0003107000300c000700053300040007004005001000000004100100000f10000001440337100c00c3000501001030100c000cc03104000050043f031000000030701730404430001430cc000f5310000c00c4001c00301c0010001c043400003000000010000413013c30f501c31303000000043103031c00101040004c00300304c0c050c0410033d440100400c0100c00003f0033003010000c0540f000c00000001530140030300040003031400000300330300000003404040c000000500c4301000003341030041000014310040cc014f110c000301310500430000001300000330c103000030cc0313000c00400000300000f10000c000c00140000105000407c00300c0310071030001010d01000310000001c1330ff00000000301034c001c00000300000301010f0300000c00100103010041015100300001c0017010000303000100d031d3430400000000;
rom_uints[836] = 8192'hf3100130300401000000c070003150f000004030001011000037035070040430300cfd01c400c0c04500c000000073c050000c3d00000d000400001001300070f4445000501004000001403000c04001413035c00000100040f1c0003c00300070cd0031304c0101d43c000400110000030300100c00c330c0000d10000000ccc14700000400130400100100c0c000143000000000000030c010000440c001c0300f713000003041033001015300c10000c14000d0041000c3c054c4c4000000400000000040c070000000113070000340013330c40f00404fcc00000df00cc00c0040000010000034105f101101d00303f0d30040000000000c000004003400f0c0000070104031f300041040433000303030000c3c040c0c000300000000f0c400000030000c4000003c3000c00100400000c40050030000000000c4401040000cf0000004037001c000000010c0f10c000031404030077c03d03003001100330010700030304000000000cc3001300c0004c034000033c1f010101040407111000003c000c03000130001013000500400400000300100c00000f0000404034534c3d131500440030001f1311300c03001304031037300c030000000313c10030071f434003000c0fc000000cc0010c3410304f00001043000f0d000c03041033150c00c3040003000c4c010003033333cc0704004f0c101300070000031cc1040cc0000c0c00005403104040000c0003030cc003131c0c000ccc10001104000f040004000100000140005000040004000000030404c0041f30000004cf10000c13000c04410c0700000030040000010114c7033030000f000301003301450c4004000c0d00030000c04000010cc40d000300441343c00c0414000000030003cc033004000d140304000c50304144043433c00104c0d00700000343010704000130300d41700003300103000140440f3007000cc00400000000034c000300c0000000c00c000300000300011c07000033f4d003c0033c10000f000301000540050c0f000303000300040030c470c0f000000405cc0f03000040c0000430c410100000040007c70001010000c0040000000000000c00c0100000130c0404003100000400c440c07400040003100000041c30f00000000143d1040c00c501000003c0000f040004005703c01f043000030300c37cc0f000340001070000f714000004cc5000003034000c0000004003040304000000311c314000004d40013c0c03010c0104f3301d41030003f00014100c0c14303f0000044400040c3c07001c000140010c311d3100c0000004c00005c00344000000000001000100fc40000003730c043c4f150100000000c300c0040004c1033301004301f501030110050c070003370c0f300fc13300410c0000030030047d0110d3000c01100000000;
rom_uints[837] = 8192'h3c30c00c0cc00000040010c000cc000c00500040001c700001000004500400c00c040340c4100000c5000400000050011000004404011c0c0400c0057000c400c0003300c04c4c003000ccc00000cc4c7010000000043c30040300000044030c0044c0c0c0c0c00c010c0000000040040c400c0c00000c000f30404100cc00000310fc0004300c00300400140030004044000c000304c05fc0300c044431344c000000047c003440001000404050040cc074c0000c04400044c040047c0004053000c3d000041000c00001501044105004c4c40000104404047004dc70c01c00000000004000c0d4000c4c504040cc0400c1007000000000000007f040c000c0400cc0430c440c0000c00c430100440400d400f100dcd003c000cc40c0401130cc300000c0500047005000c40444000000c000034041c00c000000040f033043c0000000cc4cc004c0401c04cc0000010c00c1d010304c00c00000c40050c00c1404d104c3140cc00c000cc0100440c004c4000000c0404000101c00000010ccc00000c0704c0c00c0000c50104f1c044004dc000000c0440010c0f000040100305cc0010440017000001000054030c04300040cc00c40f01040300c10c0c0c0c07004c0c1000c0400500c000c0c0001040c0000000cc00004300000cc1c5c50030c3000105041c041cc00400000d0c0301cd7013c04000c1f000000404000000003400c00c0c1540fc405c11c00cc0f00043400c0005000000413034c00c00040040c530cc00140000040c0001401c040c1c00000533c401340000c0000c0c0303f00c41c100c0404000c100f0401140107000030000000cc0040003c44c0003c300c41c001040d000c0c300400440030000000000070001043c00cd0d040c0c4010100c0c00c0c00140000c00c0000004f040c000cc0400000000000d40014f300d0700001f04000c300c54c000c0cc0400c00cf01c0004034d0c4c000000300404000000c0c0400c404001000003004405c050044cc007030004007404c00400c000053c000c00c0400c040440c40000410c0030400c40cc05c04cc00d0000050000000400c0400000c100400c4404c040c03001c040400c004c41000044c004400010400000100c000000c0040c0000404c00c00c0470011d00300c500c04040000c000c0000034100400000c10400c0c0d00043004000000d0010000c504000f433404004044400cc004001000410c003000300000ccc400050c0410000400300003004400400000c4000c0cf40400411000f3f40400000400345000004000000405cd01d4000004000000040c0001140c0000c00000c0c40000300c0000000cc300cc0c40c0c0c0000c00000c404000000011004000040440010001cc04114f004ccccd0f0c000f0000001c00cf0c00300000004c04000405c4cc0400;
rom_uints[838] = 8192'h104c0000003cd1010033300010000000f340c000103cc000000040410c0d3000c01c71301c110001000000010d00000c710300d00030011f313000003711000031051310010300001000c000f0c0c05000310010110000405d300f4140f3c000000304304000000104453400000f33c71010010300c4007000c003c30f0c03031dd30303031c00000c10100030040f0c4c300010004000000030300003331f1001c0100c4110f4d100000041403c03000340100400031c7000110033133c03000c1c001100001110cd0001300000010c0330000d401100c0f000004400100000000100301cc00d00000103fc0cc3010030011d01010c00000300d411000040000cc300110100cd001003000333007740010cc110d435ff4040040003400301300004000010000433f03000c0311d400011c00300c1100000300330013300d0001040c0101003040303000c4030f33000011c01000c0330000000374001030030f000334001410d0003401c014100331401033300d004c010001000000f430310117010310030003000404303100030300f000003f0101100010f10540130114100040103100c030c003410c000d10c0000303000c301033c0000000030340d0ccd31c101140f0101013004400c0103333c030010010003000141000040003d330c00c41001c30030100107400144404cd301000f00010d00000001c10100004010047034c0000c0dd1c00111070d100400100d057100010000014d000c001f33c4c303030000000400000001c10000340cc43100004010031cc01103c10000500404344c000040000030007000030000430000c03011d00d3000013c000330003ff1010075140000010330300000300101f04f0330000301100000000400000000000000005173013377110010140004307c17010000c340300041100300c013030110044c00333000c00003d300004351000300001001104cc073000300000130100c0000003000300100010000000410100040443d00330c14300500c40f430c0000003c000f0130c00011000c0c00304005404313d10031431c073d0f0104310c103333031c3100013413004101f001d30170030037c0001110c0000043c3130300103d037310004ccc000034d000c000010010300111100005330d050d710c404d0d1400010000303c010001433c0100003d30c03733011d000010000c030010000303400004013000313400f30000101030d13c301304010013000c013c000cd00f00004000410100070c4030c070500c414040030001003301c30100d10003010d0100103400fcc31001103040000001010100101001440300cc03150c00011003005377500047000c70050d400010000000034703d00030100001010007103000000301f0003031004000410113000000001c00040030100300414300;
rom_uints[839] = 8192'hc001000000c340070c440005400c044c014400c0000000000000000c00404300070c4300c450000dc300c4000000140000000030000040c00000400000000c000c04d0000400c7c40000c00000400000ccc0030000000000404cd4dc000c00cc0040003000000000000cc00000003c13000300000703001c0304003401c4000dd1000040000007700010040f0c0c00100004010000000500300403c0000c040101f1030501c30400035000cc005004000000400000000c00003000000000000040300000000000000d000c0c0c4000c00054410c000010004744000c00d0033000000001044001010cc000dc54010000000f000004c00004000000c0c0fc040040043034030340c004c4400004c30c441c3000100c0d000000000f4cc00c04d00300000770030c010001000044400300030c0000003400c1c00001004c0c00000c0130040034c4001050c00310c1004c0001000cc05c03c3030000014103c1000d13f00c1c0000c043044010100040c400101300cc001000404003c304471000fc11003ff4c0000000004117073000d0400c00c0000c0400004004000100404c014000013044004003300f00c001030001004010c0cc00c5c010c040000c43c03300000040000041000c00000000000c001000c00300c0f0c0c00000c0c00300303300cc004000c000c3d000cc400c04cc100003c300400003cc00000c4000000000c031c3000c00000c001004c000100000400c300c0000c000414c00040140000550000140030000010003000430cf100cc040000010100c100001c0040c0000100000040c000c4400000000040400034d000000000000cd00004043004c0300403100100100040cc304c40004030000430000040040cd01000400003000000410000400000c000000434f0030f00013140070004c01000030000540c3040c044d03000001430c0300000000c100040000440000c0040000000000000000100001100010000000400c00000d43030c0040000100000000000c005400000004500c010000000c0000c40300cc004c0c10000330000043000cc4c005400d0007c0001004704444c3000c03000c01044c40c040100700000040000c441003000c341000000400004004dc0000000000040410c71017300001400000010d00c00000c004000340c45000000d000c0d0403000100103dd0c00040c04004033f0000c04c00c00000004504100d40300040000433c00044104d0003f0000c00000140007400cc00000000000040d00001f13c5d040001ccf0000c0c0040404040100d010001040003000c0000000100100c0001011f00c000c04000400000300c300000d403f0000c330000c0c30000c00cc0000000c04040c404c0000000000000c000000000000103040cdc7000000c440000000044034c000340000100c0c40c0;
rom_uints[840] = 8192'h1000c00d00001034000c0010701030003003000400004000c0033034000000743044001030001000c00000040cc30c3c303003001c0303000c01400040000410000000000700000c0c0000c10c0d0000014400004004000300004100040000310c40010054004d10000000400100010d4000c10130430000c004cc0c0104000040070004010400000c04c0ccfc4410030000003f00013300137154001413040c0c013d0c0004000c000000034c033100000c0100cc0440000430000000054300003003000c0d00314d0000034c0cc1000c3000000c00c00000003140000404000000040000ccc4003000000050300c07013c000000400110000000000300c40034040d00300c00c1cf0c0301000d343c0c1040004331333cc0ff3000100100000dc00000c00010010c7000340c0c0c0000003cc0000000300010001110030000c400c1000000cc0c0300070000f000040c103041410fc0cd00000500101c000003000000100d03070000000c0cc00000000f03000000cd00004000040000d144430004000000cd0003c00d00000000000000000007000c070000100007c55330040f000f400d0c300000000000300400c00c00010f000000c00004070100300000004001000c00100c40001f0040000007030000010000000cc0000100100f04040100030d000130414130070010003140000c004400410c0c0003c00c04030704000000000140c03010040cc0000000013003d0034134c30000005c04c000c0004010c140000045077c0c3004000000000c3000000300000d0403c40c00d000003400010303c0000400005c0d00000400003000010103700030030d0c0044070534000003004370c3400007013000300d0000004000030001c50100100f000000004c000055cc00044007f00c0d0000000700010000000004000c040c000400000004000444100c0c40000001004000000000400f3000300c43400000141f030000000143010000030011000004070000c0c03003000030cc110330c00000000170000100000c0d300400013c0407000003010104000400003000000c500031000000030c0f3100c0443000c040000000040d00000514010c3010cc003100000cc0000c0000000000000000300cc33f00011401000cc400100c03100103440100000300000041c00300000010000c13c1143400000cc4000400030c4050c001030000410c0c0c0000000c100c040010c404070040040000033300000d0007010000040c00400c00c3030410c0050c0001000c000434303443c53d00004d0103300430f100010001000003017103000000c0000110010030030031300000000000030d47040c0004c00400040001000000000000140d3dc00100c1400c10100000070c0403000000010000f004340100300101500c0030034c0000300;
rom_uints[841] = 8192'h4cc00001040c0031004110c40004000300040305170001000303c10040001c0000c0c103000001000c040100000000430003034cf000070013c00000004300c0004053100000000000000000c0010f3c0c3001c0c000330f04030501001703010001003001050000003701000030c0000cc00cc0000033004103f1030c0000010500c10110430003000000430104c0031410000003000001050c40c303005000410000c0000000c01110c3c303000f00030444000c0140050f3100d503011000030c000d0000000007400f40010300000004000fc30003004d40c3003c73010000c0000005d0010000f003c001030113d0c7c100ccc0000000004ccc030103030000f0c001010fc100010d0010000c001c00000003033001c00003003100c00000c1000000330cc0c000110c7003c300000331001000130000c004070000c403000001c50cff0303c000310003c0140003300500040333030f00330104c00110433f304f5000031c130304c0000003000004000040010107000004c0444dc1000100010304010300070000c000c000c31300014000000035000000c300000000000004c1033010c003cc030cc330c0040000040003000fc30010000303300001000fcc01003403010fc00c044003030330000305c014000000c4c503c0c0000443040c000400000340000743f04000700043070f0503c0003100010300c30400010c70c50037003000001001c10000030000c000010303044000110000030150140410100d10000000c0000fc0cc0001c4d00040030317130000d3c330030c03000044c00040000101c34303000003c041c100000501010003c0c00c1c0140030700014510c100c030c0000000300103451004cc0140030001005000f0c3c30000c3c000000301000f0d0c37c30d010303cc00400003000001040c340003011c0410000007004000000d01c4c00000c030100c0000000703000cc0000010010c01000010000c03cf0040030001034c000000001000030301c0000000034cd001000f014000c003c0001400000c400c00d0004370c3c303000000fcc101000003c040f00001000c010301001000410000004000c3110c00cc01000003cc00c0510f000403c400000000c000000000d1010400030301000000000000070400400301f4000101c040100040010dcc10f40007000000004100c003000c00000304c0000c031000c0010034000c40c003c40300034007c71000030300011f7343040303f04300c000c000404104d3000030010007c03cc14400013cc07044c44100030d0030c04303c14014010f40040003000c40110f300000c40004d0000010004004033040045d007000c001cf410303c500030300051041010300010c030300340c300303c0000103c30c03000000440341000000034300c03004010300000c0;
rom_uints[842] = 8192'h1cc000004c4c40400000400403000010c03300c4310040040040f5000401c4400c0000d04f3040c001100000c040c40000300040450c00f0f00040000000000300c0c0000040045c000070500000400030c010413014d010430300c40000c0c00000400303003110000003000c1c0410cd030000cccc00d100430001c000000000014500500400c000000040030100043010c000004001444100000004cc00000000000000005c004001404100f540400c00530d00000011003f00001c00c000c004000000004000001030100000c00000430000000010000c14c7c0c05040440440000434cdc00000c000354403000001300001004c000010c00070c000003044404cc00004f00000c100000c40000ccc0c0c430cc000c0c04000000005d000000c300000c30045c00c444000c0500403303000c001000030d000000300c000fd01c0fc00d004000004000ccc0043004000000040f030ffcf0004c00c10cc4d10000130400003000c030cc00000c0000000000c000d0c000c4cf001c0000110404003300000cd000c00c0400400f0450000010040000313000300d0000c0000000040033403407000c00040104c0400040040014c00c04000013070004440c30000dc4c000001c040053400cf00000c0000500c03c45400001340c000303f0040044c040cf5000c05000000c7031000c0013c0c000000c00400000c3100c03044440440040000c1000100430d0430cd000000000340000040fc00f00c0033004040cc3d10010004000007cc04003500104c000c10000c11100000000010400cc0300c31c04000034000001000000003c0100041500000400c0c004000c0c100400000001cc00041005010f044c000340c5007ccc030c04000005000300000000000c0100c004003100100105d40cc00c000000004544c030003310010103010c00c00c1300000c003f0000c001340c0c3040000c3100040c000c300000000000000040000007044530c00300000c05c00c0101c4f03cc054000004f40400cc00100001000cf400c000cc00c004cd10040000055000040000000c40000030c004c0044300c700000000000c00400005004400000000000000003400c04f01003c031000045c3400c040003000040c040cd004300c00c00003c010c00f003073004000000100c00c000010040404000000303003000d000403003430000003400044003c00007000f34c0000c01000cc30c5f00000001300050d040400004100000f0134000000f000c300cc5000004035000341cc0503000c0c0c03d0140cc0c44000f01c0000040000c015103140004000f04000c00400c00010000303000c3000013f0301cf70000001000004030300004f300000c00400400c0f0c0c000c00010c00000000c50301440000000cf004000000cc0c0400dc140c00040000140;
rom_uints[843] = 8192'h30c0000000000000000000100000000000014000110000000030700000d40040000030004c70330003030c03c0000c0000000d07dd0004d0300000c004000c000303004c0000000040000051c00100000100004ff0000040c70004030dc430000131000c400d000000041000330100001000000030c30f500cf00d0013000000cc14000031400003403c00c1000010004330000000001401440000034f00410cccd00001000000c0000010001cc003300100010000c70004000001140330100040000000c0017000040303470c030000000330000c03004004510c10000000c0000000000300000003c00cd4010003004037003000400010400d00000000030f4c00000c47030c1010c03c000000040c0140000c0c3003030000005c0c0cf00c01000004000011003000c1000300dc033c0070003004c000000c00007d00010000c00000004c04040100c4000003041003400030001d00000000d3030004010000c05130000cc00c00400400000c001000000000040c000431cf300000004004040370000033000001000c40000000100000470000040000c73000003300404c000004001c3c000000000ccc05301000000010dc00c00f7041130400001333001c00c00003300000cc00d040d100040373440037410404c00c07000c0000343003c10010000100010001340040000003010000530003000c011000c001000c00400c1300030000c3000400010044454100000c0000003004300070000003030001c010000000004000010304300c00000100c0030010104100003001000c0f43001000000005c000310003400000df00040001c00030000c0c0001c1c0001033000030c0040000304040000304040000003100004000310c0003000c00000cc3400c00040c0c00c0104c030040005000000040000c000000003000000100050dcc000740030040000111c301300030400004001004c30000000400004070000c100c10000000004c0004040000000000c431000100330001010000000113300100040040c0c03300000310000000004d0300c410047000000000000f000400003c000103c004010110004c000030000340000000300001000010c0c0000304030c00034004003cc000000c30dd40000001000df000000000004cc0433cc3000041000c00000000000c14c000000000f0000000c000000c300100300030c00301000300401100000104300003004c300401040003300cd00000400100037330001f041000400000d0cc00c4c0300003c10040003c0c30000430011f7100340001710cc0003040001400c00040000000740000d000000000000003000c0000000000050400040040000c100003000c00c000000000c400000300411430133043001c000004000004030c003000300003000300000f0004c007000000300000000;
rom_uints[844] = 8192'h4000c0000c300030c0000000004003030301030303000dcc003d04004003cc040007c0000300cc000000000003000f10040403303300400c00000000c00c14000130f01300000cc11400f300440001044cc401434045004104c003c73000dc0003c04d03500000074c30301c04030c10101050f1c30410400c1c001007000000400cfc00c410000000000040013000d0030000300001171c1c0c1110cd03300c3cc0fc003307c00f0000004014000000413d0d0000400430300000000344000001303c0040003050030000c0f30130d700c01103400d0000c0c410f43011000cc00c00010000c30003000003403f0033000040c40001004003004000100000103c001c01100001c01c100003000003c03004c00000304c000004007034733f000100000040010c0303000cf00000410300103100df4c04000000010047ccc303014000cc007113011000003000130cd0f01d3013410300c017030304c0030440404c000034c35c410000500300403044dc03041100530cc0000fc0c01000d3310330d5004107004001000300c3dc01100f0401000000001c413c4030010c400001f310d0004000431100110c030d00c430001130c1000c01000040001c000f00c0d00430011003c0000c00000c4000000f0c0050010c4d0c01330000f0cc00c30043030d050440cc00c4dc000cc0000d500013400c04000c0c010c000000c0030000c3fc4fc003004050004034000140310400000001c0040010300374c014004c7303c00c400300000311040d00410440c07000130040030033000f4f000435040c00f30001041030000d40701104100501c0300070030000000001501140003030003c0000007300441c44000110c0013300400470000d3cc0000cf000c0400000300400340300531444c03175130c33500041000130f70003001004400c433cc0c4d001300c10c0030f443c00c070010c140003f0050000100c100100003f3700011440000000c0050c043000000030c0750111c00300004000f3c0430170030005013003c0000000d000c0c0033000c03c3c33004000cff11ffc00300105030c010003030001000000000c00330130f0410014000001c000c0c04dd003cc4c10100070300040004033000040f0300c1003c74303030d040c30040054c004000300003cc04110000cc00c330300ccc0300030004dc00c104074011000004f1100c0000c000300004000410000d0000c01000f031053c001330003500c010010311c000004f55c30100c0003000000004000f0c3003f001703030c44c0040003010070100500000c0c00413330f3000040440374004000474400000010001c000451040000000c30c0d030000300340c000000000c000001050c11000001003f00001c43350030c04101401c10000001000000d700cc3cd41c0c0041031030;
rom_uints[845] = 8192'h1000030000c1f0fc13c0c30307007300cc03100400d04100c00010000013100000c11010c3c30000c0000c0030000000100000300305000f010003001d3000000010c0100334040c0000003031000100311000033041cc504500001010303141100540f010031000000003005300c00430000133f0c01010c00dc300c0000000c000c401401000041010004030000000111100000040400c1f13000301f4c1434300003000403133700c3303c03c00330c413000000040000c1041c000000000d005000001000000010000c0003343104c40d04000100000000000c1503100333333303030300070c0000740f0001100dcd301100d3000031100000010000050400013f00cfc00043030003000100000300f00003011c033004c0007d300300700c0c00000000000c15070000cc030015100000c1130100000001100f350400fc0450000c04000000103300000c15103c000034043407001c00033c04000103040400000cc4034013103c3d4010000130000c3011031d003c1f000c3301000347041104c10d00110130000c040330cfc000031003000110100c4c00110000010510330c03033000700000f3400710053c000040107c100d0310040c0000003543370000013c310003300330000300030010013d0000c034000340001330010033000103511c3f0300dd00000131c01c07300104000300301300f100f115000d074c00310300003c010c3707001cd01d0c0110151100300405000d1c0000003003000370043cd11010001401000300010003c000300010001011130303010f0dd00d1c0501c410030100000c000004030100310330340c00111c001007113440743000001dcc0100c400004c341430030cc004000000c1c113030010000000330000c0c030c000000401034000130100c11000c100000d0000073c3000f0070004c30000001c040c001077001403405300000000300730300d001731003410013400001010000101013104000000000040000410040c0d103014010c00070c100c00000114004105500000017f0070000300001333010001000c5303070dc0301110301c00770000040001343001f703470d1403000001c030000000030f0000000dd00100d03c03300f001c070000000333001f310000000033cc010c0303c31030300003000100073330033007000000013430c00c500dc0df340104030544c430cc001700000d0430001000c00c00000007310c0c010000000001010100101103344030000000050000000014030400015f0000304d1305011c00100dcc010001000000c01c1400300301103000010004300111000000300000000034010003000400400541030030001f0400000c333000010303004c100301000f0d40c3c300000c030c3001cc0d1c300001010034401703000d001010d00c0cf30003100;
rom_uints[846] = 8192'h410001040c000407c30d3c3c0000430005000000c00c440c443c4f0cc0700000c34c0c1fc0c13c17000000cf0c14000c01010fccc001754c4c0d034c01040100003000044045000003015370000400510100044000000c10ffc00404c03001040c00c0040c0400c0400cc034004500c00fc0000c070f00000007010400443d0cdc1c000f0304000000034c03d1043c4fc04000004301f0c000000c40c00c410cc0c000000010040001014c003001000c1c40000004340c00400c074041000c33400000004c04c0cc13000045030c044f4c000441014000c301000101c0c4014dc00c000400000c03000f3c011fd7004003000003000403003400c0030007134031c1c40005400c30c50403140c0c0001c40cc30c3fc404000f04100340c50ccc34c00fc41340f5310cc00000001c0010c000000c0404c00040c00000000040531c070007000001cc3000f0040c0000cc000300cccc00c7c00c004c040c0314c000051fd0000300c1010c01400043c000ccc7c100c0040c0fc00100404300c0cd4403c34c03cc000034450cc00d00cc00000001000c00c00d010000010c3c00404c140dd7c0c00003040c0001dc0004400c40fd50000031c1c301c0ccc3003c400c43c007c0073000c4c001c01100c1710c00340f1c030000cc4c04c000c7000c00130c4445cdc01005c004434000010c4f30c0f00c000000c300c700013d144d00000f00c0300404010ccc144100c30300030c0000c4cd3300001101110040d0c005030000c77100030c0f0c0040053100000c0000350c030400cd0003c1000004144000100d4041c0010000c343f040410400c1004000c400cc0c10003041444004d5001343100c030cc0003000c3700000c040054000140f100c40c700c005cc0004000400174344f03c0450cfcc0c005001c0dd0cc4000f0000cc0c0000000d0000015f140c001fc10000011035cc40440400000000c40007c000000cc3cd0074000000ccc000c0300013d00c00000c000c010cc1030003f50305c13003000c4cc400c000cc04c0000400003100013f10000000c00dcc5c0003304f0400dd0530041c000ccfc00c400000c00c0c4040310000004300ccc00100000001f13100010f0004000440003d0cc0c4c0040ccf000304f4010c54c300430c0000d4034cc3c0d0040f47034405cccc0010030d34c0c0413404c0040c0004c00c00000f0cc0d00110040f0001000c04040403c0000040030ccc000000000c0d001c431c43c000014d000f000105cd0000d4100c00304000d0f00f0f0c000cc30004c001400c0001400300c505c040004001400dc000000000140104c1000f000c000403c100cc0c140ccc40c43434400001c0c0400c0004c30c40033130140301403c1700c000400000047040c30c0c031404c00003000040d0c7001dc4000c0000c;
rom_uints[847] = 8192'h403c000070013030dc0040000104f0007040103000041c0150c00f00300c0100100400c00c50d03000400407010030140f0003dd0300000004000434010c040400c01000c100cc1c14000c000000334c373003c535f31c303c0330f00c401c00000000150000003005444104000030f43010010c00140c00000c4030041cdc0c0003004000303014004c047c440000000001d0030c40d000c054051400f0000047cd111004300040004001c0c04f35030004c547007000503000c00001d003000c003d003000030030000001c0004100433040c00533303414f70c1f144c001003004003000c0013400cc004400cc1304c04000000003010f00c000c0003c33004c0f30000f1300000070370fc100c0000c000cc3fc0cc105c40000000000c000000100000000000310440100417000f00100c000000004c3030d0001c400040000c0f003000030cc00c01c014000000044c0c0304c75fc1303100130110d0305000400d531401000040505000444000f4350010317cc00c04347cc00d0c1400040c4000040414430000c4003000303000c040010fc44000570030401cc400f1415400c0c0c40304350300103f01400d14c000300704c410000354001000100045c440c547447c0104401410c40440013540c105044c013034c00f0f00c0cccc40cc03f7fc300130f0033004000000f4004c01310010010c440c0000140000fc0000100c0001c00c40f0007000130c40403dc0010cc4c031305000010cc04500010010c41010040001104033fc3000000140100c40104000000044000103370010f04004040c4c01001400003140d40f0c1d3c0c3541000353d00c0005000410730030000c3000500c0000404431f00c03433c0300005c0304f00503000000040000500c004c040435c0300003005001000c0043004001000c30170c1403c031c0170000f10c070d030d0410000104c040fd0044003403c04405300d50000d1114004010010c00003040f00001c00d0040fcd44c3040004340540030030014010400c03410030000000100cd0cc04c05130000f0f400c3c0c400000433003010f0000c000000000101000030c10030c00030000310000047c050c30410000001d0303040c03f000300c030000403015001c00000414030c00040340cd40c0701000c3304171704400c000c30c03014f3043c000110440004000015f00c00101303000c3300f003010c30010c403ccf700004fcd0fdd0000107f431414c04c5c50500dc001400033c104340d070400334d0c30c00c130130010fc01cc1000031c01001c3305c0c03d403c100001f10c00030000000c0cdc00000100314001f00003c00304000c000c1000100c00100000400130f1400010c00c04343104f00000c7c00005c03001c030043005c40000005000f1004010111430001000;
rom_uints[848] = 8192'h300000000000401004300310000040030c40f000c01c30000c04030d40c4d030c0c7055040300403103004000000355430c00c70400c5c3000000011d0c3300fc015c0300c0c4000000c014f100c100c00101730d3400433030007d00040c000c0000c0404000400350c0000470043341000010300d0c400003070f0000040013010c0c0340000c404c0000c305004040400000005010c40c4c14104047000f03010000000003100000040040c3000c040100c000c400303000014c70100000000c000005000040303000400000fc40100f100000040000004030040001040103c000c300000300c03c00c3c3000540000701404003000f4030010041000000400040010000400000030f0f0c340330010d00c000f13007150100443c00fd0c000c0100404d11030000041000003000400000c040000000040004000c004c401500000000001c0c0000c100c000000001c11041f113133000c007043000000400c304c030010140100003c1003000000103001007000001710004140344000001005c0403430040000340003000000f10000c100c00004030c00041310d1c400143c000c03c40c4400000c30cc001c7010c0101c0c101433001470343010130d404010100400031c335c0001dc000c00004c34c43000104000f3700c00c003100000c000c0030300c000f01433531f1100110f403d70300000130000d401c00c0004471000000314000300000c3df300cd0054c01000c0031017c3c31040c004c0c000041400000c00040c1430040003f0df0010000400100c300c3c400400007010300040135cf05cc0040c00f0000400400000000000031c5013010130100034c00c501000070010030cc00c00000004f01f000004f3001000000013153c0000c1534001000014440030003000d4001311f0c010000c0000033000301070000350000010040000000d0040c00000100030010030c00004303c0000c0000c0040c0d00030004434001000401000050000000010c3c0041010001303104013f300030000300004000c0000101f70c73c300c15705030000000140c734030c000c040cc310000001c000000000010000440c0003030000c00100000001010c1cd3000000c0300fc110cc00c1041c000040cf0003004c0c1040c1001c03c003014040c140c0400103050300c031000000000000303003000cc4c0000030111400400400300c00004003c000014000000000401f0c0c007000334f00000007000f0f044300000004005100c03c000540043003c43dd000f0000004000c0041010d0001c500000301000303004fc000c04000f0000101001c0001010000010000000030c350010040c000007000103103c4000001010001000f130300110c0000cc00000f000000c04000003000c00131004310c01c014000310100300003000000;
rom_uints[849] = 8192'h31000407000d0c04000c0001070000000c010300000c040000000700037c030000000000300c030405110005c000010005030001001c000d01000000110003010001131c0d0004050300000000030400010c004cf1c0011303c00c0000010c310303050c30040010000c130c0001000c000f03040303001301f40c04010c3c04f5474000010f0017000f001c00040c0000010307000000000000000000010c1f000c0033004000030c03000c0045003c0107110100000000000000000f0c0001000f000401300041000c010c0f04030f030001000001c000000f0110000f300000040000000001010d0c130d100300043c0f0707300000000c030400000c003c0001010400f00003100c0c100f340000001303330004010303310c03010700c50010000000030c4d0c000c0c3c00110c040701000004110001033430100300130700110d040000040100041f0c03051000cc030304000047330d4411000c001c0104130c0c07030c00000d0c0700001d0c111000000d0c04000f00000c0c0004000f010400030301000003440c040057000c000c05000d000100010c01041504000f10000105100003003010013100000f041505000d0000004c100001000014040300c00030040f00411400c00001040d00010c0000000705c500000003010700000104000001100c0000c00c000c0013000c050304030f000400000500040031110c00340000000701040000010110000400003c0003003000c40404000000c5000c00003c0c0000000100310c40c0340301000c101c10030d04004c00010001000c0c00000c000303010001371c03000f1000040403000300044c03035103030401000043000c013c0c000c00104000000310133c03010003c0000c01030400000c0c000000000103050c000c3000013000050004010000303000000d0d00000000cc000010010c3c000501000003010f0c370c0303c000000004000000010003100f01000c003004000000101c00000f0400c003c1030410000cc1c10f0d1d000c003d00000704010d3003030000000c000cc100050031000004010f0d0003040403100103030c00001c000c0300400000000fc010010315034c04030000310c000031140034003c00000100030004003c3c000407051f4403000511140004000c040300011007040c050c3c0f000005000d3d00030004340d0000030c01000c030100040c11000000000000030004000130003f0007010300000c030c000f05030f000001041305000300000700007f000f0407000300030501000f000400000404000101130c0000030d0000d3000f0d0c3c04010100000300100f1c3300000c040107030000000303000001000004040000030ccf040c400304040f00000001010f0c000d0003010c0f0c0100030c0100010310000430070c00000f00;
rom_uints[850] = 8192'hc3000000f711303000000301003010c000001100000000004040003700040310103c00d00d0000303100004c00f0c173703010f0cc3c03330000c0f00001000030041100010000c000330c000003300001000410000040504d173340303050001010d4f0c000403003040000300410301c300030014400000001001503c000040010400c000040400000103033d00000040010000303001134110070f003d040cc43003344c1cc10400001c033031430001000000310f000000033301000004010037000000f3000c000433300403003f00001f04c0430f0f1300f011c30c30003100005000c33000010f73431000c0430304030d3000140000030000000cc0303003f013030005010000000000000003043d0010004003c040001f104303100303c000000c0c00101d00030cc0344400113044130f000c1104000c10300300000303400103000000000101000003c00100001c401500d0d0df0c100000c00000100003343c400351001007cc410c7013070000000c03330ccc0300300001010c00030331d0050300001004000001001000310c000040c0051044000100c540003dc500004003c0000410130c0040100100040103003000104000030004450cc4440cd00000040c3030f00d0c0c3000003014c137010c00003c300004000000000000d7000300034053100003300c0c5033030040400f0ccf000f0403050001000007c000030c000c0c0f0000c40c4001001003000c303300003700000001030710d00f034013000c011040000c00010000000004c444000017000c10003400c00c0c030000000300043000001c5d0c4103c00c070c00003003000c0c01000f10000c0f70000040003d3d11c0005c030401300000030030f000c00704341000000000000000400c000010010d0013031c50030703cf40000400000003300050003300000c03130000304cc0c1070010000110c000033000c00d000c070d03dc000c00004004000cc0000000cc3c0000301731c03010100c0043c033431100300005000c3004000003c011330000170043040cc000070000f0300001cc04000510113c0d030001004000000007c00100c035010005f0003303500000000010c47410100300c100400000000000000c3340000400030053107700100033731f37000000000003011300030f31fc000f00140c03fc3110cf3f0303300000040100040030003c00001010400d010300070413700300000000070700000015d000040011d0000000cc440030f00300043c050030003344fc03030c0c003013cf00103c100000000400000001050100030070110000cd10000f0070003000050f04000040030cc00c04c40cc1000c00000030070310004c0d00100000541400030003413000003d0030300c40010004430001c0cc000d14001f311c0001100000034;
rom_uints[851] = 8192'h4c0c000000003d137000001010044c1c040d0c30c0353010047030c115c0300004010cd000000ccc034000c0c0030070f40d3037003311ff74c00030001000000000370cc0030173000c0041c040c00c10000c00c01c3c00300fc0c3040f405c133010311005000cc1c000003010c000033030330c4157100374cfc03070103c0000c300003000400cc0014370140c01401000d0000c0c04f0c50100c350c0ccc0c01c0dccc040c04530d1c3f473737c17d01010004c44c0014f4034f0340c0c303400d7c00400003f00004c40000c01704c33700710d1044300303477300000000004013043030000f03770df03033c40c10dfd000004f1c03041030100030ff5113100040d477415fc0c3c00400c00d00030c3100301301c03c7103fc0000f10300000450c00300c10007d0c0700000350401c00c0003400003c0470f01c700cd004f0040500540cf1100c1107300c10cd000c40c003047447c13c00034440000c03043030d0c45fc7f434100030cc00500c70400035c37c453c3000cfc0010010740013330c00004000c0001c503400000c04c0013c00000400c0005005040f700400c0c00000004040000140c03c300f01cf0d0c00001dc1f404000703014f401011c00000d000cc0000004040044000003c350010304f0c000ff0400c70303c1043043c03401c7070c0004c431cc000c04f4c500f34001cc00c10031c3000c333c00000c3c0d41c30000070c050c00310110cc31400ff400cc7433ccc0f0d05300c0c0001300045f04fd13000400000044d07cc00c00000103c44043300040f00310c004040c000c07000cc440c0c400004d0c03031043c1030303403404c3030d340c04c0f0c01c700c00434c0007c0440c31c04f0d03cd010d43133c00000007440003c0004004430004000031000000004c040000000000c030140004400c403c4300144740000011440405cfd040010f100101430707c00c0000000410fd000400430030cd400000cc07c1c044054041dff000f3d04040005c0f00d4000c004741440400034cf5c0430003c0003c1131001400c035c03310000cc5c03004c4050000400000044000100300d0f04d4000c00440f14c004730f00c40734f00c00130000d0001070440cc370004c44300000003101c1000000c33c43154cd000451c0303004c303003110400000c30c740400014507c04407740400041c30314d00031037100000004cc043c30000073043047f00ccc700c0473043d0c10111130004c501dc030cc104711710001d50300dc50000c300003c005c000003c0c0ccc003301440c400100000f0f3104333d10000c000c3cc00000340000000100507c0c003cd1cfcc00010d1003f00000c04300400c0c3100c0c00000040c1000c00073cc007030f400100400f040300075c01d440f140470dc0100c1001;
rom_uints[852] = 8192'h313000003d30c5c0cc000000c400401044030000c00101d00143d10000030000000f1040070000c0c105000000000001400301c000330c100340c0000000c5011001707340c040004000cc41040040010001000110c07c0041d030c40010100cc0000301050010000c0041030500010100433300c0c101300004000c1000000004f13000000000cf000304350000404001000003000043c04c4c0c00c04030040007c0000001440010c00cc0000304004030410000305403000000041c0510001333c0f3000010004013c00000c0c30000c044c303005300c3c000003530000000000000f01300000000003f00f000c00c0000c3013000d0400004014100000000fcc103cc00d0f0f4000031014000000150d34000c04c30cd010000014010d4004500000000010300001140000040c1300040000f015c0040cc0c1000000c00cc40c44000000c0004040f00c0404f5005000010c04d0300070330310c0340100103c000030cd37403c003004cc0d040c004c001000440001cc000000100300cfc0c1000f043cc00cc441000c00335c04000000000014100030000010001430000d00000c33000c00050c30100c0000000000314f005c140f00035100001043010c04000f0000310000400000740300c03000000441000f000c0104030000301030030314c10c403010000010101030000007153c01010000fc01000011030310371f00d103100c3004410000c030001014c00540d0003001040070300303000100cd300404d00c5000104300500400003cf010130f001c1fc000300f100c030000040100c01000000c35040004000000105d0c0f30ccc1fc1c0c30300045011d400c0c04f3001c300300000000000c001410011004c107303f00f0cc54000c30014311110430000100000c4430030cc01c47c4000430cc3000001001000010c0510f0c0c0030400c00030500431c00300040100004004101017c301050303700010004000003c0103410003000001f1000c0f4340c34000430100c740010040130000c0400100c0000000003000100013003fc5c0040001c03c0000d340f400010040000f03c303c4000101000d0000013000001c0001000170004003000000440f000043034400d40331c00000cc00c000300300c0130145000c000043030c500cc0c33010f004010130040cc07300c0730003134d00400cc0000c00433c001300f313000f40044310400304000041c03033434004f00c4440000c310001000110000500000003c5040010140cc001c30c0000f001440040f00333040c001000f030d030c043010001004047040111000343103100301001300000c0400100c04000000f710731c00d00c350d5033010c00cc0031140cc03403140c003314c050700300400305f001000c00500400040000000141030401400c10030000100;
rom_uints[853] = 8192'h143c3d000300140ff0000c00000010c0000c040410040c04d003cc0c0c0d413050f040f004d30017000c00cd004c000300400010000c005004c40000c700f0300004dd10043004101000c00c0c0000f040470010043000134304d000400dc0c0d0c0c3040100404cc0000c04c000011400d00304c0144030004000d1400c00d00c040030315303ccc0d4c00c3400c401400c300000001040100500004414001010004100041c43c0100000000c1d0037400d4000000c0000007000111100333c00dc01000000034033130000400d10030cc0000c0cc44000c0c4004fc0cf000410cc00000500000010001441d4d00000410c0f10000000000c0000d0d30401004d001111000dc43f031c1dd01003003000035d7300433007c300000c0000f00030000000140f0001d400041330c030000c000c00c414f0400000c0000d04c01010000c000cd0d70c70113010300343000054300400004407c00c400000d040c0703003004d0c014cc113d0c0f7cc03000000000c30d3000050dc0cf4000010001f04c30c10140c4c3001c01dc000f4000700001044000004140c000000c000f0cc0dc10004c0d040003c00100000400000043040103300cf04014310000f5000000d0030d000003c0431f00007000cd0370010100001303fc00000010500000c005d0040000100f04000043704733c00d0304c04104000c110d00000000010c3010044c4c3401004c00100703c0010000000c5443f0104305100734c000d0740000c00100405000c04d0d47000004133010000000050100c40c00c0440001df00c077014104000004017400c00d00dc00c334f013c530300fc14c041c10000c00010c000710c700440000007100000315c00030000131403000c00c0c037000cc0703000000000c0f0301c10c400c010303c0010030d0c40301c000030001051f0404000000000d00310dcc003000fc30000000345100c40d40033d4704c00033104050c0000c00cc00400c0000c0003100044c0c3004c0100000c103c4ccc0f000004403103333fc0010400400010503000317d000100000000540c0010300373000000f510107c0f003000c100004040000034000303000c51100000c010005d1000000c34700c4000140040cc1c000103400c00fc500000ff0400040c103040c434031cc44cc7301401104c01043000044005040c0030d0c40c00104c430c011c0430000040410030000430000c04034c100cd040000000000000f0073001d0004c000c0000c4430c04007f300000d00c4000c010d400d0c0d000044000100c040cc310401400070001010000103c001310c3040000c0000010000c10000341000c30100300d01400c0ccfd004000550000300001000c50c30000c40000340003300000000c343040003003c03fcc00000101f0040340004c040400000000;
rom_uints[854] = 8192'h5300000000500300c0c053c000000104100040c011000300005c30033374300003f030d401000001001000130000d4d30c00cc4f330105303030030c00030004410140010000705400030103f0000000010000c503300101c30030c0000f00000030034003000100401f7700001c4001100100010001c5004400000000c4000c40014010100031000070c000031130303100c00000c00103c00013c1c00000010000000330713405c0000000d050010013130000001500000000001010c0000000704043000c0000030010403c000500003d10300c057300133000f0c343040cc00000100430430043000700733300303031000000400003003000033c0040001010400c10c0330004001c333033030c001404733013000f000001c00030c3f000cf100000000100003003303000c00000700300c00500050000000001033033000003001010d004c003400400000110035001000f3c33300003f0d3c0030040100300007000344330004040101031000010c30c4040000073001000034000000000300d013101030000c04f1300c13040010000000003100c1103c01c0150c0d3114c0c0300100001100000000070003003000030300000400001001310000000300005000011c041030004000013000c051000000403d050f0005003c0c10c30000040010033103500303003c0100000000300c000c003c0100300f000cf000040000cc0ccc3430504134000714040000001130001c01430030031c00cc30031311000c010304000030000d030303013105004c041411000f0030050000d0000c000707014c00000dc0c10040500d0c501c00000007030000000403450030dd0700330c0030000000300334001c303001300030000000ff03040000000300c05f01400013000f0c0c0010050c31f0105f04040300040f3030c303c00000104334340c0000000cc000f4001c013400c0030d0000003030000401c0001100c000005010000000003c04003000030d0c000c0101304100000c0004f000001300030040043c001030000000101404040050010414000701003d0013003d030500000101073c3703330000000c003f30001400330000000040000734000dcc0000310000010130030c0c0007040030100000053047100c000007340013070400030011301c345c010c0d0400335013f40c0f0400370c110031c33000004d030c007000000000300000004cd0040c000330313400311053000004130040011c300051003550000003000c00005c0f013033000400010f0f130c1100300000010f30f300033f0000c70110103040034303ff0030001c0c00f000000c340003430c30005004ff000004c004003c0c1c000000303300000400010c30000030033001110c0100015000c010030330000000c3000c03000003004c30100d0c0530000010;
rom_uints[855] = 8192'hc000000001c0d00004c01004000034c0c3c0054c1100004501000d000154400c0010d04003c000000000c7100300d3031c40000070004040c300c1340347c3000fc3343443047001010003cd030001c7440c030447c1000c4344300700110000c5310407405300000074f001030f05c00fc00c15000c00c0c0300001430004cd34041300030cc0c001c104c000010001c003004000030374c0544d03c30f010003030f0340000f0000040044f0f0f0000050040100000f0104c000000fc340c0c0cc04414000010013f000c030000300c10003c1100041031f000433c1f1c00300c1000007050043100500cc01c14c0110c40f000000000001000c100000004f0c030000c10c140000cc01c1300c004c44c0400000030040033c0030404c0c7300c10000030f0000000f03000700c0c00f1000450030400003010100110000f100000000000100100300144c540c014000003000c03440c0030043c400c100000000d300130cc00c010700054004d430003344c340c0044cf500c0010030c1001340c1c00c04000f330000c1004133c5040003030003c004000000001c000101000031004513c000001300030107430100001130fccf00c000040c04cc03400c050173301400c43f05c0c40343c0030000c004000010c543003300103103130c0c40040d4c1fc50340c0cc3010300001030030d40031130000000004c0110f3017413000053004140330001401000105c01c34c00000c30c440305c000c1c400000000100c01c0c000f3f14c0700d003004c030004cc0fc01700cc00010103700f000030c00040c10003703cc0f000c34001c4015347c130f0c00000c10000c5c305113141300103000001430c0401143fc10dc4c13000cc000100400001010c000301c4f000000400c1c0c3031104004c03c1c331430470004301003073c0c1cf104141400000c0c05000cf1400c4c37400c00f00400301000000000c0000001d0030000000c1c03001000003c100400000010305030cc04000030330c304003100000100c0c30fc03003414100040cc003411370114000000c00c40dc14c03c3c0c0c01030000c0400054000004500df3c00000000000000353103c000000040c3030004c403001140010000c001040134031c03430040401031c000500703310131dc40c340d000d000c0050301010743400704c00101c330c000104143000000040c03000000454700000000c0011300000c101001040fcf0001c0034f010cc7000f0300000000000303c000cc03041003f34035c40001000700c07d0400c0050101c10000000400043d44010c0100010007cc0043000501000001c130000010004f030371040100000c3001000d4c30040c1140d01005000c73c0c3010c400043000300000407c00100c4c00d03d1000004040c300300004001d300f003;
rom_uints[856] = 8192'h30440000300410000c000003430004cc300040100050300000cd40000400110100100c300001004000110000000c4000050c0300000501d05c0101001100c000c010d0f000100000c0000c00100000000001c000c0f0c040d000000000f00000c444c4050000004010000400000304c300300030f01010400c000000ddf304000dcc000c003c00400c0c00000000140c01000000000030d000c4100c4000000c7000000000330c0c00000000050c005c00f0143000c0110400c1c000fc14000000cc005000010f0c0043001000007c000004d133004004c000d1000403f300cc000f040000100000000000030443003c0000300040000010cc10003f0000000003004000003c400000c00404c00010c010c030f40040040c000000c0404440cc10c0100000c04cc1c03000000150c0c043010014c01000300000f301353000001000300430003c00c4c004000000000030000000c4c0004400c00c0000303c0030005cc01c0c00000000c000400400c0110c100000c101000133c044101501100c00003c430cc0400000d03000103103cd0000014000c0000000100f00400c0100007000540000100000044030f01100004001000010000c0004c00010000c40300300000300300c00c3000005040000013000f0c0000740000c1000303070cc401040cc00000400003100113010004311000c0001000000f03310000c0001103040400c4034000400000370004c0c00c00050300000300030001043040000403f00dc40000400cc00003000c000000037434000044000004000503000003c10c040404c00000540040c00003000c00004104c3370403c000030004105c0d400d0000000140000c073cc0fc10000040c0c00003000000c000c04010000100100c00301c000310004c00c00c0c030040c1044c04c003c00c400000000c0c03004d1000400000100000000c4c000304c1f1000100000000001c03000400c0c0000301040c0030030300001000000c000cc000000031143000030040c00000c01000100c03033000000000010100030110f0400003c00030000001040c00c3c3000004044000000001000000010000c0050430000003300c1000cc74000c0100001c00100103000000700030004700000000001001c0000000c1573000050044c040c404050c4043040c04cc000000000400040003310f30c0f0044c0000c3003c0000000100000010c1c0400405000007040000004c03130003000c0000040000030000010000000145c0c100000000c0cf0000c0004035400c0004040d00c00000004704c000003c10000300000300c0400333010f00000000401400000303000c000000c0000010c0000cc30000f3003c031000004000000401004c00000400410c0d1000c100ccc00300000c10000d0c00c000000010030000000010c00000c;
rom_uints[857] = 8192'h50700000003fd0c170000010cc0000000414004c501040000004c00010300c003030c00c00010000001010000000c0747010300cc004d05c700d0070300014000000104300100c400c00000030000001410c100c7c0000300010c00400101410000f0300c33000000c3c70000130cc400400c0403cd500f00c04503155000400c010000000000034c040003004c010c70403000f003004103f000400044000154c01d000100000c000041000315003d400fc1c0c000c00ccccc40005cc0744033043003030000304004c0004303c700054044001004f030c00010100030100c1003000104000000030301010011c00d00400c004cc7700104000c0c0400000001000500f30003d003f4440003000000c30c310c04000033c3d3000300c00000300010c0000f00cc000101c00c4c000103014000300100004c0000c0074c03cc0040c100c414f00044410000dc40030c0c00c0000400c30403710c00c000004040013100c00f0c1340110000c1000d0000003400c00f010000000f700103000404000700000030400430000000010300730000000000000004f531140003003030f01003c0c00000000340010005c0000c303100003c0cc170000c0100000001010c41c0d0000030c1000c0000c00031000700004000300400000c00c0c07140d00100cd1000001000c0004ccd00000000d400014c3030000703c0c3005100003d00000000003040c303300c400100c000000100000004004c004134000305400000010000c050001100440000c00300000711c000000c04000d000030c00470cc40c0000000c301300c00004000f440400c0000004000000010f030000c4703000c50f0c173c30c0000010104c044010003300000001c010003340000010f03303140d040030100034100400001040000cc0040000301403000c300c114053040534300000043d0000370001000300070c074c03403c3dcd00400000f33000001400040414000034f10c00003040000000f0004f04440440c03100740010000414004000400000000cc0410300d0000cd0000000031000000000540000003f00040f04c134c00077c514004c00333040300000104c000000d00f003403400040100500101040040d0153000c000070004011c004007304000cc00c00000c000000fcc03703010c140011331f00c03c040c70101003500004343c000004000c040000031c3030000004040000cd0040004040404c0034430000c1000410100001001010040000000005f00c01070000110000003c0000d000c0001000d5303000c0010dc0c050c03c000000f0037014000073400c300000cd00c00c0040473c000000747000403c1d4000333c000000001300410000c0401500000c0030043034010c000004000004100740cc3000300044000c3d0030f00407001c1300000000;
rom_uints[858] = 8192'h4d0000000d1f40c300010d01000700100c05400070f40000340700134d00c000c040f15101003c03100013c17001c111000003001cc34d0000c0c44c00000043301100307103300000303430001101c0010013c0f0cc0070c130310040110004700cc041cf040303c0100c40dc100000033010140440cc4c143dd40003c100f300c000000f000100d300001303333000c0010000010000001c000031dc30103140003000031100000040000c00004100cc1c7100307c03c3130000fc30000c100003113300504010103041303400310003404300f0103000031040001c010000040000ddf03000004c003d0f510c17104033050c13014101404337000003300130000c3cc1033c3511001340003003d00dfc0003000430fc3030c3cc105f1730050d0030000000300000330c0c10400010000000041300300400135f0014340740475031300004c1003431003001c0fc3c00040c7000340100c40c000c00173000410c03400004c00431010003100c000003300c104030100d700041003000010fc0330035000000411000350001c0d30000000000c000033050f133010c14030f0140d000004000000d10003700000c000441c00040103f4330001d00300c47507c003000d03100041001411030470100000d0c04150000c000c0d3f17103043100000300133430f045cd3d001000d01c0d50c030300dd000003c474370350410113003010007000010101f000c00030343100f00700001c00000d013300400007c40101000034000010cc030c3033001100001010c0000310c040000300300c500001331c0140001030000300000500140100030001014f3000410004c000d430337c0001007300c04f4310005c0f000013000c4104503430000371000c4007d0f00c4c010c000013030c300c3f00c1005301cc0d3cf007113001000000170c41010c0301f301f0403007431103000150c0030c1300000144c310c00010000000300000000304130000031cf003401443403173100013d000c400140074113000c035d00310000433003030f700c170003010043330c313001c00f00330030300005000040c700440440003d0400000437010000030c03c030000100000040000000c0530003003d000010013c000100f041000000f0cf74103033df41cc430000000300c40173453c103300c4010c0000fd030000110003030070100cf005000000c00000d350000730f430400571c04000003015141070001001013100c1004040d31003100000001000300330400073411000000013303000300c0304100710034d0c04001000040003c0330c34c1004f30001700100030001300130100010004304110000000400c0000c0100d00000010000003d13c00ff003030f0000040c03433001001f30f3400001030103000c10013dcd0c433050000005400;
rom_uints[859] = 8192'h5035001010004fc037000c7d4144cd03c7000000131c0c047c535011d4310403c73411fc3000051c3c03d4030c03040304c004030c01c100300c0fc10c0c0c0d01333f0330433c0000c0313c015c110c0001c1330d03cc4c001cc10030000f04070d0310031f110101d7000c04cc0400c30d700c1cc4c43f013c03040c00043dc00031010000030034000d7c00400f000d14c000100104c3c033403013034f05c014000f140037c0117c1cc40c0c01001c4d050001c104f0110134d10d00300d310c00043400c040340040040c510000030f3300c00d013033000c34dcc0400c4400c0c4f000017c7007ccc003000010035430030100003000040c0000003040c043000030440340000040000000c03110044c3f311c03cc0c340410431313005c0f00004000130000c010003c110c40130010030703000300000353c7334c044000073030c101010f400101f5c005314cc01d0000340f01f44400001f3cc051004000c010030d0000f01057dd03cf00c0040c400c77c0f043000030000c730c31f04304440100c4ccc300c03300303440340303c0fcc431000000dd00c000d1310103004f0cc0000010500d4470000c0010013cc130c00f003d30d40d00303c3104103037c007f03350100400010304c03110001c110400100d0003041454043500001031033000705f1c341010c4441040c033f03400c0c3c000df001703030c33c00c0c040004f1110430c3310f0f030c01130011111c0144300100c003ff0c0515030000fd000403150100c00037340114300d0400401d04007c0000043f370300300c050d00004c013cc30d3010c1c4000015330010f3f04010010400c033001cc4100c1100c04c0f100040cc17014c7f030c00000704c00f300003040004310100000300030c0004c501c400cc00103f401cd03d0300cf00f0c03010410100fc07003c3330100f3f70d4001f037ff304340000403330070c001d00000d0c31001000c40000030000030f010c00701c0050c00f040c01d0100f10000c0c003000d0444100c0cd04c5440334040c35dd4d1c430c00c00141003f43450047000000c00f01c40000c1d7cc10003f340105cc070c310c000c0cff01070707310304043330c04000c40c0d01cc0430043c01400c070033040300cd301c00005404001011000c0c1130033f10c0c40c150000c1010400c0c047cd04005500011c00c40c13f000f03000011404050700431c000400300f30000d003fc03440313730f01c00303114000c0305101153000304030503033300fc031400ff00003300004c1ccc0403c1003101000000300f000ccf10f0001340041004000010111340004047000003330100140700110000301304151014000c00c10004400343000c0504304c33003c330d0c007f041f000c0c31330040000c37d004000010d30c;
rom_uints[860] = 8192'h11103010103100047003400fc40001c0d01300000cc00043f0d144003c00cc0000400400500334003003300000000001f4005310c000015c0030307c00000cc000031c00003040c00000435414100003030c4c1000011f00c70c0000d030c3000d00000700f4010c40c4030373003c700c00c1034c310c4c030003030430cf50cd000c000c00170000d0c01c0010000041040730c0304c000303010100004304041c0430c03401000300000c3d14030070044330030030d04c0001403d003101003f0300c0c300101c0d00c040c40003001fc00c0c443033f430047034000000c3030000c000f44403000fc034c340000000007c044000ccd040000d300c300000000110000001004000d100f4c0553101d0c001c7c410f0d03000001f0100cc00007000100703c7000d10c0010100d0100c0c04030000c010000cc340f7c0001104000dcc031c0c0c0c40530c400000d000cc3004d433c00c41004c3010c044c000000000303404c4101030734c10504007100100c3100040c011c44000031310f0c0011000005c000000f40000030000370001031c1c400130000c074104040c4000007d04014000c3c0101c00c4000051310100030040300304031000c4030c03cc03c0347100c003000c101000030c50c100004000340c003d000000051100003c1000cc0c004040004074c00313c0000c30c01c000cc000c0004010fc000c0310000c0434cf1f4010d31ccd0000035d000c0300d0d00054400333004000073003400010301703f4000c31740300cdc3300000c104c3003dcfc10c001001400400c030cc410c0c71310050340431c0f4c0313101000303000d5fc033c000004040000710c11c031000745000c3c000100430330130c003c0c1000400040f100047013c3c4cd410c330001c40f0000c300330f00000f33107c041cc40c00c00401071c0c035030c0000f00cc00100cc30010f4c30d3000300c0030010004000c00c0f1000140000404040d1010034c10034104100014c30fc004000103000c00c310040000c003c0441c44000011010c3033c0010003310110c430000100dc0400dc300300c0cc0c4015010c01c0d004f300000300030700310d700000004070dc34030d310c0f00f001c77c3c40c3f00fcc0c034103f3047000105114ff000c10c000400c00f03004000d1000003300d11303403000000c010400000050c000004045000c0c00030c0c100443030030d01711c0000511c01d0cc3001400c00c40400030000700001041007c0034500130003cd0400c3c000ff301403c0cc001003100000000400c0c000c11000c000530000030400004400c00004304d3055dc3410304d0c330000000035f300000000300003033400f31c0074330400400043df3004000c30000ccc0000cc00004040400fc100d744000040;
rom_uints[861] = 8192'hd00c300010c00c0c0030f000004c4001c300007c001300300c050000310c3c000000340c073d0030c01c04003500000001030f30100d05100000000147004404c41030ff0011c014000014300300c010d00300ccc3051c3003c03cc31040041400130101300c03000110030c00107f0100003c4000000c0f000700031c11300c04400100d10c3003000000f04500040430000c030000000103000003401c1031000c44c0100cf000300c01d3300000000440000000033503100000300c0300300000057030000103003000000c0000303d00050c0004c000001103334f3103403400000130711400f0cc003300c1010cc0030100d004000000000010cc000000c30c00400300310f1c01c004000001cc0003004403000030cc03300c03c0301f0003000010001000000700000c010100003330000000110003c05c00fd030033c4c0000c14010f304100001101c00314100404f00c000033dc13073c0c3c10c100c000004300c004041301000400001c00005cc0130100c00003f7130fc001000c030700c7000c300043300c00304330300005051000000000010c130c10101000d053c31404c00c00003030c401c100d04004031330030040033f004003c44c073c300003001070057000000700041303011000000400001001000104f40ff004c11301003401141014040d000300040c0003030c00c001c0030000d300130cc01003c0130300143001003c0104101d101700300c00c00014003400010cd301000f0c0c0030000f10c1300c01033300000000000d0ffc0c30c10100100c1314010043040c000f3000340400c043000000410300013310003fd000313504010c00030000400c13fd0001105c010103003f1000040c30c000000c05100444010003c0003004000cc70c110000c5000f130340331300131013000c0f1000030f0c7330040d00d40f04003c0cc400001000131c3c7303300340151734d000130001000005f100001000c034001100100300c0fc034401f00500d4000300c300441001000c400033101500d03000c00300000000c040300400103013c430300000101c0005c403c100430400c300f00f0035305040003401c70d0c1333010105000000730004c4d0033434c017100003cc140c11300400cc07130d0100c0003f03003c0c003430f4103000030c10113000000c00000400c10347040f0000707003300000034c0dc1001001300003f310c0033c00d30c00c0330047040c0740340000331430000010403000030030f00007030001003c3340c0300d001300c0dc00c03f0300003c54d0c30c000073c1c0304000300003000010110c33c400010c003c00007150c3c0030000133cc30c400400330311003001100400000c40043040340f000000301103500005c54000405300001030030000330411000f7c0f000003;
rom_uints[862] = 8192'h410cc01d101c4100007000c4300340330403c100440f001030050000c0c4434000040317c300007755c0c3470340c0d101400cc00333000003c0cc4044cd0303471cd30010030003000f7cc001c30c43040d031f400001003c0013100c00d400dff0070410340c010313030c00730d000100030c017404000d4103c03510dc0c10034040c0c0d104030c010c4000c5f14000000004c10300000004c0c100c01c474040c0000cd011c00c4000c1c004334d5000000ccc4473030c00c30d000c40cc1001f00043c37000004743c01f04c0cc0c0000440301005c00050031100000cf0c30ccc000c33c75ccf04441043cf54004cc40cc00c00f100100030000c4430cd30000301000040101df00444c031331010c0147f00040f00010075704004000740010410000c00100c30010c301d001040103040000c5c0010c3017dfd0c00301d00051c071c10f00033410c0004c70cfc3c3030fd10d0000403301000f400c111c0303010135100cd10040f10300310400cf00000400000010000311100340c37010c040050001000c005000cff300044040013010cc0f0f030040f00401c30d0f0c0000001000011100c1c3c1470030004300d00111ccccc0003330003ccc0304003003010033130044c1c001c0104305fc0d40003004500343340400d30000c040c005000043c105000044005c00c4f314c030403d000c401400d14330000300c3000407d373300403d003c0003301440003700004c0f4030dccc0740fc0cd01404400f0000040010700c0430100730000d4c3040450113000000140000404471470033017410fc0f34cc0000300c0004034d3c3c00c001dc1cd07430cf10f0035130043004330003000dc01040f7000f04454cd05005041c00300cc0d000003003000003c04fc404003044337c50c40100c0030004040004dc0000100c00cc000030401cc03c17001001045c041000c0304430513f0cc0700400040313003001100cc070334cc1700f003401f11000000000430130400c30401cc410c0000c031004c04004cc0303040cc000cd00c00cfd00300034007cc3d0443403401c13001000ccd3f00005400c4c303311330010300330001c0000d4000040104f10c00040300040c30300300c3010c00c0070047c3c0000001dcc003004707c54740cd0010470104c3dc1043c0c00000040401040d0144c1110cc00100333400100000000003f100c50f300000c004540cc001c0c1d3000000000000430170c001130d3040ccc4c0300f11454040c10111004fc000c4044373440004000015c0c0450404c4113300400c1304c0c30000f0c0004000400100443000c000030100c441d04310c307c30000100004c000010003010c004031c0030d1300300404407f030d3003404f34310f040007400c0c40ccccf1015c44c00014c000400100;
rom_uints[863] = 8192'hfc0c00300c110110341013500d0404c304033c0000300000c54c003c0000cf00001700305030400034041040003c3c00403314310010f01700d0004700347010403cf0300000c010001f10070c30c40430300044d400003010f0000cd40c000074d1c40134c030100070003c00d00000003cd40c33300d100300d3c430000051001000d03c3000005000300000045f00300000000c0d143cc0c400c0407cc03330000040000340f0000040041f0c011050c03000001000541c00004004000c10c004101014010007cc04140c0c343c000400041000100300701000000030c50054c004c0544000140c00000c100014100c000c30000000003000000030103105003050500c134c31fc1cc00300000c003410d57c00f10043040000101c3430004000000004000003303434400c00340104004104301030000c4040c4c3000c00341004100030d0f0d4340c000c001004d40000043c5030300030004c04c0c4000c00100010113c00340c0044003030000c103c0c3010001c1c404ccc000c0430104404043030c0c00034000310c0000c0000000000003000f0003004401044cc140013c004301000000000000300300c00303c0c7000004cd0000004000030d0113040400000f0c40000303400c0300d0010301c00053c44700000404030740c000cd000131300000010343c00300f34c000d43c1000c0c300000070003f331400041334000010000cd5001c030040001c400030103000c013140434003010543c04d0c00400010030070c3100d0c0105010003054f000107070301000140f0070c330001c00cd004c503000343000000c00c0c0004133310454d0c0d41c0c30170430c00000003010c400443030c40c10f13c07001f0004003c044c05003c500410010000c000004000c410d0007000300050f0001000003c0034c000c40004041000cc1000040c303350043c303f0c00003c00000070001401330c000003301000304000c00c30000040c0303030c000303004135010c0c10c700301c030300014103504c040003c3000000c104031334f7000004000030cf030040c1c003d404c0c34c0000c300c100400000014c01c00003c30000040001c0313003000c014000c40143c00003d1010003c00001413305c3400000000700030001000003000c0300030703000c0cc4015c00c3c00003004340c0c401004000035c04400d00c400035000000d4041000100040cc7c00300c0400070cd0430c1400300110fc44f330001000004000103c70007400001370c00000343c40004c00040000100017d0000c003000010c001000003040000110000c00fc00c4000c000031000400d0d070047cc03413103c4c30d000000040030dd0000440000010d0400c373c40000000f5100007040014000c01043034001004403030c400000004003c0c00;
rom_uints[864] = 8192'hc000c131704111033300444070c001f0d00000c1c7c00000f003c300d300333040c3304f000003c040034103c3cf0031d0cc050cf0cd34000003013005001301c0405c000cc0004000c400c0303cc1003500c0c13c03c0037f044103d3000000c10000dc00f31103cf3003dff40043307430dfcf000130040073cc0140410034dc30314c00000004130000f01135c0c330400000030401040300043d000f10ccf0033000cc005c034001cfc00030403c1030000fc05130c0000c0c0030c300f0304440000440030303003030c310c00330000111040c03c04007313000001003000000033000c0f0f000f11c00c00dc300c44000c000000001030000430033cf3441510170c030330410c0f0034333f1d0544f03f0f01110c030d100c0c0f0c1000000001c100130000100400c00033310c4c301110000040000d0c0c3330100d0001044c11030370003c401017000f00000030f1003004143fdc300004000c0c0c0c00c13103c3c0c7071001301303330000043f100c43fc00000cf30300f000370c0d03300c0404300c4400034304000f0f00000000030ff0300103013010070304441d0010400f0d000f031c005003041030300cc300103c40cc04700041003f0400c00001447d3000000003000000041d031044030000053433430003f0001105f00c440f0074100304ccdc00333dc04340400c1c0f3c700cd10d130c03007013000f1101400f00c50403c003031340f1c0400f0040f003470305c0034300c000cd1510f0000f3c133730010050051001000cc0cc3001000f1000dc130c140000013300030c110d1c0c13c0040c000300014c000001014150014fc000f33000415333ccc0300470cc000030400dc330001c4411030110f3010f34047100100c044400f0000c010000c300d0c07000001d103fdc3000f13100001c003730300030103cc41c0033310f40000c0301030300cc0f0c0c1003003d000f0000d0044c300000010c00400c0010000c040c0430003c43c011013f0d300cc13000040000003c00000c4000031c031c00113d000100300030c004030700043055001c001400000000034000c30040033c774c13300300040c10003370131004001010100000111413003c13c000000004400d30c034030d34010010d003333c44711cf101330007033500c1104c10310f03700f3014031d031c001d0300f0010d0c3130003410000000300710000f00301001c3c010003413030300003010701303c00034300c00000d30303f10c40ccc0f0c1100c0000000000434104000003050fc3c11300000cf3030033001037400070044000013000d10040c13000000cc0d0004030030c33cd1010c0d11010000103410d31c010100043001100000c00c0033303000f0300f401310040330070d003103043000c00c0330331c3c0f031000;
rom_uints[865] = 8192'h5001100040004c00cf00140c1c4040000c003000400c10000c4303001301000000c004d34343400000f0001004000c030400c0c40000030dc0400000c30000000c0073300000014c4000000404001c000c000140300000c0c30053300005000000c0401c00c00700c0c003000400f00404000014030f00c400c0000c30000000f30010c00000000c000c000000000000c0000000001040001fc1140000000c00cc10000000fc00300100400c0000004cc0000c000030000000c0c0004003c0c000c3000cc004400040c000054000030005000c01c0c00000030374c0fc010440c40430000033000004400045300dc430010003c000100041040c0010dc000000410c0c00c000c0c13d00000c30040000070c005000003500cc0400c00400013c000010000fc00100000000000404014000c004c0000c40000c004007000100c003400000c003400000f0013403000100335c10034100c0cfcf00c4cd0004000400c004000010010300100c00400000000c30300cc337100c00001c004700030040400054c700300000000c053000f00040000050000000000000003004d0c0070c4000c000300041000000c30000000000000c04000000c000050c0000c4030014c1003c1f000000000140001c300000400140000300005dc0c3000300000c3104000c4100000030001fc04000c0000c000000040000041c0c0c0000c0000c0000000100000c00430c000051000400304c003000101c003050c3030033010c0040004000000c00000000d0000304000005001100100040300000f000100004c000c00c0000c010000000147030000c00104c0000050340000c000441000044001003004030c0c3140f405d0c3000000c000f0c000130100000010000c34403d00000c0440000000000001c000034cd00340fc100001001c0000c070400000500c7c40303004c003050000004400cc000c4c100d003000400440010400030001005004403c000000000040010c040cc10000c00400001c00000c00003304103403000030001000004000030c031000030400f00f000310000c00c0000140fc40000cc0014010010c00000003000c00041c503003000000c0c37000700d0c000400d340000450000000000d304000173400040404000c00000cc300c01070041043c0401c70cc01c00044100304440cc0000c0014150040030040c040404001000c00003c700000000000000000400000c40000f0003030c0030c0000010000400cc000000c3000410c7150000040044300000000310440000c000130000000000700c0c044010301c00c00400001f0000004c4c00f000704000000000c0030f0c0040000014c0000cccd030c00000000030c30031000000010c00c40300001000c0400001030000000000c5000040cf0c44000300030c0000c700330400000000;
rom_uints[866] = 8192'h3070000040000c3c3c000ffcd04c000040c0cc00d0c400000004c400c0d010400044c050f01043100c001c00000cc1010c04f00000030300c0c010010000c030c000003000c000001000cc54c00014370000c00000f03004df00f0d00100700000c010cc00c000100000c0c00001c07c304000300c0cc0003d400c30003000001310440030300010300004c44c4000c000300400005000dc3010504050000000100030100000701c00100004450400007034f00000401c4c000000c0004040000404f0f030101000003000000140c4c01007dcc00401100c003c70c0047000f00110004343c0301c00c0401c003031300030400000004000400c0cf4403013440040c0f00c1c000000400c30f0f000000010c0004000300f3cc0035cc41cc0c0010000000000fd40000010d0c00004c400c44000100c00000000401cd00000c0340c0c004030400004c1003c1470405410f010000004400030004000c0c040c00441000c00003050c0304030000010c0003cd40300000cf004305c000004c0c0dc40d074300000407010010000f040435000001010007400c4400401c00000cc43c040fc04c000000c00c0007040c034040c000000104040c01400004040c0fc4c00ff0c100010c0c1100000400c50f070501300010007503010c0003010100000300c740c00c004f0d400000c00000c00000c30c010007c50c0cc04cdd03437000404f0c0000000000c001040000031c700c03030104010d070f0000000000011cf53040c1004c00040003000000cc0000030c000101c0000100000f0003430007030ccc4400000100470044410d0503010c0c0100000c04000c1004010100000f000ccc03030000050cc04000000100400c03030013000300000304030104001dc4000c0c0c0000c00d040400370301054403004104cc00010040fc00010d0000000c00300013000441c711043c01030c0000000d000c0d0300400000000c0000010100000000400300000c0007000001c00001030305440340000300400cc3007000510c4c000000c1c3000300430100030d000c400003000000030dc00300000501310101010c00c4050c0f000c4d4703000500040001430c0c01030c4104000000000f4f0000004f43000101000c04001d000000040c13cf01000c1c00c0ccc00030c0400d010d4c0001000700000c00100c040010c70c00000c014101d4000003400301c301000004000000000f03400040030003034440c003404440c7c0043101003000410000c1030000355001034100030d000303d330000c001004c00c00c14343040107c50700cc0c0100cc00c1300000c300c00000cc0d0700000500c00c040c3f00c304000100000f0000010000c0010cc401033cd700000400c40000100000000014c34d00001f0041000403c00771030104000140004400;
rom_uints[867] = 8192'hcc050000000400110077c7400f10000cc4010013000c0cc000540100c4005000004c040743440000c0500c00cc0cc154170dc0040c07030000000c01c000033003040340000000040300100d000000cc3c0c0000d30004000005000000004000c3c3c000c3000041cc4335c000c00f00f1cc30c0010c035cc004030311f04003c1300f0040000070000300410d00000030000000000000000f03000c03cd7001c0c0c000c00f0007400110000cc10f3000000000000043000fc000c0c40101000f0c0f300300c3031307000400030400400030000c3cccc000f10c300c03c1c0c0c4030c010001040003c07d00d001c34d40150400400000c3040400c00000410c4000c0fcc00744014404cc00100c040100031cc0c4100300c10040000003cc0001c3000c031c0dc0050c0fc4000401140d03303003500c0d00c0004500c00000c00007d1003cc04503140f4700400000070140c301037101410dc0040c01c0000c040005c000004d30440c040000000401410000000330000440010000000304000c10004cc010c00f000c3003010c0400000c4504cc43c04011c0c000400401034000010300c0000044000000000000400c0d0d0c00010000c00f010c1dc000c0c4004c430003cc03140000000140003040014300d01000c00000c001001300430f1400c0cd010c0511c0743400040d0401010c0c1000400f000000cfc0c4100030000d00c00f134117d000000140cc0f0c100403c504cf3047c700000000c3c3400300c1000c01003d04030c0c010034cc000004cfc000c0000c000001000105c03044005040c004f003330fc0400000c0c304c30000000103d00c0004fc30c0c0c0370400d3c4c3c3404fc101000300d0410f00f0c0c300000cc040c7000050c100040c00000d310c00000cc10041310f04014c01c100433c30000000c011c1000003400c01cc5040100f0f10010cf14400000c000c0000447003c00000c1c0010000000c00c4c30c400000010fc005000531c4fc0300100400011117000000c30003cd101500004513c73040c3d3cccf30c0c30000c300010c4000000010044001400400010c4040040c040047040043410000000c000df30173c40041033c0003dc440503100400c00000401000c13d144000c00007d40140c0003400100f0440c0d00cc0040dccc0c00000010300440c00c03400010430000013c3400d03050d0000000007444040000004c0d40041040c1010ccc0c000040000c300030c700137000000070004000144040000cc40c3000c000433300c03000004c4c0c1c1cc3350400c41d1001f011c13c3000000f0c0000c1000334f0001404340cc11c00c0303c303cccc030740c400cc40030000004000fc4070cc07cc0000400f004440041c0003c0110000c30c05030f00c00c41010c105403000c000c0000;
rom_uints[868] = 8192'h1004000000000c5000403c404cc01344fc10001700c10c4130c40400551d070c00cc000c3040000c4100000c1c000c0007111000150000110000cc001d003300000000001000533000000c103000000003d0330000100031cf4c10700003c00000330c10100041033107c400300c5c000000000530c33410100d34730c4cf100000c1c00000100f000310000d000000cf00c000c0000130f10c04304330734344c0000000000fc10c00000000040300000cc000000c33c0c10000f0d0c00004000d0010c0c004d001040000010000c031010330400410403000004001d010003403c0000c00c000c0c0100d0414f05351110013041f300040100c04004d10000000c7140003c400304c30000f0003000500000c10303d3040000000300070c10001070000001d00c00000c0003400001000100045051f400c40000003010c0403003001001301000d54010303300510033010010c00001d101d00cc30340c430000040c0100010103000011101001014000300003000c010000dc001003503401c00055331000004cccc0033700c30005c00000005001f0c0f0c3011010c04440c3c0101004300070030000010cc00300000c00104d00005033004f0000c01004007010034c140000ccc130000c0c33c030105013c000500400f40001000000f00004000003000c1c0000c001154040cc10013c4005370001c3c30431104000c1c1001400004d0050105000033010d3013f031104130030011004170341037041c000c00001010d001c055100100030001305710001000030053001c1f00dd31c00100441000c300003f53010030031304c010303f1000051510410cd43003100001004f11400500003000300110040c57000340c34170000f0cc004c501700f41f0f40031041040c70003014c1030410107d050110000070010110031cf100cc05001cc00030150d010fcc100100000100000c0000c001140301300c00c00431c0c34300000110040c10034034000700000140c003f1400c0040c00044c00007000400000c0000040001447003c0100c000034003300010000304013030300000330000300c30f00300030040400070c00000013f01c300300101300300140d0c3400000135f004d700d00010f3000003cc15f330331043075000c040c03014555000000030c0451300c00c0000cc003000000c1050300d00d11000001310d3f00033000070113c1000d00030030300401c000000c0000030000000d1410000134043003300c31400003c3004101c0c010010c00000c1005000510031410350d40000544005c000f003c005000404f50001040c0c0010411010c100000054000000001030f1304c40043300000c04140d100110010c003c4cc0d00040000000000f0000c3003431c01000000000410cf030000c00050400010c00c010000000;
rom_uints[869] = 8192'hc010040031c044013100030000001004030dc010401f310100ccc1001001100430013003013c000051440000c0307340c0cc4000d100d10cc010004c00040000300001c0003010000300054100001100300000044011000330010030400010f000000043000030003010c0000004000330000300300c305c0031d004111c4c00c01047f0044003c50007004370100100100000dc003300c071f451c0d030007cc350f0004170300004100000040013c3111d0300000300140030003c51c14000030030030000f1000000010334f0c3100034f3cc0001c03033000000f04f000d0000c0c00310f110101c300d0433000c30c00350000300003003c0cc401000037c34000df00100000c0f35c00310000331301001711f3000000110530001c0300030cc00000c00140000c103000c0000304c0001c000410010100c0107c0f030100343f040000300d0340c310c001c00300001d40030000f41100010c3d0703100c0100153c00cc3c0c000d0cc300c011403c0c0c04f40010010c00000000d005c34400001fc101c0c300041000000705300004000003700fd000530c0003100133400c00070401f00331100300000010dc000000c03103300c043c1030000c31dc0000030000010300003005001d303031001000430d03300300400d3300f400010f011c0033c00c04c31000300d00cc410300000013340104c3400c04000c0c0003300c1010cd00300cc4001c0f00000c00c0000000300010cd3401000cf00333400001303334000f0000c03103004c0d45000001030030000d0003c0013010f0074c00000404010031d00c0000710004400000cd330c1101c313070301003340000d0d50001040040f3013300310003014000403d4300c00030101c00100000c0c07101000010c0c0c004040010404000403d400303000000000001c010c04c0d040c00c0400c13103003301034130030c050014010414100c1c0030000f00c001010000000003000c000044003c430001c103000cc500100c000007c100033001000c01000030000c0d1c330000001000440c3f3000000131304410c30303000410077030413000010000031030053100cf000000000001d000040440030c0c000d4c03c00d0113000c040300101303003f30f750000030c403400c330511000000000410c300d4303f1014417d330cf0003057d00ccc01c40110c10df0770001430000000043013401300c0c0c3d00033c0c0f04010000c000403c0d304301044000000031373cf30100c10003030001cf7403131003010001c0000c0f100100cccc304cc040030c034cc50c00c000fc1010f00f0010004100050000000001007d00013c000000034100000c00c3000000300004033003c1000000ccc100007000003000004c04000c00303c104300100400043700001c0c03003300000;
rom_uints[870] = 8192'h40c400014c700000c3354000401044cf0004010044f34c00000d4f1014310700050c14140c0100040003c4000401004000300013cc30304730000f043010c00003c44c3c0c0d00700400003003004f0440c331003440405005044c1500c010c11733c0dc1c330c105444c30004440d04030f401000cc103000010050000151041000f34c0043004010000004cf00003c030c3004000c14fd30100000043f0d0337f00f000c077f00f00400c3003d001d4f03d33400011434041004403710041411c7330c03053c3c00c01400040447d0140010000c0350435d0410c0000f0000043104000010003444c44005c0370330cc0c1445000000007000c30c0400000071044000005cd401475017430f7010f0c05c104c30443010304004044c3c33fc0043000004000040ccc4d0d3051474c0000ffcfc043f01000c01043ccdf3cc401c33000c43043050430304731c034c040343000005ccc3000000cc04044000f00000000cc1001340cc044400004100c0000100304d004d044434c00c014044003405444d374c041cc300000c44430c300103d0000000d0c4340040053c000004c7740f104003003000cc070004040f40704c0c0403c73001cc01501c0030000c0f00c00f0404040400fd00001fd0040cc0001130000300441c0f1f00330cc5300007c0c31014cf00c4415c10c107c0f00304740030530004347000040004c0300c4000743c071dd013dd03014000c04c4300cc30034034414c040344d44030c17c30001403050343001c43c007010d033034c0001444c330c0c30030043074031f030000440c7010c30c03c0000c3c000000004c01044030000c00000f4c00040003000ccd4c000444004030000044d03500400c003100300c000c0c004110f1000cc05100c300c4cc7d00145000347c34cc41400300000400001f0040004074cfc4040030713f00d504fc0c370300331140f0c03050c473400131301c710014300c1c5d3c00000f040f00c304c0040f17dc710530040f3700033135403001010c003300140040c0000034f3400004001c143053034d100007007304143000013c07500c0d7053c05fcc00300001c30054040300004007400003000c33000000400010c00c430cc34301cc00003c0500043dd41c0100001cdc0d000010d00100300c0c50001404f0003000030c15040000fc00c00007304c04030000cf1f40044c0000cf00700070d30004c0cf04c130f14434300c1d741000000010cc07434000101c3f14140000070034070dc1301041101c04030c0fc00414cc140f0015000f37cf3373000030cc10104f00404f1f004500303300c40c0004c00014c103004305070d004003cc43300033f00c013f000c0c00001500d040dc0ccd13cc00010c04c104000304c13c104004300c03100f00144403130c4d54310fc43cc0003c;
rom_uints[871] = 8192'h1140000034c17030030500c1dd70000cc00001703700c0cf0031330300c043c0c000003c30400140030c10000f0f0030c1333c5033040430c040cc10c33000c1c5011010c04000304c00004c40001504007000030003007c700f310f0d4000000c05034c0000cc00c00c101c001c1000f0c7334300701c3c00f100113f00c0005f10100c000f304d00c00040f3100d0d0c0f700000f4c01dfc0030343cc0f14401040000045440154003000000dc00000003000c00000ddccf0030c3dc4040101003c001cc40005000030000dc1000004410cc1140f01f30c0fcd0703cf034340c150000155cdd0c0003c00110c13734ccc1374103c0c0d10331053733010030f03cf5c0300c0074004010050f003c0003c030400400c17030040040cd11c0000430c00030f070010c101430100cc7003033c3c3700c0c000410031043d00c0030004d11f303f730400040000c40003f0430c100351501003f30577fc0103c1000437170dcc0170013340c1dc5dc0f03301000f00c4fc0001cf33030c3000f0130400007337cc000c1710c010cc404171c000c0c04000c000c00001c00040c0030034034d0c0cc0c0cc00037004c4330c1004c300c4037c1001070dc0d370f004305000014cf1c30131415014400400031400df4fc0c1377007cc0031103c1cc010001741c0dd0030f003030000001c010700f0c1c00c0f043030c00300030f1044000f0d300c00000004411007000c0000310300f10013000000dcccf34c10c1c000000001c033f0070cc3c30001c000001010043340c04140110100000c0cc0f0301d110034f001cf5c00c03cc00c4cc4d0d505570140c30c400004003104c0cc300041000c3d3703131003ccc131070dc040041c4cd3404010c0034c000c00c71104cc00c0c10c3c0c00c014c0037330300c0110f01000000c307d400443034c3003300001fcfc047100c4000000cc0d005000133030c0cc0ccc30000100c740041000000f043fcc503c0f0dcc3300014f00100407c01c000c0c0c03440cd1000005c70f000341401000001c00c005500005001c10030f43033003c10cf00f731c141cc0c7c0f03000c00000fd00543c00040d1f003000004300000300040c110000000d000454001010c4001c0005c10cf4500ccc004c3c510000c134c307433300c0300350031000cc00000d00400c001d00c00f0c00434031001454740403000c00030001c333000100700c5c03400030100c01040f0000000f03c34d000074437430004c03000004130000454dc0030fcc077c100d000fc0cc7cc0cc0f41103003cc0370f17005443d000000f00d0110034000c0300103c0004400fc0f0100330c037c0c70000f10101f010000000477010404c430c0c010030f30000400001c0c10c00c30040c0003000c3c00d0000030f007300c3300011330c0100;
rom_uints[872] = 8192'h43000070031000000001c3301c00030000c311014f000000030000404000000040300001c0000003000030f30cc0d0433130013000c0000030401133401003c030330000000001000c010c000003531001001010010f3300dd703005100301015111130000030300000000031100d3030f71100110003000300000c0110000f03040c0010300300300104100010700103033000330141000331300c00c0010300030000c4000501110000000300010010f10300000110000100d17000000000300003000d343400300000c00030f33100301003fc37330c1011103f31003010430033001c310000113003040000100005300f30000000000000000110003030030c00cf7c1c003710500010000000013001101010040033300c03330730010f134000000030030000041300000004c413031310300000000000101d1fd04c000000040f005c0010031031010330000005304111000011301010000c0733010300031c003001001000000031000d10010000040304100010300c0701000300c0101300300300030f000107000033033d001c000030100010f0000444000d000f01c001d0353000000c000000010010030310300310030100133d003c0c0d001000300100300c300003040010000300dc0100000003373f004100000c0c007110300700000140c1001350310c11000030010051031c010000033c003010300301041c0000103010000c0030005d33010004400001000033300c0003c000001100033d100051010000000d0110100c113c1410001033010314c07033010001331000001014001100005300c40003300c05311c0333040c1000f30010100c051c3d0c103713331001030030033301007c3130100130004c030113c104000130330004100110000c14003000013d001d000000000000330010003c000011003100104414000030301cccc004c1400c000000010000100030300f101c3100000c0000000c0030000030030c001000100c3000330370d500000307040003303070400d000003000030f000400d340400010317303300003000010c03030051430c033003000330c03007000010000c3c150c3d0301000030100110d003000f00000330100000303d03040001c0100003030000010103037c4000c530000000141f11330011000000030053100c4334010001000700041111034304140501003030000f3000300f00004d1d1110003c007d0040050c030310430c30030010010c000033003d3000100304310000031014f070000400311000510000001100103c100000503305030034000000000f00300301305f000c3f0334010110000001001105000101f014f3c731001300033000100433003001140000001000400110313000301d0d0f31c01c300004111000cc300007000f001100f00000000c1c07000103;
rom_uints[873] = 8192'h10040000000353df4771070f0010041131004100000c010040054004170000c00134010c03000c00cc0100110c0c1004410c0f0f00000dc100000d4000c4401c0300404300000f100001000f000c003c10040fc374004140000000400c0dc404014100140c100400003013404314004340040350c00004100030130004004034fc00000c03000d30330005000c0004f1373c04000000000010c0000040030000430010c0041c100c4000c00c40f00c0c04c5500001000f3100000f00000c0000f0d040000007000c05000400c00543010f050c0104000000140310d00040030cc0c000000000cc0040d44c330f430404040c0071100f0000030000001cc003350cc0140d0c1443030c410c4c0c0000034034000011c007000c0000430c4000100c30000d01000c0001000300c001c50100c000000c1c0301000001450031000000c1040d104c100003000c0010010003001003c500304d1000c3043d0000340000f100031070100f00000431003503400c004fd0101c3300003031404570030dc004701030c00000d0054101034307000003000001000404c44c7014000005440403000c4001010004010000ccdf03303040030040cc0530103141000007f0000004001c41000000d701400c400030c0430f010400cd0c00000000030c30000c030c0f0d04000031130d0000c51c00400100000f440003030f00030010c10c4d040304030030000013c010cc0100000001000000030000f000113c74040401030c00c10c1345f1f000034400000410000c43c0001d03505c015c0c0310440300100c04000000304070c311000040c00001000001c0100000400000710000331034c34300034107c4c3000000c0000000d13d00000c5001011000000143030c4101cc040040000001030c0404000f1f4c00000407030d0301c007d0030c0d0c0c00104300033350c040040c0c311100340003700000074c050c43030105300030c0000001000001040000c0000000030000c01007400c13003040040c00c50000d00000010c1034c000c00014c100c101014000c00000000070c0000500001001c030c00cc0000dc000010c4403000305313000000d010000000c40c304030d0c00400000c000c014c10c3c0c1c0000001000c0f00370401700c04d0104dc001004040100100004100300c30000053100015c7000054000c00100304c000040cc000001030300010000010404000410001010d003300000005140000c03700000410741050000c045300d0c000001010035000001400730434c0004c7400300010000d3000c11cfc00000044000400000031014004001d000041cc0000040000c0440110011d170104c0303000710030004500000001014000c004c5c010440dd54003401303000340530400000001000700c0300c00003c730dc4c70c001000;
rom_uints[874] = 8192'h430000410c4400c1030c00c00c70043f04f0c000c00404003c01000300c7400010d003007000c000d0000400c004000000c4054c00000000000c0005000c0010001d040c01000000004303cc000003c03fc40cdf30c0c3c01103c03031cc00000100030000c1000017010001c135040c00f0c54003c4c40041143c01030f00c55d3004040000f000030050c1003cc104000004004c004cd0000000c041c340004f0d03000001000cc000407fc500400100440000001000c001001000c00000730d1c0300c0000000cc0000cf40cf0c037040300c05c0fc0100013c004400010344001040c0004cc0c3004044c54511d51403300c0f000004030c400000000300400c000001000040403140030c000040130f0001f00300c04c1470d544000c000000000cd305001310103003000c0400413c54c1c0c3cc4000dcc00100300000000004c0004000c001c3000c000010011300d1030300c0cd004300300ffc00310000c4cc03400001c54300010043030c010c7030100400030c0300c40400000003d0100043cccf0c00000000000003100000cc000c10d0c0fcf0c0d003000040070001110300c000010001f0014000c3c0040000030014030c00c0c544c1010070000c00c004c01110410000000f0100ccc000c10cc30f31310000c10d13003000000000c3110c0ccc0c0710c4000c434041000004c00f0f04000c01d1100c35000005f10cf003000003400d0110c01001c1c10400cc0ddcc4c0f3c40017004c010000000c00c700000404004c3c00000c14003c30000500d0000003000111cd450c10000100040000c0c330c4004030f700c1c0cc000000000430030004c704c1003cd040c003000310431400000d3f01340003f0c05040c00c0150140000c000300c0c1000141000c13c14f04000001c04c1300c30d00000c501110d0500451117c0301315c00c0c004cc7000000000140010300c00400403c70c03003300c000000c1001c000f1000000000004000400c004433000f0c04000d300000c0040007000c0ccd0d003004f0c0c1cff170c0c07c031100030fc0dc000cd0000c430400401030400c4c0004cd00d41000300c303d000007c00001110c0000044c300000000015c007c04c1004c030cf000c51c33dc30c000c143c404030f04710000303cc0c010c0101000c0d004fd33c0c0c101d040001c5c0000401c00300c0403c000030c0004100cf040040000100300d010000c004170013000100044004cf044000c4001040040000dc00c0000c00d0000304310c3030c011cc10d4000c00070000c304054300000000100004c500c10c030f03000000000000401001040c3c500c000007051300c0f00f10110100150c04000c0001c073440000cc0030040f015003f003c0400d050fc140c00c4f03000c15000100030004d000000000;
rom_uints[875] = 8192'h3103000034400303334011c0030ccc0070c001c3030304000001c00145c00340004011c4001301000f0300c1140003c070000000330300c0345004130c300000c410050330100077d000000000000c00c303100301410c504500411c10c040000330c000003000103140300001c0103001000000c0c0010c00400cf343415000150c1000434300340003104140034c00440d000000010d01735100001f0c00c404030500130000c01040c000330100c000030040000100cc0001000dc35300010000003500100401010000030c07030000100100010014000040c100f30300010001000c13101000014000130d0340405304000340400000004044c003400030133003d03001033000500130034c0c0703d0054131c03400331000000cc031000033c000034040000040007110004100000000300f330c400c003003407d00c000c03070000d3000430010301c404000c407000103c4407410030001073030d0010040405dc403440000c0010001000c030043400501300000050000c0004030dc03c000400f00103033003000330f100700d1000001410000f1cd010d00c10000c300c070cc01c3430104000140000d03000003004040444003d40001f01df104c0c140d0001041001300011300c00c370c030341001c00c403300130073171f0003003311cc00330100140004301010103030000c40074c0c30000433330300c004003c003c00f045010d04040001051000c000440030140007034c0440104c0c11c30105d001c00000f47c001000000030d010301c0c0031101c3300451004003f0001045000000334071103c01000000c10010f0c001c730c0434d00df030c303104430040dc01c04003013000010c0100c40303c0c0c00000003345d4000100c0100000000c00ccc1cc0c00c3005043f00004c0001400004040c130d004500c000fc00000130000304003000000c4d43c30001c013000014003010100c510001010f000c000c344000100330030040000004400500f43000040c0c0401d13000000c100010003d0033000cc003100c1030504000411cf0003c0c101004040000c404f000047530003301010010050c0004000050400141000000c00007303000000cc01433300030100003001c1000c1d11443400043003c04f0001d1dc3cc00315d0010400051300000310333111340c1d0c740003004710004030011003c7430000f00030001000530300c000c0413070310d4300314c00034340314404cff4410000c0f31001000310000000000103cd70f7000031400d00cf0010300d03c700000040330000017001100145070c00d070004100034001000100004000d30130017300c0c0003340310001400007c0030040030d040400c01030f4010301000140000101f04010c0000000000300c0c0004051401c03000001000000;
rom_uints[876] = 8192'h3030f000000c40c0c0041100010c000010010141c00c0000340c00d300110004030cd0000051c000c040011c400c40044d0001c00543cd00000000004000c00004014005004c000000033c00000cfc400300000d00c4303000d47dc00f00500307f40300f4000d0ccc03000c0030d00c040003c300000000004500c050014000c0070000d00000000df0c01300c00031000c00000000503140104001130043410037330c300303104cd000f00c000d40c7d0c0000f004000c3c000c3c01004001440c004c000c10030c00000c0c00c0c0030c0cc05c3d0c41440c101c04003c000c00000c05000400404004fd00030000c343fcd100c001400000c0400030c70c300c000300010374010d3400004074003030343400300041c300001f000c00000c00000011c00504011000c1010cf01004000f0400c000c400000030104700444301c00050030035c004430100c300300c0334000100c4c410730cf10040000d000003050c0130040304d0000001000030010370300003c104c0c700000003c033c00000040410700000c0401100400400d040c100c0011c1ccd5c005dc10040cc1001100cc401000010000c4c3dc000050000005000033330cc000000cd00c00000301c50013000010000c100c04c00000000001d0d101c0c0d000dc300f7300000430f0100000004c401140f000000000000c4c141140c000d00c03133000d0c014c000cc40d00053c00301113400c15000c00004c050d3430307100f4103c0c410f00d100d00040147300110001000033cc0100c300000400000f0070000010001010300100c0f440100010030340001c00700cc000000010c004000040c30f10003400000c00400044100cc0400000c001000410c34030440c13000c0010000c00c010c00d100044000300d3030405c7005400003000000c003dd00000073f100401c000000047000000410407cc011700c0d00c0f0140c010c0c10000001011001000000301c00c0c000000400c0400400300741c010000000c0044040100000cc151c0470c101433300d044f30003cc10cc000001040040c10003f00400007c00d010145c100004400000040d10040410000004034f00000000340c0541400c000c0040c00400f0c0030000010c704c4540000000c0c30cd01000070c040001100cc0005003000ff40c001040140d40000400000c4c30000010000c0000404c50d0c00c00c00c0000300400c440000040404000cc3c3000104004430030c40043000f00040003005001070370ccc000c00330100cc070040c1000003003cc0010050c13c0c0000c01c0c0000000004040700001c00000000c04c004000004c44414713511c0c40001470000000031c4001007001c3c4cf00010410400040055034443c35134c3c0401c34001040400000404dc30c44000c0034004fc;
rom_uints[877] = 8192'h11000000c01000000c03c300100ccc43c00401000001300004007431c0c000000c370c000cc000000c5700300300100c74c043c0f0000010010c00330040004c0000c000010000100003037013c1300004000000307000c70000000010c40000000004d04c0400500c3700030c1404000f400410010340100cfc300010003000f7f0400c10d3010403400c00003045c1cf31000000000300d0c005000114430c004000001043dcc0003001c004c0000000c431000000404044000c0004400000040303000003070000c00000c003c3030004400c0051000ccc1400000300f0c003c00c33c3c00cc000340df005100001040003c443c00307033c0070c000004fc0430c0411040d00043110c14c0c4000ff403030d431c00401400d0c1c0330c701100000cc311004000300c3c00000003c0074c330701000400000cc40003700400101000044100c04000150340cc00f40c0040ff403c0003dc3f14003300cc000000c3cc04010340000050030003340001c0d14c30c10c405c03131c00010000d0c037c003003c00000733700000004d0004000000400c0c1c004c0000d130c4c00440000000040000c34c000050d0110001400c0c4014f0000300017c044c03c3100144c700073df00c00410000c04c000100030c000c010004034c0040c1000c103040c00030403141040001000cd4300cc101003034d30040f004400004dc003f345340431004c0f03cc400040404070000040031c0433140c0000c0010034c000000301004401000c53403d004003c0100003c00000c4cc0001d000c0400110000c0040140137d3c107003c13010050d0c004c300000000c0000000004d04000300030403c04c4c000040040c010403407c403413c0710c400573030f00cc355013000000c00140030c000c5000130c00400101c0100f4400033001000cc3c0cc7c00301103000300073001405403000000000c4401000c005d40030340d0001071c00004030300000000400c40c40c0c0073cc13cc4000d4f011d73300000000033105030000c00100000001003003000c0037c0030130030f3f4c100010c0070d100040f00001400300000307310c043f4d0001000010c00040411014f0f0040c000040f040041000d150000c00d004300f00c00543000d1301c4034003100300c010100c431403c003034400000c430c400004d030c000000030c0c00c00001c040000c40700001040030403f110d1c03300300000400331173000c0700c140f00004003c30c00c340c30400c03003000c70000340c000c04040003c0004c0404141401351000000000435700fc0d34f001c0041c3050000400040000000004c400c70c0c05300c00c0400c0c0010110c00010000001c0c0c03000000000430030434400450003040d400c03c143034051040f0c40000c000000000;
rom_uints[878] = 8192'hff3000000c03f0044f00300c340cc000c0510400c0300000010c00040d150cc30000140cc5340004010100d0000004003c5403001c010cd007c030003c0014004001000000000c0c3c000ff0003133140c0004c0030f000414cc0c0c00000c0000400d3cc10340c5140c0000000c3c00010000400c41113c101000000c0000000f500c003c000014400000f04350c0000000000000c0000d013c0c003c0000d004c510007017401400100040000000300f44300400c3040c1000000034000c303dc0004000004d0404340c01c00544000000c03700030d00000040003c0f0011005c00000f00000c003c00cdc0040f130d000404d44000011000041400000000c1100d04004c07031003c4040000073c0001040000003044130c0033013d474410001000f01401000cc40c0001040c0134000c3000050300000044700703cc0040001040000013003000440c0c0400001040000d0054004105d01000003040cc1005c40c0c0003000c4130c0401cc300000c010c40000000300000700404c700c4003014000c0c040c3500000000000c0c0000000504030400000000000000000030040000000101000370c44c0030cd003000003300004c00301011011300f0c13c40401100c010103d40000500cc34c000304000000d310033c4037cc004433000040300c3430c0004300c330000000030cd00010c0000000010005404000f0c0040035c00400000cc3c070003000fd003400400c0f03c1d000c343371300000c40404000f0c30000000000300c000c00c030c0c0500000003040140004000300c30000400003001440cc30c01000c013d04433444100054d004f110c4f40c3114c0147f100c0c00000d0c03000053c00cfc1c001f030000c303044d00400c000000c00003040d0c0010000fc00310310503040000033000004c000c401030001c0030000d0c04130005300400c00040c03c0400cc010003003d0030f0003c440c300c00000030044f0000000c0000004130010df400c03430500000050d01000040000100300000000d7330000104311004cc3d3d0000303c310c000000001c010cf130000004100000510040003cc03c000004c0c0300d1c000100000004010c0004c7300000000c004014000300004c00410400500000004000c03c000001100000000700030d04c0400100000010300000c007100d0c44404004004030c4300101c0070c03004000c41c040000440f0000010c000f7300000003000c300307d4510000303004000034c0101331041000007013040007000400d00c0004cc00300cc40000dc11c00c001c10003c040073d03c00000730000000000c000000000c170030fc540040400301d03073c00030000000c0100000001045000d0c3c00010c0000001c0c03030000cc10d03100000001050000d04c050400004000;
rom_uints[879] = 8192'h4c50110430430400c00310111c3010043c101c0340000010003114001100300400331410041314001f13101030411300f00c030c03431d03141010003003300010103d3004131c1f3f0001d0001031040330343414300003301c340100001000003400030003000000d00c103110f73400003cd4003003cd0030101003300130330c50c350303017100034033c0004040001000300001013c0041100f410004150003000403f03000030000003d0005001330430001c041cd0400000f034cc0c00303033300c770300500c0f0c04100100430d0003100030100c0030c33410141d100000033000000400001c01133004400110701075100030f00fd0f001001303030000d01d00f007301c3400111404100c30317c117010030c011c1f000d001000010010f100411044017343000000301031103c00110010300c403f107400c104df3310c00f003c00001403310f1d30c11034003f140f040001000cc0300010110000110c00303004c70c054c34000110cc00f00000103d0c1c0500303000431007c0d11003010c343000340010154c00011011343c300000000440550d005333c130103404300000cc001031001c00040400100001073401333003003000d0001c0d04f010300030301004001000140014c000303543110c140030c1100c140c107100c0010cd001400710cc1c13440c4c1014300dcc3430001003010010730003c055010401001400000c1454004c000475c3331003c0cc3d00043050540c0c3c03004030c00000d30c3505001c001c1c00000330013010030053003030fc0c5001100000c0000c010c3314030c3c331100030000003401000070300034000000003c0df0301043c004040034c4dd0000c030011001000c0030040d0000017110c001004000333c0c30100c100c1cf7740000f14c1f0053cc01310f0c003130103330d1f00100303010700000103c0303000c10001110c00000000000100000103040003000303010100004c01710305010443ccd1c05000dc00030350c3c000400303130300010d0c00c1030004004ff01001500000c3014300d101f3030d3000003000030103010df04f00300f404040050031f4100010133000000c0c070000111003404311014141000300013440070301f3400f1400c47144c100011001c003c0500031011fc004040c01104070401000700c30c10400030cd1c100403004d3000003c343010143d103c004040cc0f3031030140c030cd10f03d00001073300f10300075100c700133300c04301d03001030007003d00001cd00110c030c103004c40f00000c3010044037000010100c00d4000000d0000030cc033311c00f0004f340040003000c1c0100000c0c03003030c0000c3c00050cd000400000300d001c303c0430343430cf3030101004003030303130140033c00010;
rom_uints[880] = 8192'h75010001474c371314c30000000000030301414140cc000000c70d00c3040000030131c050034030003300000030cccd010171f040d4004101000300f34340c1470c000003c51100040000c30f04430000000000c0030101c74300000000000000511004c1f110c300c0103303c3104003010015110000cd40000c010004000003c3307030c730cdc000000404030040c0470000003030004dc1300033d00cc3030340000071130303030300033f00c50313014000c04103130000cc3c000003f034000f300007c0000300d40010030f00033000413d000003300cc071474404c010003400430000030000400001471301000003050000000010110330000000010001100d33c4404300400001003000c07041530c0304c1dc403331013dc31d30301c00c501c001c0340044c30000c000d3000c0030400100000340d50d00000331cc0110300001730043310041441003100017400001d10000030000c004c41330c000c740530703000370c100c000001c0c0350733000040700d1000100504010c5170031030301c00141c100100003303300000047004330000000070c0100c100410300c00040c0c103403300000d01003fc337003103000040c0004430c30030000c3dcd410300130000040343c100030004f0c300104000031000010100000cc300f013c0d30f5501c1d7c100000043030310c003000004004040cc0000400511104310c300c0140770000c4c40300c00144000334110010d0044c1c033400d0100c0340d00010c0103c300107130c0050000010d0303dd3f40000431c30d41c1c703c00300415335730000fcc0000003c1030047c3c30373c440c3330010741354301030030300fcf4034cc04d1043d3c1030c40d4c03300001010c30071d003000003d0c1c003c331c41100c0c3cf404030c44f010117000c000300c357c0050000d33c070003c330c0c0000130c0c10070c04330000300000040400004303001003004c0c04001c0d0c0f700034cc0c07130004c00004043403003f000000341c105070403001101054000400000f11031d70030030000c310400105004005c10701c04300d00000031003c01301410001100044434444000d31014343300033c131104005c103000040010153c304c05c50000030d0c000030013c5d11004334340c0c3cc0474430311000000037000001000005d001000040100010303d00131000100001003fc003001c0440d4100000c30140003030133000370c040100100001030c04033c300014c03c00334c0103c0033f3cc0033050044001140c0000c01130011004403007015004340d07440c0040010010000051001004f70f10300011c0010014001d47c407040c000030000c3003031c0d0c0100c43c00c00003300040140301304305301353043c303004370000010c100c00000;
rom_uints[881] = 8192'h5030501f1030034330300000d0300000c0001070001c107010d01000000100c0000101cc71c0300031400010f0001000c300100004f0cf3000000010c0300000c0c04030330030d030004000d100000040d0003130d00001c1c0d01033d000413010f0430000340040003000140c0030133000c0101000c030c00000003c0010c3414000303000000100034003100130003000000013000001f0000014000010131000f01030c0003030c040004c00d3130300300010f0003c000010700030c0103010c0300730c100c003003000c0500000f00033c0347000000000f0300340101033543400000000300c407f51000c3c30010071000000003000100000003303f0dc10f040d000103c33137030010050c1c01001c0c00c0010100300000000c05c30000fc3003000033100d010037c0410c301404030003003cc31c040101053500034000c3004c00300000000303cd04cf001c300140cd0031000003010300000d03000c3001440d0f0100030307100040000c01330010c1000000400c010f031cfcc101130c0f0003c030010d014700011331001400101000003001cc0c33070114040500031c400f0134000100070f0c010100010f001d00000000030030104004c0030003300d000001031c00011303030f0f010001000401000c0007c100070533003440c701100f000000300100333c10000c0000310303050c00340400c103f1003030003d1c000304100000150340cf0000001c000000030c040001343f030c00000304000400110c03000313040410100d1c04c50300000000004f01000307000001c17d31040300700000140c4013c001000c00000c0300c30101000d004c01cc040000000013000100340000c000010411300000040103000d03033000010000007c0c000007430c014c03c100303d30000c00c000010d0410017003400c03c0001000040c000005010c31101c03000130300ddc3400300f01300c001300001c0010010000030f300130500c030100050304000c3c01040c3c000003000c0c0f0100000c4000001303000007310100000011c001000f001100043100050000030000000c33043f0c0f00f0003003000c00000d000c00100304330000303500403000000003040c4f0003003704300c1005000d3013000c01000007003f010001400005030c0f0c10011100110303030c0010c003004c00030f0c101034000003001013030001000d0005010303015000010005031001043100130501f00c004c00fd00005011c300330c00c30331f40100111d000333331010010cf1051fc000d000013010000000c4004f071d13000700000c00000303f00300003c010000c104000c40100f0000040005300100451330100c130301d131f304000001000000030fd4c0000000c30003000f41000131434d0c011004004000;
rom_uints[882] = 8192'h30000000304300500001000010103003030040c0cc00000011310114014f303001000000400410f34500400013c44033041000c3010c30000001030004c0fc00c000033000001040000010003000f0040030fc30011000d01010f00010f0000c30011400300000c000c0000d000000000000103050003000300000103000001f341100c15000070304000c103103005300000300c43000d3c00d033f733054f0340401000c40400000000430000050003005c0000051c000003130fd0050000000003031500040003c0000053130c0000000000300003030101001cc0c0300000000001340000000fc00ccc703003000033003333c0000040c003400100000c0000034100d4010c00300300c1345000030111304c40000c30c0000c000334030c030007434100311040710100000c030170c00103000003000301010300c000003000d00001000001c3c114003004d0014034130cfd313300f111301301000f10053000330030040f000cf000010000105000011c0000010000310304010003001433013c0010033010300310010015f000f1007001c043001403030004100013c303003c73030100000040010003dc00450f40010cc03343010c004003000004c0c143000000103ff000007000031cf0101303100000100303400cf00c050300c07403000c000040010101c10000c04001c000010000300f43030000110cc0c0010303c0030f000003c30001003f0d00100001070c001005300000c10d3013000000c3051000f00c1030050304c003000f1340003003c00c030000000000700c10000003030103000040dc307440f0011000030300300f0cf00301c400110013300301d30003004410c100041f000003000315300300f330d4400000c030300000c00000000004303c13033400c04c00000303301000c000110000c40530c404c00f1300354030010334c0131000c0410100000c0301300000dc00d3000c0100010000000d003f007c00001004034c000303401cf400001300cc0000343305c00300000001130c000130c0c0000300000301c0c0300000000030c4d0301003000c00c4100000100104104004000000031000010310d01000000031c10001031d03030000003300c004000000030304114301c0330001030030000300011300000c000041007500010010105fd000030043700341c0010cc0400000003100004010403f000004c50000d30400033003400003030113000400f00c1cc1000310c0000130c000004703000001400001000c3003c00f5000010100034c0100130000f100c00330001030103440c000c1c0030130c130005000c000d0043004104103001c10035300400cc0030400103c00400300000310101d04f0044030133300530000c0000c10000130c0003003030030000304c40c00001300510300c0c00;
rom_uints[883] = 8192'h10000100c1400030100c0c0000c003c0031000c0c003001040c000004370c000c011334110030004034100f000000003d0015033030040100000033000000041030030c00030030003c30c0003000073c00f43c00000000cc03c0000505100c011000400c0f0100ff10000017001303000005000c0030004403040c4f300033014000100f000d00000004040000413031000000000034c000000300041000f1c0010003000010400c010300070004733cc0000033013303310c34c003c000034004010000003000300030000031c001044500001c070c00000401000f0000040000000c3c130000000304030c000343005c000031000430000104030000000400000c007c0033030c01030334300303100040003133000050305134033d04100f01001301003c0330003d0414141030300000000030000000d00c010c000040000041030073000c03c5430000000000170c7400100331030403ff103d30004100000c003c0533331450100104c01300001c0303000c00310f0c0000000000cc000000100000010301000c0c0400030300001f100033c1101104300f001000000000000415030100000c0530030014c001000c073c10000c30001500003000040034000000000100100400030000050000000c0c10330104c33500d0330c0400043000010c03300010003000373d000c000010343310000fc0000004003c001400050304301100033301d10004051010000430030c3c11040300c530041f0000001c3c0c3f000000000300000031030c0100000105000c0000c103300c13d000040c00300c0000104c043100003400c00000303130c30c0010000030000003f0000005000403030000041001400c340c03000000000f30000d000033040410000100040100000c030c0c0f03330f001115331000000313000000000000c40c7437000010300c000300007f0103003300030000003cf03001000010003c0000000010000400400001030013001000130010001c030114010f0c00030000400404000031300c00050717d00000c000f00000103404041301300307300130000000c010000110013034003331000f00117d041330f010370f031f0f110c10003d177c000004d030103070301031300c0000100f04003034140003030011001400300010000c010000040400104c003c0500000c00004c3033401103003c001030000104c7000f301300010c00700001300100010c0000d0033030003000030f00c0140300000000c04030007d040c3f430f0010303000000c00130c01130f00000c0000000d000003000000310433043000100c300300310010333000000c0c0f000110c000313300c000030c0cc000001cc001000070300403043f1c3000031c0000100c030c03040117d40101340310000c000003030033103f00c500000000;
rom_uints[884] = 8192'hc30400d0cd000004cc000c0100c040000404100c00d0140000000410cc0400c00c0034c0c000040ccf00000c00010300c000140c00c0c4c4c4000340000d00004c000c0c0400c000000c0000000c000310030c074c4f04c00c0c000140400000c00d004000000000004f00000f1400000c0050011c304f000400d0430cc10004040c404400c031000f0000c000c0c0100c00000000cc000c01cc4401034000000c400000300030001104c000040000000c14c00000c0000300040cf1100400040c410001000c01304000000c0040040003d1c40000140000000000001d000450cc0000c005000c003c00c000c44c0000000303441000000cc0000400000c0cc400c10c1700300f0c01c0004c0100000f4c0d0d7003cc007c000c030cc000030000c0003004000c000411c300c40014300000130003000040c0ccc103430000000300303001100440c3c0c000000c334c10040000100c000f000c1700000c0000440000cc4440000003040c0500000000034300040cc000000010000c000000cc0003c3000c0c004c00040005044310cc000c0000001000001004007043300c0c0300000404c000000301c4c001175c00c040ccc0100300000cc40000500d00d00440000144004c00010000500050cc4010c00cf100000700100400400030cc0000030000c0004040000dc0440f400005000cc40010043c000304cc0000000004c0c04fc10010c00005000c0004070c0c04007d03000004c503c00400001400c000c00040cf0003000001400000c000c104004000d04c400000011000000044400f0000000030c4004dc001c00c0400000444c100030000000030ccc0040c3c0000004040400300043c0400000000010f000001000303001030d0c00c0004001404100001000c00300cc003f3004c034317030300c3d34300c00c00000010c3300cc04001400f0000000030c400401cc400c005000c03000c001100000c0000cc00140000000000000c000c000f000400000c0c0c05000001c003cc434cc40c34004c00140000440000004c300000400000030500c000cf0000140cc0cc4c400000cdc000c34004c4044004050f00110400f0010f0440014c00005014034000000001000c1004030400c40000000cc5300f0000000400c44300000300c00440300030c5dc04000000010dcc00c04c040001010c0c0040000c040c000150d7000100044000430000010100037300c000c0ccc00001c00340001300000c04000340c00c0000004400fc03004103000c10c000c003040000000c404004000000000c4c40007c04400c001000000305441400400003404000f0004f04000c0c03c000ccc03d00400cc4004c40c10440004c000cc040000c0c04c3010c00000010cc070000010c004c04000400000040030010c0c00f0000004c000044cc03000100;
rom_uints[885] = 8192'h43c40c0004004d14000100100c00144c0104c0440100000c00103c000400c010000c033110110c000015000c44c3c4014c00f43410c5c00100d00c30d3003c1000170c4c000c04000000100030300c3004c304d40033003070d74033040100300f300400000031710000030ccc0433000000003fc0011c33040404f10717c000c4000034000d003c00000c40f1001cd00004000400331004f0304400cc151c10c0c0303400303c3101c00d000000031404340000000405d405d4f00cd4c004004c00dc0c3401037341c030041030c04c01044c00300f370c003003040003043400000030000c031400df3c35140ff100003c0c40c04303103400040c04000410d00400ccccc10c3400c0040c40c00400300c000c70d000103ff00001d400c71000030c000c04000400c30f300400340c00c10000c000000000000030010011007c0470043100010dcc000033300004000040ccc0450cf03c300034000003301404d01d00000cf10300030000000470400304c000000c000000305c3c1000c0c001140d040000c00304000d00400000505000cc0c100000000317d030d4cc4000140c0400000c401030310c1434100c000c00700004c0000c0c043cd01434c0343c0400040c0004010c0704000c3c14310d140130044c10000cc01400300000470000104cc00c00c0000fcc0000140404dc0030400030000001000c0000050010c130003cfcf00c000d003010140c0c00003c3f10003c1414000010c004344c4c0004047d4cc000400000c3000000110003c354040c140005cc001c070400330cc0d430000000c43c0000040c0370410c14004c300113400c0cd000007130041c451f0404c50404140400700030c0700c340030005000300c00040100c3700c0000000c11003cd4373100140f10113cd0c4700c003c0400c701c004000f100500f1f4c000005015dd0d05fc0c4c004c1030d0001c0301c0d00000545c00040c0001001c013000000c0f3c100c14703000005d00441300051400000003c0000d04700000000000040c00040004000400c3300c004d04000c0c0007cc30411cf0347104130070000c0534001003300130510c000f304143001034fcc000c0010004000c1014c443cc303c033030053c0c00010c1041cc30c000004d000c00004d0c04c0010c10c0c47d0401000c040c0c0cf0cc0007100000c3dc0c0c000d000004340013100000000c10000c303c000c0c0003040ccc3d004c330c0404170303033c00441cc0000c00013400d000040004c4000c00cc340c1000000000000d003c1333070c000c0c051c10304c000c00ff0000c01c00000110030004007d711c470ccc04040030304c00330433004c00f400c03010000105710000030ccc0c1704000010401003340000100f0c3c0004003541300c000c40303d0cd371043c0004;
rom_uints[886] = 8192'h3030000303100410003000d030070103103000330c0000000130030003130010000f031c000300000103001310400031000401d4100107303000000330000000040303000c030c00000c101410044000000300130110000103041d030400c1100f34001000000007001300000000331401001f03301300000c0430050000000c100100013300000d0304000dc0000c00300000000007001003010004300100103334000000003300000000070000010107d00310000001001003034031c0000300000100000004100c3c13030c0370700033000331004000313003101403000013100410000000004000345d1310100c0d003170c00000000001000c1030003034130003100c3300040300010001033034030101003300c1141000004f01000014000000300100400f0003130004c00330040110000000000f00c00000c07000341c10103134100400030400000044000000000000010003c0011cc30c01100c00c1fc01f41c010d10040410001007000c0d0013050003400f3fc010003071371000000cc100003c0011c3030000d130040c0d0c000010000f00c00410000170130400030d100cc0040000030c1004030c0d000000d001310014000030131c1010370000000c140044c00403311c010d300c000034c000010000000dc40c303001c0110000fc13000d000400c0c0cc047404014c304130071410001003000013070c030000ddcc001030000c0c000001100d000cd0000400040c333fc0000c0403d30003313311000500340030000c00033100000304701c0000c013100031c4010000000113000c000000000000000031000f1300000003100004001003003001000000130c000000104104000400140c0030001c0304010f000003300000000100c00001100005001001c10003000300170000041000d0000d000100d300040000040c10c430000000117050cc3d030000000003001000000404001003051000003d00100000000103000003d0150000000d010c7103013403030403110110000000070003c0c043143000030000304333300000003000000c330c0c0710010011410000000cc0000000c0071000710c3100030004110054434c00100c3000003000000c4c3130000f0003005300300c4c3d43030300100040030d044010300d0101070003000c0c0c100f100d0c030433301000400030010001005000c007400c053003100010010001340000000030000c00d0041c3434c003003005f03f0d034500001c000c3d173d01040cc01c000d07010031000000000001000000041010010000c0c41c30000450003d00000010070000010100011f0000371010c00005110004031f0304030c03d000001300000000000300100510500f00cc01000004000131001c00010040cc000cd003070004001034431d1f0003000000001;
rom_uints[887] = 8192'h400000010340000000000340040100300000400000d3c0c3fc4001003030c0c00340030040030000c0004340045cd14c404010344c0303c04000c0c00000030004000003cc0000c000c00000c1c00f4000000130010000010000c30100cc00040000010000040000000400001400000101010000c4c340400000c0c3c0c003334000c3c00000c3400101114040031040c043000000030040000303010404000300c00140c0c01043c00000000003000c01c0c000041000400001c300000040c0c3cc000301c40500c00c03c00000040100c0004111c00000c0c0400c0000000000040c4303c0400700c0c1005104444000000f0000410004400040000003000000c040004000415dc00107c140430cc0c0c1c0c33100030d4003004100434001030000c00000400004c040c040c000004101c40440430040c000040000000300300140000400cc00400013c300c0c03c0000c0c3cc000c30034100014fc0c14040000340000000004c01000040c0000003c7c001004040c0cc4c0000000c040303000000c000004503c043c04000400000400000000400c0c1c1014000c0c047010c1041040000000040400004c0c003011303704003c0403000c040c0c0134030c004014301c3c040000c00c00013c00000040c05f0300040404103000700c000c00c03c00330f300c00c4c0000c00100f00473c0c041000300030040003001000303c000c0c00301c3000cc0c1c0400003cd73c30047c0c4c3c0000701c400c0d00040010410010000c0c0030000440c4104c145c043004040c0400140030f0c030040c0010c4c4000c00444034404000000c000400000414001c000c40300c5404300400003c003c00400010340400000c0000001c0c047c10041c0004007004400000140030040c00303c730400000c0c043400f000c404041c04000003001c040030040c0000100400000074004000c4304000401400300c0c000c00150c050c3000140030000000040010000004030c1cf00c300c10300010144c0000001000400000040030100c00c440041c00000c003c000c00304000017c07007c04300030000c304000f0000cff000c3000000c0c000f040c100400040d00401403000c170c001c3c00100c0010000c14003c3c003430001c00103cc0dc003c04000c0c00000000c0000400000c070c00c004304400307010c00000000cc00c100030103000400d000c0000c030c00004000c04000c0430d030041404140000000440340000c0103c000c303000343c0104040c047c4c04000404005c330c001000d000003000c0000c0000040404000c04007310000c141c0004000c000c00000011040c315004cc003500040c00100004000c100c700c003004340c00003c043000003030c00c0004303c0040d7004c3c0040040050100030000c003c4100;
rom_uints[888] = 8192'h130c0000404cd00044c03430130011c003c0c4070000c4c300441330303c0003040c0c03004d0007004c001043003c304c100004f0014417040000000c10c0c700c04000c1c0000750005c70fc007113100404100043034ccf4700cc0044c40c404c001004cc0c0400c05c44100cf04c41c070fc0004400100f4c0000440000070d04407010f00c400c0030000c000714000400400000c075c00f001c0c40041340d0100044f01cd0400c770c0000034003f10400040000c00430440cc0030033007000c0000c3c1ccf44010c004c10010c1c30040c03400f00c0c00005000c0c0cd3004c7130304400c003c01c04400000d40300004000c5000000043000000c411033f40440c4001040040c0ff0c00414c40700c4304c00f0070fdcf05000300400f0030300131300533453cf000005c0104f140104000c33c005001014d000ccc445d4c0d13007c000010c04400000000c0000043c0040f30017c400003c30400c4530c17007000c7407010000c1cc3c0c0000300400c437d4f40c0004c0c107140cc1d3c0001cc50030400c4010413000400f040400440f7c0007c003c3c3010c000c101c00300000c0103c0f40030f000c0300000741000000300d0743c30f4000cf400c0410cc1c000cc0070c307003c00cc003011c043c040c4c7410cc10014430003d30010404f00000300340ccc4cc0c00cc0044113c300504c0cc3d11430f3c40005c45cf13c1f13f1c0004050c04d030c000003007c303045403004503110cc7140100440f010c000040330001001041107010c4c1003400100400300100c0c0000c4013100c344f0c000001000400000c000c0c30040d104f300000c00c07310031f00030431cc00750304f050c1505d0040000c000044ccc0440c34040c4c400030c0c003034003cc1000c00000403440770001ccc0c00070400cc04000000001000f00044d50004003470000003040c05d003037d0044000003004f430c1004040000c00f0001c03000c100cf311f713f010513c3c005cc30c0f000300430000000c000007c04c3047304003400044cd400000f500c0c0700053304000c004f0f3c400033dc0ffc0f30400c0cc0303400440004f0033040040c045000050c300c50004000310114c00000003300ccd00300c00c30000410cc0cddc3c055101030000c1400c31041c010040117cd04400004c0050030000c400c0000313cc40004fc0004cc4c000cc04d04f3f0030c17003430000c00030000434f003000400700dc0c00c001001c0404040c01f10c1c4001c301d0401c3004c1d3000c0030354130004034034c04404003031004340131c000f43003c000cd700f0c30c004c01d00000010d0103300c0003440000c0c05403c04c00c330c7c1540f10c00f437f3c0474f0000004cf00030040c1c000510c01f00440dc00cc00;
rom_uints[889] = 8192'h10000c00d010d000cdc00000fc701c13040114c0000410f00040330040300cc0043034000043400010d000430353c0030033fcf4d00c0007d4101030c004700c00c000f000c01000100044dc03000034103153001340c510304003000dc0000000fc0c110000303010c07100000031004000037030400000133334c1100330050f41d4001d0040330703305044c000340510c03000000f01c000c0c3f310f040d1017300c04c1000003f30d0c04030cf100cd010001044d0f0c0c3710000000c41ff01303030030044d330130030f0730031470100041c0043030530f0040003300000043d4400000030300110d0f10300000700070c000010000043340100041cd000303400030f3030003511400000f3400040000c1140300000c00401000f00053000c3001c00040001100c0013100040000000101400003000004c0530007000c0c0043030003000000003c01000cc04007c0045007c3f01c0f0f010c341103033c0103000530c30040443103c5000103700700f13d03c100300040000c143c3d0333314000000010000050cc03c30007430000010400d0050010010100cd30000000504500400000c0f01100030c00313c3cc1133004000007000c04f00003010103c000333017431301500c001131c14000001045000c31c00fd30100c0100d0c1100030100435030005c1401cfc30c0573c0c43041cf03000c44003141c0074f4f300310030130c000c11730010043113cc30131000404700130c04140300530cc0411c330000c0003070300003d1cd00000c10c015d34c05c100040400c100013110f00011030003c005300001c1003000f30540300003005c000000dc700033310031153f04000003300030f3000c40cc44d70000c01c00050034300043304001000c010c4f4450140f003f00703000c44010cc00033d0071d00c004c7cf03330050c130c00411c03c00004000cc00c05000000140070c0041000141500033f10001000030400470001000c00301c0c013c0030d31000331c0377401000cf104100103001d1c0d0701030004100f100cc14001300c3f00c4c400300470000c0c004dc5c0c00c0f0c00701003cc030007000001c0c3304404030003474040000130503010cd3040033c1700010c1415000fc0034314301101051003310f0c4430040fc0000300030034cc50033c51551d000f0000030dc004f001310c3003fd00000000003001c00c0040cc03c1d01144040340100000000c5f4000003000c3000030001033030100f003001444000003d0340000d3c1500070300d013c1000c003044100f00000300c041f0007005c3d00010100001040000030c0130000f0c00c0f100d030c0f000137001000000c00c0003400440c13700000540f010743070c0001300100070cc00314431000070400cdc4044cfc4d573403103;
rom_uints[890] = 8192'h300c00003c10004003000311000053003450143000c7400030010001c400100010030c141500113010000d00000c0033011c00033cf0f50010303010000000c000400001000003100010710000f004030030001330100100001cc73000040010d30403003030010000450000004303000001130000045c001d3410000333000000500000010040000c0031304c01cf150000000000043340030000c003001100f4303403c0103d0101c000313033110000c50000f015130711001c041310300014003c004000000303001f00d3111010103100000303000044000000300040000300303f00000000040033004c30030073f11100010014004030100040001cf30c030113101000013000510c00010030c001f43731030c500010000c30330000130300040100070300341c01000300311030f31f11f400000004c403000000000030030403500031f000f00c003001cc33f010f7411005050cdc1f00030c000cc41000400100000c140003f37330c0000c700000c000c00000000014003100c1000000c1533001031500000000d04f1c00013000040000c4f01501300c000000111000703c00300000301130c33044000003310000040c3013c1040000d4301011100034343d04433f43000300000014101030f03300f00000047c00300c130040054130153033104100c00004300c003030001050c040300140000001005303001c0c4dc341000cd1c001f01031000330000100c330c003010c003c000403c30c0101004033150000400c10000150ff01300300f5100004404030430030403000100330000000c00fc00500100000d0140470f0d14f000100c03000100000170000407c01400000003f0033300043c0000010100054cf0c0c10000303105000004000100114330040011010101c011101103c300c3000000c4000c0c000305401f00000c0411430100030d03000103033171000000000431003000033041f4c00300000000c000c1000303333cc040051f0000000013000c03003f00010040000030cc3001031033000000c0c1500001430c033000000d330100001130c00344033104310000c30040030303d00c300c000c0103000000c3030003c40441434401010fc3700c1103f100000103130cc44f1013010130014f3030011c40001105300000c0430000011530300010034004000ff1030400010f0004011000000c0003c4000030300140100003c3030003130003f00003fc0001000105c03333000041000030000d0c503c305300f7001003400003030c4001c4c1401f04003c030000c4f001100100000c30c30001034013130504f00001000000500010140040010f01030f103041030000c01003030ff043001000000c0101c000013144333c40010000007334c30033c30040c3000300000140310f0f0c1c3140cc0000000;
rom_uints[891] = 8192'hc13100013dc1031300030310030003103300010001010d10010701000043300c0f000450d04f00001c01100007030f43300700c00373300d00004000c0c3c0000f0c111d000101010000c0000000000dc03040300c030d7f03040c4f40c404051131030301010440c003d1000304d4040cc030d001f300070304010343c0c001031303004403000d00010041c003c0f403030000000040c4cc04000000c001030c0300c4c000c300474104c30f07030403cc400000c340030c07000c0000300303c10000000003c004030303100000330000430000011300304f00c331f500cc030300030000010003010143007d03c000000043013c00000301010c07c00301000f1100000301c00171414d00040340444c5c00c7c30500df0f074cc0f7c0f0000dd0000dcc00c30130c0010f0041030100033003000c0004000c0340c001000100000d1400c3004307030143c04003cc0c0f03301d00740c004fc0400307000003000100030c7000f1030434c0000100034000c40d010000000cf1c0000cd0400c03100f10030301300fc01304c300040300004c0000000030000c03000c0700404107010c03c00004c043000f4300c030034300cc010100030c1007030c001c34030000004003d00404000d000300000000033000c73c40040304c0c300050000c3d100c403341c450c0c0003000c04440711c00000c103dc00030d03030cc040c010073c03014c730357004550001000370700000300cc0350000c00117007404000f04701000001cc0403000c500100c7004000000300011103f100050030f4c3c00303c10f0104cf0400cc030331c00fc0000010330f05000000004300fc00c310470c0cc34d0310c0004301d4304c0c400300000301c0400cf40101010c04d004000000c00747000c0304c000004c0d0100000c0001010400530c004040030f440c0d5c03c3000740030001c04000030001c000070100030c0000000c05030140040001000340000000413c1c00004300f70c4300c331010103c001034000c00000000330c0000130c7c10300c300001000c44f001f00010077130340040cf40000100c0f43001030000000404401304003010003040d043010000d0000c700000705407100044c00100f000170173007400cc100403010014340030fc0c3114000010c43000001c1030c00410c110104c0f500c001f10300000000030c00c0c0cd00035007030d403701400103011041000741c00110000300c33441430c1c00030003304300cc04430010cc0cc04100f000310003c0030303104001300131000300c10c0001000f001003000010c013f100011000000100430f4cfcc503010103030fd3100c0000031000c100004500000003000003f5000103c00000000d00c3100c0334040000c0c00f000100000c070c0c00430101c0c0300000;
rom_uints[892] = 8192'h300010100103c00400313000040000004070c100000057c0401001c003c00004010404100c00d0133000001003f0000003003000df00001000000000100000c0131c3040001030030300100004c500000c0740c3000013d000c0030000000074c00400101003100000000001004cc4000c300100c5c0004710131000005300c4c0000110000400000000000000400000010000c0000030040004000000dd0431100040011c10040000000000030c05000c4000000f0000000cc30000000c3000c00000000000100000c00f3100c40100137100c0000107c031300140c00000100000000300000c0000f00441c000300c00300030040000704001000010003000c0400000703110330000400001005d3003c01000040c0000cc0c300c0040133100000400000004c000310304040040001014007000000003f4101030103010034f400000f00000110050300000c1d4c0010400100c0030f030f0333300100004004dd030301cd00003310c0033000000001c0c0310000010f3403000c000000701c74430010140000310000c30c30000001000003000d010101000c3000c007030000114000001000000031003300400300311300c4440c0010003311040303000040000030004d01004300c3000100000304100d0000040010f000000101070100003001300000040c0300000000001c43070000030c0c0100110c000400400f00010cc053050c000c0400000100000c0110000c00011004d4000000c300c04100103100400000030f1f031033043101000341000c5135c4000000400c0000003001cd0000000010c30c0000000000033011c030000301400030030c100c7400040000000c00304c301100400d00004000071130001000d00000004300004003c0000c0400003030303100d3010c4c0c01001c000c0004000000304100c010000fc00c01000c000c0300100400110000000010000c000073c0000004004000400004000c41000001300030033005104c000103100040001005ccc10100300000003f000005000c000300004000010004010004000030000003300000001130000cd3000303000433c04c10304010c0000001070000c04d0300030300000dc30007000000c000000000100c000000300010000404000c01330000000300d10000000c300c0cc0400705510cf00040000004030110110c0530030003000000001d00030d01030440001c00000000140003000c0c400403400000030030c0003041045100c00001330400001001001011340c10154d000f0044400c0103044103000000c3000f0103001030000007004c000cc00000030000c00003000010004c00000000001d010c0304c0d130300000000000101000033007000033000c000c0000030000013000300000c0100400000300030010c00c01000100dd0000;
rom_uints[893] = 8192'hd1300301c011000003005c00010c000cc3c010d30f40000001f700000443400000c3430100c0000c330f003040003010c30c1cc00000350c0040304041d0000c010411c000c310dd0000010d300f400101401000c1731011343ffc75013dc3c03313040407d0004103030000010044c10005f0d1030503400cc00cc301400c0f0134510400c0000000000400000000430170000005000c47000700034400c000cd44000f03040d300300300c30d30d0134050010030dc37d0101c4003000010004040130100100011df005000000f70000c00400030337cd10dc3d00050400c0c0010c01030000000030c370f7054c03000030310011000101050001000004004fc43004100000147d00053003500000c33000000070300401304303731003000730c00cc3100307100044d00c10010d00401fc0000c40030c43c0d310300403004cc4304300000c400037400001303401030030073043f0c40c7303303100110443571001000c0305300cf30cc04300cc3c0001010503047c03030c100300100cc0c10f7004337100031300f4003750c0000003000c0000d03c03007303f00441c000003000c00000f4014001f030041000347d0d103f000003430001300000341040000c10011cc74001030000c30d044133001c000300cc10010003df7ccc100300c00001cf0d034f4303710c4cc44c014f30040c043343301000037c1d30017000cc00030331031d0d007f0c0340004700000100507d700d0000010c100000c3000130104040030f311d3003000405104001004040100f00ccc1300011004300cc0401000c30001c30cc07000300d101404350340000370c040113c01d300000000c400c003c0034030030000000000c300300041d00d3d0c00f0c3004c01041c00000030cc0d3001dfd01010c3400c00001307ccc040f1370470df10400000101000001f0005341cc0141c1d3c1070c00d0c0300cf03300c0c0013c0103510c4f030000000001c0033000ccc0100573003fc0030400c0043f0371401c070000043000000d000003f11410d401f350000400c0d0000100c00007430570150000130f3dc30340c0000cf00500c10441043040c0000300337444400c001005c040010370001000410105007334000000330040c4d5140000100010003101000300300105003440011000030500000000c30c4fc11100113c0d010f1503000100000f00040004c54050c70370030003011407d1001440c000401c0cf00137700c45001f0100c007310f00510010003d0303710301144cc0ffcf10434433040003050000c00070f00400010010400f000ff00040414c00c4004030000000f3000f454cd3000f000000010010c04300140307000100001c033f000530c011cc0d0004034f10000130100300cd0c31fc11110000031cc07000300c34010040100;
rom_uints[894] = 8192'h300000c1310c00c000d00000000010034c101040c001300000c1010000133c0030040f0c10c40000c444c0fd400030c34314fc000434c001110c003000400c0c04030d300001000d0000c1430000c10031404000c30cd0004c1c700c4010c0c300100410140000001c0001c304370103000033ccc10400001011037304000d0c0d0300404030000500000041ccf0003d00170000003004000701000000503c013003003c0000040100300000730c0033010c0500000040c0d000000c130f000f4000000100103000404500030040053010c0410100c00130c0c3300100330010011000033010300001c00017c7ffc4101000d4c000740003000004c0300000000c40010000310100010d00f103000f7037440441c003000df0c100c30070101c0001c3000450c040004013f0c3c00000410340070031000000400010301031000d0100cd01000300301d1c01400034d0c0033c1040c00030101003700000000005030310c041147c030001d00c0f1fc000c3073001d04000114100000010f310c40313c001303004135003400c101000000040000400101300440300100700000300c40001004001413f0c00500c400400000005070c0d0040000040470003010000000003400044001c0000c401001c0003000051c14df0000310110c1104100100400300dc3c00043c0d00c0000000010005114c1c0f004f000001030300000000001f110001c33134513341000100c00100000c0133c4010300454000c104040713c0413000100100c0004c0000370100031000500000050cc00f00000c0c03c3040c10400fc0010fc03400100300704300304004c10c40c003401044030c10101004d0000003003040c30c10011c03000041000dd3000430070000003170c01030100000000c0cc30133c35030c050410000303370c300050c000304130014d034003011340003c30fd50071010300000333c01040d5c001143100000030c000f0300000000730411000000030300000470004c000000000c3c3c0144c43c000330013d00000000103030000400410000f11000100040f700010143041400c30003003010071400030441330010001010010f331000034c01d000c00000144050004030000d4000c30001000010000c0ff0c33000000f7c0001003140d03740f10c00000000054030000400000054331c01f500c4003c01c00001007304101000357033f00c003010037d0000300010c0000c300000c010c0003004c000044d050d70000040000000040f01034c57c40d04337440100030c1000003c000c30c0c13470001030c7000040000000010074300f3300010400704100c70330030d000031c301000030c0730040070000c0000107000040300103033c00000100003310001000400f01000c01000300015030010114000400d000011000000c00;
rom_uints[895] = 8192'hcc0030404000000034003000031033004300000cc010c00000300c004000403300000100c0d000705040103000c040f0000000304133000f0040000010000400007003c00000000c300043403000d01301110000f000c000c04c03001030101000d014040100c5330000040000300510000400040010310400031c3070100010400040f0c074000004000010c5330c10010000300030c0000314704011703c407017f0000000043cc0d0100030d0c000c1000400000f004340000000003040003010000000000000f0c0c03000c0001000303001c0101430f00401c4100433c0007300003030003300d030d450d314004400001030700000c30000700410000030330300f700000000111004000000c0c0df0004001dd0010c4000001000f45030f03000c0001050001c000f01003010c000c43100400000100000003c00c000c000000000c05700c0c000003010004000407300d000401000103341d00c3000c00003c07333c40030300010003000430030000cc0c0d00001d0c01c00000000134000007300003004003000000014747000c0cc00004400003c3030c040300040d344c0403403c100f00004010001331030c01330440454c00c000000004cc170000000fc0000c030c003305304700c30400000c030c10030300000c5f0d000000010333001000c300013111005c000501110003040f0000040004300105003fc0005c004000400f071d00301503c001030000c7401c3300000c00ccd00c00000000c00c05000131000304000004030107304000033400c00530033000037003010000000000c000013c10000303000011000000030c0303400001040400010300000c0140000000000c0000010d0105000103040d01004000c700050f0730334d0310030010c10700303300c3070003004f0c014443070000001003030c003000100d0000044d01470000cd0c00373c000003070c3005040c03400000000001000000000000000f0c00000003000300000007004103040dc00f0fcc01030300000f010f03030f010004001000003303000c04c00c030000300100770003030100310500003007c3000400010054000100000104000400010c0d30000000c500000c34000d100f0001000000040d33030101400303c3730001000033000400410400000700c00000c000000c0001010000000100010c014000cf0000034300c0000730700f0001030c100004000c31000700d0300f3c001041000c100d0000040107c03300031004000031030303340c0100dc00100c000400010000004001000510400d0c0c05030100000000c000400d051001000000000010c0000007040101100003000040c0041f00f43c00010003c0054000000004070103c0000c00000403000300000f0115500000000040030301000007014c0c00000100000d000;
rom_uints[896] = 8192'h7400c0000000000513000c44000400c4c4010004c003f0000c0c00c50310c0c00003c004000000c44010004300030c050300c030053044cc13000400034004004000c0f1c00041f4c00001cc404004404400400403c003c0304003c1450440400145044c710040c300053000cc0100030310350040000c40400000c01000005003c0cc00c30c014c4c000f0000000000c04000000000c00055c01c034000cc00045000004c0c0cc001c000000f00030000447040000cc0040030030f0000000040400005000f4cc00000c44004c403c0c0cc00c030040000c01147c04040cc451c40400000c3c0c040000f14400000c01003405f0140000c00404003005000cf4011000c0ccc0000000101c00000c003051001033545000043c040c00500400c00c1400040400000c0000300000000103000c040c0c000000000d5004030c0c04100007000004000c0140040300000c00040c0014440c100cd13c00004c000000003011ccff043f0c0000000400005c000c01cc0c000000400f540cc0300d440000500c340000000450000cfc000033f00034000c00040c10340ccc04040000043c04040c004c0100034004143df1011400040c0034040500003c000c0c0504510c0005004c34300000500c50004c3000000c00000040340400000004c004f0030007f70000545400040c00040000f00004c00c1014000000040000c0040000c0003cf00040000010cc4034111330000cf01004000044c00000f0004400400c00040000c050003000000404010c0001045c04040c0000000030c300c40004cc00000010003c0c0000043030000c3000000400ccc000c00000c00005000c500c00c5c0001c3040040400c030cc0100c0c013040030000404043000003004c0000014001401000004f0f400303411103c0c41cc0000fc0000000300001130001d030c000000000030000c003004330000041030001c0c0000040300c0300400000000000c100000003c000470c01003cc00030c404030f0000440f000c0300301c0000007cc0000370000040400c44cc054103cf000000000300000540400040cc0341410f00d000c4c00000c00f00404000004040f00401504030000050400000ccc000000103050cc140005c0000c00000c043cc00400004000100dcc4000540004040400000c0500000c0c4100c0040c03000400043fdc0051300031100c0c300000400c00000c00045001c400043c000c0c100400145003fc0c0c040037c04001003000000c50f0001c143000c3fc40003003501000000c00050c30c40c40005004300f0c00000030003004030040000c14003000000400004c00010004000c0400cf003c40f000500000000400000c000504003400000c345c0c0010040400040c00000d000c003001040cc000005c00100000003000300004000000000c;
rom_uints[897] = 8192'h3c0cc0000df3c3044d430cccc3c004f33340070d000001300004c3010400c00000000704034300c3100d00000c004300113000010c440733000003000c00c00004000003000000000c0004c3c4000007c0c001000000003c011cc000004d0c0013050704100c010c0f005000030350000000f00510000f0100cf00003100004501407c01040030100c43000011030c000c070003000000000100000007000000004f0000001c0003001304fd0c010d00c0130400003fc300030c40003000000c110104c300c04701010000c0301130000d41400000000104003300000143000400000001403f000000c00035040701c0c533cf053000000300c000030100000cc4c3c400300000f0010000c00001000031030cc10000150c3fc143000101403c0004000000030040000c40000c00f140054000010cf3000000030f0c0040c0000004000500000000000000001d010c03040401015003030c00051c3c000c300701000000070f00c000004001070c100000004700c000400000313f030031000347000c0003030001c30000c00fc40000330000000000004c07740c40100c4c0000f700031005000300010c0100510100310003c0ff4c00111c00070100000355c35400000003000040405500000433005700c30100501000010cc3014030000c0000c1f300c0000300d30301000c0c301330300c0000040343040000310f000cc4040040000004000003000f400c0c141004030001c30c043100c4041c3473000003c3100010c403000040015000040033030c0000000013000f0f01c3014c0d030d000000c00001040c00f03c0f00030dc500430001403000040c54000d5d00c000000001001d000103c70004001043c00140000f0003143030000c0110000000000101030c4c5c000010000300433f4c1100000000300c40404c000f0c0d00001404134d030cc1000100001003000100300c0000430000f3003d0000140c004100000c0000010c00000010001c3d0003030c000d043c034001304100c3c0004000054401000005001f010500703cc05400033f330301010330040003030000044043000c00031c01000c7c04300003000000030c000003040500004c0000c00d010300f143c0d50004010000c40003c3404105000000000104003300150300c03300040000000000003d0f44070f0000000140c0000c4c00000c40000531100400000c0401000307110000000000c005c000700100040c01040000cd411105010f740000000c110d00430c0f000f10010313400414c000030c7000c0000003530341100f0000f0000100000cc00001010c0303000004000001000007000c4c0011030f0000014303000c3300044000400d400550c1000000c10040030f0000c30f0f00c40100030501c01000000d0000000cc4000100000fc0003c00000003;
rom_uints[898] = 8192'h3311000700dc04c4000000d4cc4010404c051530000c000143c10003440010000300cc0f0c04017030000f00404dc0040107317033404c51000c007740d0704450c0d300000030f1000101100cc0c000110003410000544000c040003c4cf700d4c30f3c03070045013303403000d0300300fc0fc003c40041000003c30001000d151001c400000c100041040010c4050000000000c000c7dc00c0c110c0c040030000000040f030033300103c033000070c0000404143400000130300000000040c000001fc40030c000c41405c0c0040cc441d000c013cc37c0504f40f30100000401335c00000cf0030cf000300000c0c01441000004400000c073000040310000417001c04003404c047c000c00ccfc1000370030000c7030034c100c010000000d00030cf03007103300c31000c40004340000dc00001c3004070c000c17000040003c30100040f0d340004004043100030103000fc30cc000100030040c1cc0134100070c340cc47c0d0000003c7000040003c0007331000030100407000000340103001370100c1503043000000c0441000d4000410017003103000401d0000710c00f0004c000c10f31741030001475000030400c745001000d30400070000044000400000004400c000f74f5000035004007143000d000d1430033140053370c5c3034004c1000774000000000403dd010c40cc304000041c5313c104c0d400140c00c001d0d01004000704c400340704007d0330100ccc04c000c31cf0040334005500403000df00144000040000000100c3c353410010007400000300011c000c0031c30340001051cc00110000c0050001103f3f000c00413c01400000f400340340000fc00000000c44000503c0301710cc130000400000104005430d7000000004000000000d000340cc11000000105400c07000f7c470103307103700003030c330104cc30f000000001001000d40000c404300007c00c34c000100000000000000003343c340400000050c0c014000330503034040004000001340000c040101000030170c0010cc10005d03014000001400000d0004000303c400001cc0055400010c0007700101044101100071100000753303c40c03033000041100000d041350400100004101030c00330c13c1c1f0000000010c0010cc0c41004174104c3c0700c00105001040cc001dc0c00340010000300340010003040c0000000400c00c41141070004100401000c0d3d040450400430d0f01000130000040f0c00500cc01c30744000000c0000050000303031341d3c0300434030cc00000000000040c0403000400004c7134070051000030000001000003343000540c70000c1c001003403001c0000400000c01000d0100c0c01f514010443c40c30300704040d4c00040003330f0410c040000400303000f1140010cc0;
rom_uints[899] = 8192'hc0c10100000cd34041cf00004710000100701000301003c0034300f0c340000100114434514300000071010403030c31f11033f40041004cc00000cc130c0d010000330f000010c0c0004100d000404003010cd3f00d7c0c00330c0c401400400c314300c1f0000130307d0040030040fc040305000440c30004f3c4000c00c00d00c1000c3c01c30103000103000c033003c00000104043104100c100c00f03030c030040004300c3004403000c001403004f33000000100c3104003c0000000103000030004f010c3000400ccc340000cc45000131000c41f1010c001001d7cdc003c00f000cc0030c00d301071c00d054001000c0000040000044004003035403000403000014030c01f001040030c043000070434000330000d51c3104034100070000040430000100017170c371000f0c0003040500c0003034305100c3410001030c0103000103070f0000000f0f43c100034cc0040d01133171c34cc0c0010400000113cc000300304000043dcc0001030010300000000030403103034743050013000010001005f03d0000d0030041c0000043c0330331300100f00103030c40c0c7004100c0c31f01c30c014401c54f0c10004101c0c10030004307000000030000010307000030300001401010100000300c000103000000c00037000303d40100f0cc030f00051000010030000001370f0003c00340034100033110030003073d4000400007540040000c0000044001400cc0143040307104050103404f4000000c4040c100010300043100030000001303005040041013000c3100430330040f000c400303010cf0c0103100400300034030c1100304c1d0330f000d03c3c030fc0000c01330030001033300400c00007000000000000cc0010340500d0c03000031f5034473010c000f00c1304030d0304c041030000c03c073c0130000c000cc31101300c014130000440c03c040cf007c430013030d400c3044100000000000c0010c0001030031c3035c45003d130000040000130003000001000f00404c010100400c0000034003040070100304010100c0c0043501c3001300400cc0030c0d000001c000000100010000000000010000400c0fc0003f00030c00001031000000100403000f0c00300c4101c0f540030c44310000310000d00303c000c0030400330003d31100003000015fc54003c3c0430003041000c0c0000300030100430f400000030430000400c03113034000004100055041407c010553000000030140c103cf00000003310d00c0c1f30d00f00073001c0f0000410000003cf100001c510501400c4431000cc0031000c0000000130001c00d030040cc070010c147033000f4051301000000400001c30301c011cc1000c0004c0c004100040d0cc10051000000003c04113340000001100f00c000c710c00000;
rom_uints[900] = 8192'hc010c0c0f01001040000fc0c000100f40c0054c1301010003000000044443400c00000015c30033c44001040000040034c00000030007c00c400004341000000f0400000131000000031c03400cd400000303014034000007370ff000c0000000401303030003400040cc0040014c0c04cc01700100003300000c0003030c3501c401000400043000000000000001404c0000000c0000d3000101c07000000000000310004000070003d00c05000cc00010d0c00dc3003c4000000c014000014740c30004000003000040000304000c030d00430040c1c1043000030013000004c00104034c00003f0104c0c30f1040004f013304000001030700cc104003400303000304001003004c300000000300c30700040cccc04c13c001000d0c070301000000030040070001cf0350010000040003037000040040000000000400033300cf00000400070010000c000c310cc1c004030403130470030d5400040000000000370c040c0400000f0c1007030004c0030000000003000c00c441543c071000400003004c0730010030000f0045000103300000040cc0cc004f1001030000000ccc00c50000030005d000100400c00c17d4cf00013300000100040000011500040c0340c0700f00c003c0cc0300000010003ccf0c0004cf000000030700000305cc0003d004030000430d4300cf1000034531c0030c0010c0030304cc1c01c300000c0003f00004000c040400c00003cc0000033000000c40cf10050043000f3043033305000041440013000700070000000403010000cfc40000040f00310100000c04310c300040140d041001013000c300000000130000c0000ccc40100004c00c014000000cf70000400c004c00c00073130cc0c030c010010c4c0c030c430033440c040c030000010000000304130c0001c4c00000400337040400070010000000434000cf0c1313004010030dc4000c00040c0144c3000000000000000000000c0000030003c0c40d40c0034004c040c50c000010030004c0400010010000000003cc0f1404443cc430c1c00c00c100c0000c00007003000444f0030d3004000007c30000400000430000000003041c0d40c50000030dc30400000040000033d44f0100c0400000003c0040000000033500010000000000f4c0c0400cc11010030304004000cccf03300f0313040073c0c03031d1c5004001001700000400000010000001000300330c0304340000000c000300400c000141c1377304c000030500000c0533000000000140034c40000f30003305c0030000000050400c0001400c0c0c000443c005004004f103000000c3030001000d0c014cc00f0303c3c70040c01001103000c00030030014000040450041000010000040c40c0301c0010c00f3410130004040704000400044014c00004000c0400003470;
rom_uints[901] = 8192'h4c000c0003c0f03c030000cc0700c00100310c040001cc000040037401010401000044070c4700000c0304000404101401c34004d00043c0c000c01150000000001001000004c40c000000f3c04c0c04d4000c00040003d400400c0100770000000700014000c00f30500c001c100000c3050044004c00c000000104503d0004c0000f37005000c00400400100000004401d00c0003c40450cc04cc445030030c00cc00044ccc34000017000c474c0040c040cc000cc7010000c0400041400004500cc4d000040c1000000010c041105000f70000000c7415144000c030c00c0c003000704404000040004054147001f404c00d3043000000300003c000c000004c1cc00c4c70000c0013003c00000040000000c0c0c000000330d104c37014400030c0030040004000c0c004004440000cc400040340000c0000c004c00043030003030c07c1c104d0400f04f0c0004c3c100000d4700c0c04074044c01cf00000031004df10ccc000003c04500440c000c5c0c4010c00440c10000000441c30d1c000cc4000100003144c40134010044004105000003440c040300011000400004000000700047041001cf0304040c04004070cc00c00f4d01c3c000004100cf03104cfc0000000c0101003cc000440004c00c30040d1c0007c000c0c1ccd00000cfc30004005cc000c1400c100c001c400c4d03c44000c4000c004074000005c00000001ccc140300000d040c003c0c70700170000000c100747434c3004004007011300c00070000050c04310000004c1f000005f00411c4000100000c000143c300040c000c0100410000f0100d00000c00010050c0fc010130c4f43c10c17300040c01107c1c00c140000410700000c000004c440c300000044c0c44000000130c000000c013004001000403003000c040c0100f1c003c0c00433005c00cc0000000000f0410cc3100040000000c3000c300c01c0004000d0c0011030000f444400000cc00003c0000000c1330cc47c40040040f0007001c050c0004004400040101cc0c00000c40c0000440c40000000d0000000c01c0d00c700c00000d04440c1074c00404000000000cc00004c000000c0cd3300040000c340f0000c00c000c404c000400cc07330cc0100004410d3c30c300004c0d0303000c1c0c0430fc010cd0cc040040c040c400000c401ccc0dc001c0001040c30000cc01c0c4000c00100400007400000030000c0c0c0c4c000d30000c0cc000041c350d41340430cc4000000c73004000c00c0d00443d40000cc77000000004000441400000000053010000c0000c04c4030507330041110c0000c000c300c00000fc0f0000010cc3c0c30c4100c0c3c0cc0c00c00040430000010000000001000103003340d0400c000fc00c0c17003050000000c0c0404400100c000700000100000000;
rom_uints[902] = 8192'h4030000c30c10c1040440c0110000003f010003103cc03c003000017c1d7300d10f400fcc100010110700dc0f00013000030400303004d30130100034c073000101130c110c00c01000003070000040000030d00000045041330f0101f3f300100330040001010014cc47100f033303101c00431000007134c400130331000000d40700431c00000c0100103014100040300000004000c33033000303401010000050d0001400d10000000003300f00030c00c000070c3030110100c0003000f013031111001c00fd0c01000000d10c0010013500040000f003004000034c00400000001300010000f313fd50f00000003300dc3111000310000101000000030f000011401cd1301303001330400740000cc00307f03f000004c03300031130401001001130300000300000011040300c04331030d50000300000000300000010350000030000003300cc0330330010300d0003cc13c0d00c300740310050010c4733304c4dcc0077001051410030f300000004d100c0103000031403431014d100003113f03c3c003c43040000f00011001003f31001000100030000fc114d30c1000000d010100000000000c50300000c0cd0c301033f0d01100033303040cd00310001470c1cc1303440c00d0310c0034003004043003000040077010d7300c0c0d000f310340400034f0d71300c1301300fd3100d04001101c004000c000000333411701300000f01d110f000000400c1154d10f05100c10d003c000f3cc4d71001100c500300300300310103300011010100041040c3301500c4103010044000007000000c0c000073100043c34300300000011044310c1d331c0300c33fc011003c14305001170cf3000000013d300c303c01330111043000040010004c0000000000033c70101110d00010100c011c0101c0334c30c000003730010300100f0010f00101cc11100fd00000c010000300000300100033331133c00001f01c0c0c03000000010c0000000c00150c1c400040303001001041000000130310000c00000041300000c3010040000100034110330cd100000010071d30003300001c00331d433d341000400001010000d00c300310030000c410c451431000c00000000004300d0000c0010104100000040d00001000013cc411031d01010171010d0d1010013000c01004400133004100003000c3333300111000c0003c0f00000143000400100030003004000300d10105001130c000014c000030003c3c0334d0003000430151010303004101001c1000415010330015403301330101d1030c01c11030070430300011114004400004000100001000c00c000000100540000d4d10304433111004430000c10003004007300000004c0010030010040030c4000030c00001c304040000043371c00f011000300c44040105000344010000;
rom_uints[903] = 8192'hc3000000130300031c0030c00001044c010004c00100c0000c400c0c504c0040000d010005d0000000300400c000040c000001030ccd03c00c0003000004c0001c04d150c00c00000001c40000010043fc004c000000000f4014041000301000000100f000000000000c000004000000c3000d0300d0010cc00001c703c40001d4c5003000c00f030010000c0003001000100000000005030c14c33c00c004c100f0030110c4c0400010400d0c0304100c01000000000c51400104010f40cc00133000010000040001000c000000d3c0000d41000000001c0001003c00c303c0030100000040400c30000fcc4741030c0003000000c0010000c000000000040c0043c4044000003000c14301000300000cf01300cdcc00000c000c1c0d0c030000003003400000040c001c00400c000000000ccc0c30000cc41d410c010030040c000c0703000003400c00030001040c33c000cc004404f3c0000040445000000c0330000c000cc0000004100c0000c004004000c0001c4040004000040f40c000c0000c0010110000004c0007c1c4c4000c0400000c004000000010c100400fd04003000007000003000cccc040400c01150010c3c300100c00dc430c40400530000001000000000f0030c0300040c300000300005303f0cc040000c3c004c50030c0f04d40c3c034c00003cc400104cc040440c1c340cc000000030040010cc1000141c00c0c100000000c01c7cc0000010c103000000cd040414c4cc5400000c00440c1000340000100004001000c010dc00000001c001000c0c000003c004415000000000000440c000c00f4f00c4000000000000100000000030cc14c03304c003110c14d4000030004000400100004cc0000030c0c0003010c00400000000d00c040c000100c0c434c0000000c4fc730700c0cc0004400004110ccf703040103400540000c0000300c00000cc001c0400000c004400000c0d00c000c0150cc101000033c0c010c0000c140030cc04500100000010100000c00003000004000010f00300c0000c040000c000c30000c40c0001040000004c104300c0003000110043040040010014300c340004000000000300100010c00000100000003c003000c0504000300d00c000405140001c0c40003f00c04400101514d04100f00000000c4000403c1c00d00001000c00d00000ccdc40cc040c03004030fc10010000300d000000103010d40300f400000f0304cc4d0040003300000000c0070010700c000000000010100030f0c303c4c1330700c00000c0000000043400000400000010000000c0000070cd0000000055103000000c3000140000000000000c3143004000c30000100c30400100c0000c1000000000404c00c0403cc0c0000c000000c00304c0000dc304300007000000100440340df374f000500c00300c;
rom_uints[904] = 8192'hc0c000000c0000030500300000050710c300c414c0000440400c00004700404000000c44c100003004c00000d0000ccc0300c033c430040000300000000000c0004114c000c000400000c0c0000c10f010c000100040040c0340cc00c0103c40d000c0030000004030c140000c00000003101400d00010000c00530040c3c014400007300c0001004110c4c04010cfd0400000003003f3005070000004403000070000c00000c0c0000007403003000047c00000000000004000004310c040c00000000003400000c000130000013007c0004004000404000000c40033104100c00000004d300000f000c3014c41000300c00047c0000000040003c000000133007040004c11301000c010330000c0000740cc01040004000000c040300000000100001000000010c0014507030000c004d3c00000c000c00003c00400001cc3cc00c0003100001100d0f000004003cc440000d040ccd010c0ccd00000400001c000004010000c40c000400000c0000000040000c00000030c14001404400001011444c010c0c003001000034101000300c010004013044014000000000000304000400cc000000000c3c00cc00000cfd0300007c0001c0000100000c05130040000030010000040fc0000d400d030100000430001300110000000c0000000007f000403040c441411100003000030c10003040004d00100040000c514001000000f5050c00040c0030c44100004000000030057c10c3004035400034101c003100440000050d00000c540400000144000000000c300d00000c0c0c4400c40d0400040030c0010300003140004c001c0130070c00c4004000cc000c30301c0c440404043400000c04477c0040010400010c00000004004001143001c1010000400cc00000000f00050c300300440400cc300034030cc00000000000000c400004c4050000040000040c00004000010000000003000000004d1c300c0c400403040000000004000400003c03000c00000101030c00000c03cc0030c01130f04c0000400071014110403c0c001441003c0404c37033c1010400010000001c0c000000300cd004000dc00100c04430000001000003140c0004001300cc004000000400000c00100c000001000140c0030c00073f344d154c00000530000ccc00313004010041100000030100cc40340c0000500001073000313d00000101040c3c000000400c00043000000c00000dc00c040c00c10034003c300000303000c04d0cc0400000000c13400cc000c0340000000c0000c040000534010043d470c00c000c030000000000010011430000010005c015071000010000000000043030740013010000004404000040c4103000300000000000c000c00101000141000100000000010000040c04c4003011003100300101c0010014cc05c00f0c0000000;
rom_uints[905] = 8192'hc3f01030001330001130000000010040c300000000300710d0f03c000400301c004c0014300c0010400070401000000430000030000f00707030000c004030000000100014c00000000050003cc000330000050cc00c0030c0411440003c31c01c00103333000000100041100040110050cc0c0000003c70301f300c00d00003101000300034300130000000301000303000000c003000304040000c0000140304000000400114c0f0110c3030300004301c47000000000140030000403c400030003000000014300044003040007000100c0410004040000700100043c430d00dc01400101100001f0f00f0000000d0303c301000c0004004000400c0000001300040c0005300c30030003050000004000010000033303010000000c0400c0c000000000c00000c00000000c300fc003000300000001100000000403000001000003000003cf0003d00000070fc00003c7010033040033030303cc01400000114033000010010f01c00005c0000303d003170100030401c0cf3104040041c0c400c001030cc10703070000041003c00013000d000001000000010000c34043030331010103c00c000003030c0314c0000010140303040303300100000300cc01000000000004000110c1000730000003030003010043000301d4c00000c3c00303033000000001c41004c34000430005000300c004c3000100050103010000430000301103300330040000010000000c0000400000000000304301130033c140001000100000000000010300000000000003010003c407c34000c3c3c0037003c40441000101000001c0070c300303004003010cc40d010300f0c00001014000340001445c0003c00000070000000100000041000c4300c0c00140040010030400c300040000d10c0010c0000000010307c043000000000004000c000003011c34d100000013000c0103c0c0c30000c3c00031010101030000000000043000ccd0000000000c3300004000100000000001040303000340010403001300000301100c0043400003300007030000001040f0c04000000403000001001000010003c400c0000000c0500001000000433003154300000110010001c00003100001040c000043c00400000c0000030000100040007303c001000400c0100440334000c100001005004f01030c4101d0400400070000000cc0010003c0000000400010000103000c010100000000440403300300000000c300c100030000c00303010000c10300c000100044000007c000304000040000c004f0c100004044c141003300c0040040000001100303030104040000d1c50f00040000004400000f00030d04000040c0000100000000004cc003c0030400000400000003c00c030000000401000000c00000030c0c030000004003414100c013001cc0d0000c000000000;
rom_uints[906] = 8192'hd030000003000044cd0001c0130041100cc004c300304000000030003030c4400030001000000000001c34f3040010c3f0c0c000407001c100001000431003304c000000cc00030010000070f7004340000013450340001000c000c000700100000f431703cc30cc00c00c0c0c10001000000030000c0015007040010040700000000c0010c00004001000100000f10400000000004011004501000405030f0000000044c0405c4000000000003403474c04131000403000300c400411033103c10010030000033400100000c14000014040c04040c010c0001000c0f044440004000044040000030000003404c030303100300c005c0000000400440104000043c000c004c0c0300034c0cc404d1000000f01400c0c4030f1034004440103c007010f0000000000c0c0040303f040c0c0310000000041000031c00cc0c10c417c100400004000400011334c00000f0100d0340000f030fc0c00343030105c404000470001c0c000333000c0f004040000c04000c0434040411c3030000140035401c300003000411f45c00000043370c40000014000cf0330030c0d34000c4000104003f0c00470c04000000443300c34c043c1400330340071f000004000c031f0cf40c010040c000470031c000001340411003c04110000d3000030c04300000011430031030000c1010300f040030100f00c0c10000000340000004000f04c40c000004030c0fc0103540010000c00000045c040040000301003030f30401044c04c10000004000003c010404410100c040d00f300400003c004001001c000000d30c3300000c000007000c3000000c17c00413000000cc0300000c44030000000001d003011431103c01400c0f40000003cc00000000303000030c0cc30f410300c0000000000000c10014000c000300030c00400030030010010000400cc0100c03c3000c31c000040014000400000c30000107c40004003140041c0cc000000000000fc04c30c000300cc0050000343003c030c30044500c000340c0c4c00c04004000c0000400301004c00c33100d314c0000040c000c0000000cc0005030540dc404140c000300000f0301c50000c013c1004000c000140c73c0030037000001430007c4001c000c0340040cd0013cc00ccc03000c003403000134004000000d0400303000530001c40c0000000334154500010000350000040f04035f0c0d00000400cc4000170010040c040000f00c00d43cc4c01000000c4140000001c400c00ccc0cc303c50300000030f000010f01cc000cc00c50000010000000000331f003005000104510001000001c3401000000350c0400100350000000001470030003300000013cc031300300000030300011040300000cc0dc0334000040c030000001c40c4c04000000c0c41c000c04000c70cf04030cc04004000;
rom_uints[907] = 8192'hc00000c000000110c000c043030030003c100701cc4dc0404304000c3d4000000404d004c340300c7400000c0001c03100040101c0004d0300000c40400cc000050404000300000400000031001d0000010c01c30041347c4c004c001c43c000d3004004000030cc4011000c041c0401c04000004f0334100300100c340c0050c1440440000003304c0000c010c0403003000000c0004c10400000300404000c0100000001d0dcd04c004c05fc00073c011c0000003300004700c4f03c40cc00c5003c00001300030000c04c00030300d4030400c00300003500010301001c010000000030c0010c0000cd00d414303044300304070000000430f010400000300404000400f00d0d5000c0100c40400c00000c003f0300c1000035c0cc100c00100000c400004107d04cd00030c0c030cc37d000000c000000000c000c0303f00000000003c03070500c31300c004010000cc00cf4c0cf003ccdd000304dd0031f303030c3cc3000010310c0000c41000000043000c00000d10430033000005040333100f300031c0100000300ccc470000f000004500403000c0cc0c30034003010101c03c0c00000001c00100000000001cc0c00007340004c00000003000dc00030000700001ccc1000001c005c3040003004003400000c0000ddc0004c0000100c0000c000000c1040400000004c00113507503000d101000030c700c040000d0004c30f0030130c011050000c0037c3c40400000003c0770f0c1c00040d00f00044000340000313000000000000151000040c40100c0004001c0400f0310100000c0c0000cf130d44c00040c300100010033f30000cd1000cd000c1407d340000133010000403430000000000300040f0000c37030cc40300cc0030cc0007c03c0000401c0107004c4740c401d0c0413000c1100000c410c01c00c0400f000c400000c53003010ccd0fc0c3f00000030000003c4003003c00c3000000d107c0000000000500030000401404000c33000010033005c311301cc0113f30000003c000000030010300c3300030001f000c3d0c0730d000c00010007070000cc000cc7c000003d00004c0100000000004400000000100100d00cc0440003c434c3003700100cc400004c3c0004300044000c0000074001d00c00003dc40d047000c000c01050003014010c3c030030000000040c00300401f000000cc007000000004000000300000000030443c00034004430303017300440044040fc030d03c71000000004c3000003cf000c033c0003013c0000000170004c70003000404411dc00704031500000004c040001400031c300000000000000000c0c4041003000004004414c000d10000301000100040040010430c0300300100c030c0c00d0140c0700c000700340300130400300000000cfcf0510c7000004301000040;
rom_uints[908] = 8192'h4000c100001000000100003cd0004004030000000000400c0000d3300f330cf40000f00d110000c03040000c00001cd0c5000430330f7040310001000040c4100104d0d0003070001400c000040040c44000414044440300040011000300c14000cc0377500000147f30000f0000001044d0003103045333c00c00c014440300000c05000404003000f0004001f030dc100500000000100c0c000000cc41011c30c0004000000ccf00030040c0300010303c4d0000000430f00400400004c03010c100cc00000153503d0070040000001f04150004004030c0c410c4fd1c0000000c00000c0cc0400010000c40cf0c00000400c440000000000070001030001030c00c00d00c000c0c4000431c00000000c3c04010f050700c00003134330c7000400c00c0000000003330007000704700cc0050004c300000c0070073c1c0371000d0cc01005030cc03000540004004c01c004c4ccc00cc100000340000c50000c0010d34000d0513010013c0401013000fc70030030dc0c04300c01000100c4c310400c0d0003d0c0000c4000cc0104c0000000000401c00c00033000c4000000300014041500500f4104c4f0c000003000c33010000140c00300411031c000c0010c000d07000307c00004040004c10000010c0010f00000004030ccf430c0400440d340000010454c0001c70300c0c001044cc00c00f300dcf000330001330000cf01c0300cc00410d000400c03400010c40404000050c00c0c1440017410040300430440400000300440cc000040007700013c040400043730f104044f4143c01000045041000c34001000307c04001003000000300c0040041530c40000000000c7fc3003700000c1c0c00030c00401143000000000cc40040c031c300000300440cf40043534144017501cf000014c07000344734000c40d041013c000540c000040340000103cc0ccc41000000dc0000300030300000f00055310c4043004c140000000000000c4034104011300f010440c000cf004000000100d030400004013f00050000c0110004c1c03000c0700030100004cc010c0014000100400000000013c4005300c00f0c0300c03cc00100c4003001c00000c00cd000034cc000010000004c00004000c0000000400000070330033010100000f14010410030c1c0c000c31c0040040000000c30300c0000401ccc0cd0037000100030000c400c00c3c03000000030003000d1c00c043040001003c140430000101c4001140c0c0400000550f41000cc0c34000c000000f01040c0005004000c030300c057f0004040c4c0000040000403000c1c004c403340000441400300000444740f003105c000c0104cf0f30c00300040341d300d0000000c040c5504c1ccc40c0030300c0c000400300c00c000cc007300000000d01700403cd3dc01c001001043;
rom_uints[909] = 8192'h1000304000104c00000000313004000cc40000033100100004d500013c3000000c05044034100000000004040003004d1cd10030cd4000f00104003d100000300000003000030300000d00c01040000001000c0ff11c0d041401cc0c03001400005430343000133340000000300333400000033f1101010000d30c300c1c000d0704100001c00000000004001000430110500000040c07003000013103001404701700000003033304c3030c00c110000004001000000c1030000cc0300c0300c41400c0000401f0000000300004fc04001000c10c30540030000101131030403300030701c00400000004cc1c3000c1cd00010003100000100000001c1000c030003c3c000c3000031301c001000300c0c00c0c01110330350010401c030f70000c00004400331c10073000cc030000110400cc11000000110c000001c001011410000000100000100337000014100c1044f403000030dc000030c000c000000400001dc40370000301005000000d300c0100500300103010010c0101000304330d00c10c00111000010c007030c3d40000001000005400010000004005010301730000303000010030c0000701140c0000110c00d00d1100050000040030403c1c0f0c00c00003003330030031043011003104010034300300001330030004007c1400400f11000c00000005c0c40330110f3c0c01000f00300031d1073c1030103c000031c001000000001c100003151c0715001f17010001d10c010030030013003030c101000007011411000d0f03300030000003441010c000000010100013000d000c0000c00331000330300100c0033000c030010f03c00c0000700001000411d001030040000f34c40c000300040000011004100c400304003030000113c03cc0000331000030035000000111c10001343c0f0004303c003407c000031000c100041c00130400070704113300c0400c000030000c0430113413000010300000100041010014030000000440000110040001d0c00101f4000c0d1d1010000d14d04101000000004c0000000041004403000100010013c0003dd4301050331010710001003400343001f0307000d400003c30000300100310700043040d00000000001330331110030c0000003400103110f1003030003100003030000070030430000004c03d07030004000010343304000003cc0f301000041400c0000c10d440000104701300001001000033073dc01c000cc010000d0c0037100c003440340000000510300300100004030c4030013c430001000c0000c00c0c0010030000c10d140003000d00000005300034001010000000003110000030000c0c100000011100c0700000f10030000730c0000000000c000010030c013003c00030004000000d30511335000011f037301400300c04001cc000d3c00000000;
rom_uints[910] = 8192'h10040010104c00c040cc30d307003c040c301070041c51f440f43000c0c00300001c0443c0cc0040f00000444300c0400dc450103cfc00445000c00c00001040000003030c3044403c00001107000c4300d3003473c0310035d37f0040000f00004c40c30050c43000470c004344055000d0f0540c0440c0404c0c040f10c400143001c000f0040c3000000000001000f4fc1000000cc0c30c10c000000c00c000c10cc000c03c3040300000c4c044000130005c000400100000c0c000040040333000c04000cc40000000c00440f4c043c0c0000410c0c43000c0c000410040c41000000070004c007000d30011c10c041037c00050000400001030411030410314400054400001c00c404ccc330070001c40c000c30c40400f100100d5000c13c04f000041000000005cc0000000c00000030c30c0400010001130f04c00000140d0c040400c00c0c0030030440c000d000c701c0fc3430004c0040000f00c01000440103c30003ccff0cc041000000c0c007100001d00c03c101303040040fcc14001040c703000004000c300c001030043311000d0004111f4004c1cf000130001000c000cf4400040c00040d00f1000c000fd0440440000070000c04c0004d000000040004410fc0d40100010cc5004c00000c1c0043373c04000300c4300f0110000301cd5410003101c0500100330c01c0300c403000f3c00401310c104c0301004010300744400cfc10d07f040370c4000504000f3000000400057074cccf0000c00c007000040007ccc0400430c1000003000001c134000f00000003000000030c1c104c01000343000300300040c0c4c040000f00c0010cd00c30014c000305001000001f0c0c00400000c340110004030500000c0000c0000344c1440c0004400400140c44300d00004000cc015000000100c5003c00010c000005400000d4c4031740c30cc00cc00010000c0044c03000004034400300c0000c00cc0134000003c0030cc0000000c040d00000010c0d300005170033000c00304c0003430370c400004700400044533003047f1040000c0003cc000003004004c000010101c0034cc0000000010c100c00040370404c004500ccc00c010c00d00c0d00010c0000040005c140cc00100304000c1c000401400f1104040f030d0cd0004fc00c01001100000005c3000000030003c1c04130d7010300040403000004000c00c00010040f40c1400c400300000400010c30ccc14c0c40000000c0c341c00f03030001000f43c0050c0c10c401404004140c100001030d030cc0000000050000c0004c005ccd4100010c00c30000c0030004000000c0c1000c000f04c00f0004ccc31400004400040400000c01c40c100007000f004f71000004403043000400047040033001400000010c14040010c700004c1004041c04004c00300;
rom_uints[911] = 8192'h41000000d3cc40c00043cc3c000000005c030003300500004f41f4c00400f0000000040c4c000010c54d0000c00c434f0c00417745003c40400000010000430500c0434000010c00c000c034000c10000c0004c37f00335003000703c0c000301104ff4000000040cc0cf3000004c30001001ff0150005c00000000703c300000100f0030c000d4103000440400004c4440000000011007000c1410c440c40300f00c0054100c000400104004500033f100003c00c0c543003c300040043000c5d3003000100000000c04c0000000000014014000f400d504cc30c0043000d0101c0010c003500000cc0013705c00c04030c0301c0000000000c010303f0000000c00300ccdf0c0043040400004004003cc10c000f4401c33cc0c005c40c40000033c00d13050500000140000000c1c0017305000100300100f4040303000005053000c30133c30017c0c10c00c0df004040400440300c3c017130000013c50015c54170cc00c0c50140c300000100000330400c30c0010fd7f3f0000f43c0041ccc400140c0df00400140c1004f4000c0000340000300c3f0400404434300310100c304007001400040044014310103000341010fc47304000041000004100400440404035000400040c003730011000c000c00000fd110400014000004c00000c4010003000c400f50000f0343044040030341510043100000000540004341400d14c000000000c01dc0051300030f3140030003c70104cc4f03c0c5c00310c0c0000d10000050010c000c01040000c0040004d30010050000010000000f03103f00010010104400f00110045070400010000430d3c50c0440c0000100ccc150430504300000c00f0100700040c30043100000300000000c00300143000400c4f00007000000c040c0130341cc10400d010400000003300100c077000140c14c0000430140c0c310c17c104c104d0003004d04c3000004034c0fc040530fc470000011000001c100c00040040f400000000001070d75c374034440400440400000401040c30041003030cc03100c10f005f45100004303000000c14401d00000030403751cc404400000000c00c00d4c00013000dd030101c400013030340d100001154300000c33c0400003030000000314300c700040000c0ccf0000400101040050030004014140143000500300c3d1003c43c000c00030000340014c00c000c1007000d3003c00004033001c04000f030c031fc3cfc00000444f4c1410c1455050100ccc004004000010300dc43130030105c1000010103001030001c1700430c01f000f00030c33c7400005000f10000030000000010dc003ccd003001c0c4c03000f00400c01030143000304010100c40013000000000c4c0d4340104c00400c4d00004103c00c000003004344030000c3034c07010100004000000;
rom_uints[912] = 8192'h330500010300000000040c31030000030404003c0301cc0000304030010c0d100001404000cf0004f007004000000301400c0c0703c0c0070f0000050d00f04030045c0f00000003000000040c003c0c0c0101333c04c0730005004c30c5000000000cc075040040430c0000003d0003140c0000001c4c000040030f0001030015000000031c0003000c0000c40010304044000000000c340f0c00004c0400004c00000001000000000c00010403400c00310d0c003040c10000000c4400000400cc00000004000004000040c000fc0c150f000000430040004030010001300400c000130400040100000cc03013c104010c414044cc000c4004004000000010000040304313033c100003104c000730350d0003c031000301010014c00d014c301c0c000d400000000004d13100f000300000010400030004010300c0034f030530000400000f0005000004f000000301300000c143473001c007000c0003000100040004000000013000040c000000c0f0000040040c410100010000400000c1f05004440c110010c100000000011c00000100000000030c013000350c0f00054c007000000cd0000305c30cc33c140100c1000011045000014300000030341401010000000001c3000400100000c01004004c0401000000030704f000003d1000cf550c400c014c000c01000531001001103000173003010000004d000d0c000000400f0003004c0c000100c303c00c00000c0100000400004d300100000c0c0c000c001000400000040d40010c000f000f0d0000400001c0031430000001000c0c4c4400c400000c0330c013100005c40030000044000d050003dc000403000c00c545710000040030c000000000010c11000400004000000000c4304004003d1400001000054440334c13d41c0000cc104005030c00000000000000040001c54c31000d00000c0410700f0103000000001000000d000303004c04000000144c0000000000404000000000040003001f4001003c01400c000c31040000033f000035d0000040000c00c10001007000300154340c000d4000030007000000030400000400000100000000000dd000440000011f0010300430013d0501cc00c400003003330000000c0cc1040c010000c3c10f304f40000cc00c1000c01c01413001031010040004030000f4010000000001fc0003000014013000401105100303c1350000000cf7f1000101000300004000001c000070304000000333000f000403010000041140000c0f00c404143000000c00003300400000003001000c000000000c0000c00000004000010045c030c3c1dc00004c0c000d0000c01c0000000f03000403330000300c400d0304000c0c010011031c0300000011007000c300000001030040000c30010005010010130c10015c00310010010003000000;
rom_uints[913] = 8192'h30000004010c00040d4000070300150c3000fc03040700000c0701034d400000000037010c0000011100040300040311001000000c01cdc10004011d000301000103cd0000001700000000c00300000100c10cf100011010c0c4030001300003033000300401000001130c3d000f0301030d0400c3001001040400110c0c40c3034300111c000000c0c01c000033000000030000000c0c000030000005041300000000040701c000030700003100300103000000110140000103110c0101050000000001303f4cc30300000c0000030000110d00c13c00000f001c000f00000c04000004010500010300310303c40c0501034f01300000010f000000000030300301000000c303110c0c1f100000000703030000c5000010040010004303300010c300040300010301000c000001030401300004000100000333300c03070f0701030c303010000d4c03070000010c100000000303000333003310000400d3010011000c001300000c010c0400101c0c100c000dc30000000003030c110c010f03cd000500000000400000c043c7100100003c04000c000000010001001100050f07100c4510010c0c0011000000000f00100105100c00c00d1000001f040004000500070001013140030300000005004301035d103f0305000703100001040c40010003400004003303000c100c00040003110300000c00150c0001001503010100010000030c03c103010001c40000040004c0050011301130f40000031100f00f000cc00000000000030100040004000c00c0000300030d31010c000103010000004000000c43030100013f0c030103050003000c0c000f000c130341c3010400070d030043010c300000001001005c071000014300000c0f050300030000300000000001131d03010d0004301401f10105c3110000000003000401010c00440000030011010030001100010307010300300c0300030c010303000400011000010001000004030100c4030013040303000300030500731000330500000d1c000101310003030001013003030307440cc0050000000001000003100f0504000040031f000c0001001010000c00040d0000040fcc10000301030000c00000010d0004341c3c00013001040003030040003c30104700051040000f011d10000303c0000307050007000c0030000000000c00300d0000c000070d0000030001040c03300343001103011001070000070700400001300107001340000100310004041303000003c010010130c0000000400f000f0407000f01030001010c000000000000cc0c011c00000400c300000300c0000330000004000f04000000100c000000340410430000040403000f010c0000070100000c00000c110300030f00110c01113c01000000000000000c0d00030f010000031d030001033d10000f00;
rom_uints[914] = 8192'h300010303000f030401013d100000000d0001001001043404c030c07c0703000004044d0cc0000300400401f000d01333c011100c00c001300030c0000000000303441001cc011030000fd74000130d40100044430011d5c0c404000c00050114301d70c01000770cc000000300001300030f7303d704000000043144314400400c3000040001c403000d0004000404043000000000010c1770000303000c300cc07000011f10c000001c000000003c300000000c30030c04000344040003c001f3470000170000300c043731c10000300100140404300303110dc5100c00310001005040000c000f010c4f4c1700c073130103014000040004000430000c0130000300110100001d0c0301003100000300000010f341030710041f000c0c10001000030000000c100100300c07011400100001103c00001004030000040301303014011500000000000c0000040407053f300d0501cc10101c00400c0030000f0d1f10053c04c0400cc437c00d1f1013040f00c310010000300f000010010d1f34030301100030c00401303003cc000100300f000410040400000030000400c04c010c403010d400000c3c0c0441000100001d30100400104111371d14050dc0040c0500000033fc00000c1c4c30000001040c3141310c0c30330c00000c01310000c4004c0c0337400504c3000c00100f0c100c00fc0c33c0000f0000000000400470000030300d0c0c0130000d4004000000000c30c130070400140c1c30000110030404131000014004c00c400000031000000704100300001f000037000410010f000c1c03011404313410000c40500001033c04013c10000c000003c00110003334030300053500110007100300001c301004040cf11030070730030005000c3100cf0300043000000d0403031d1003031c0370000404000043040c07000301100f0301f1013043010130040100010000031f0010030c0000000d00cc143c0000000100000c30c40ccf000000f01403c0300400000c430303030540030004000d30300401000f00300031103107070c30300403313003004d0000c0000c1400041300c000400400300301010100300d00343c0443045000c00010000434000003000010003400000c00003100031d31070104100c000c10403c7c1c0700000400000300100c0c3031cc00f004173c00004504c3330c3000005f04310c130300301c0c0004c1000c040001040013031014303410000400003010df34000c01c01100003f04cc0c30d000040c34000c1403343c03070004003c430330004c0c3001c0074000003c050100100130050c130500033f0000c00001044f0410050d000c071444000c0cc04c0001000003041c004f000d0c010047c00c04030301c0000c31ccc434010400030403010100cd001c170013070f0010030000000;
rom_uints[915] = 8192'h4c3000c0cc0d0c101500c001d004415c040c0c01c0740c00057700040434000000000c0c140c00cc0050310000430030304c000433041030040004071c1d0007c40000f034000040000c000c0011cf3010001c04d0100cc030c040c304030fc0ccf00c000c0c130c140300003443c000100c00300c70100c0c7410f40100400c054014001401044000c1010340100cdd4f0040000000c0c0300031043300100cc4c0d31c1014c0d041304c1434703340c40ddc00041030010c1000f4f5303003337000c0f00014c00fd001500005ccc434c0c400001000334730000033c001000000040534730001cf70043cdfd0c4cf43430c33c003070c004044010000100030000003300c0374043f00341071030400c00130000d053c00c4041043340fc31400000105100c334001c3ff0c07dc0c171000004004003443c43c04c3300c34131c34c03000c0014c0040130044c100d4c0003107c0f374c4770c3cc40301100014005370341c040cc303300f70000040044143030704030c034030c1043105d010c400c4004c43000000c03010c00030030d05000c4c33dc10d0007000d4440c3043d500ccc10030544c1c3044c47c703000cf1c307c7c403105740001dc004003d311101c040104001c0000000014403c007041050034030c1f03001300c0000c1c0c043000401d4c3c30005003100cc4f4444100430404f0000c10070f340c00cf10001f30300004000dc0130c1c4030001c40c31001f0407cc4001f3000cc0000000f0000300045f00030c40c10c1df000c04ccc1c00c30043c44030035744f00007c000000c437cc3001d0440c300f040013c030003730f00171c4c370cc40710c45000343cc1003400005f00c30c04d00f0100001d40010d13440301c3004004403000c00400c04034014000700700c14040c070000d0000cd0f501044000c00030040473470c7041141c004f1c04304005c3101514477c33cc30cc75717300c04000fc100c0001030c0000d0c534410000c344303c07300001c0304c3005c00574000f10c3003f101c0700c0c00c001f0c000000005000000c10cc100000700c1f303474c0000410000431d1cc00300cd0000000170000000f00c4c034300c1000304004301c31140cc4300030103010040404c00100400c1cfd4315130d114100c004444330000d10340030033001004300104030c7404444503104c000141503001c0cc704013010053000100403003045034fc34030044dc47cc3101310000003c000c030d44003100004000110c01c1c300c0030000001003400343c0300003305050c0400c310ccdc0005050003400c030c0400c00005fc10100d301c00000c0cd0c0030c044cd5300003c11000007c0fc4353c30c70c00054cd400c0307c300c040c40f44050000044001034040041dc04444cdc04000070d;
rom_uints[916] = 8192'h30000000004c0001d0000000340000d44100400cc0c0f1c000044000c003000000730c0f1700c0000104000c000000d073030000343c00044040c0c030c004000001f3c3004000430c0000403430411031010001c0500c7301c00f04000040000000c03504000104404110c444c040010404403c01c100c00000334143c0000004d1300cc040044300000034040040000000004300005000c0000000000700000044cc44c4004453c000c3300703000700cff40000014003040000000c4110400400000300000c4140c30000000410044134740043c4003107d000c000010000cd0400003c10030000000070003c0504c045500c40000000000010100140000c3000c000c010c0f0344000c10300030fd155007000307c30c100001f300c10c0000043001040000100031043c3004d00033040c000000000400301004000000d0d44014cc14040004034004040010c0004f0030d0003704704c00c310003cc03007000101300c47000c50f7040c0103000c4c0055045400003303000054430000c00534001400040ccc04400c40007c40c0000000300710000f110003031404000c00300c0f0000000400c0030403740001044513401c1431430440004c103f3104040c03004001003040c00040030030401c00147cc33f004c004003003405000003111c000c0040140300430c10c0c04100000f010004300011000051c00340000c00d00310000000713c03070040004000300cc000300005140071f310004000dd3c00003001000000300100003100cfcc100300334c130404003c1c0c07001000003004000f0070f0344004400040000c01c0f0c0d0f1100000000004000c4000000cd01000147000000400000100001000000330000504c0000c140000c000001000043c40c040044c00041c000000030430040c00300430000000c0c0c0501000c300040150341004400010047c407f0400f0104c0c407c74007003c010f30040300000001030003400000053400317003c4304003303100cf040c73000300300c44c100c400000004400010030c030c0000c3000100000000d003c0104400d001c000003f0400c000001d0030000104c00c000000c040c003310400004d030000031040c040cf00010000cc00d000300f7000c000c440100c4033c31050dcc310f005000004000001ccc00000000000c311010ccc0c040c0c5043303c0000ff110000401f03000003c0004400300cc34c50033000404000000400400013d704400c00003007040c10040040000340000000d0f0004100c04304d000004430c0003004400503010040430000000033cf00fc00301501001c00d04041000000007500700300c0c10c0c0cc033ccf000070300c030c30004013cd1000403034000004405000f14040010440000c04300c0130004040d13c0c10440030110;
rom_uints[917] = 8192'h1000040040dc000034400104030000000c1c00070040010014400c00d41dc03011c305fd07100044c03000c0104c10cc0350c015001004140400100033040f0044000c10004000141c00c1014c0070c3347440d1100fc31c4303f04c0000c40510c0000000c03c4010140c000400310010c010f0d00000fc403000d5040c101c0000cd7341030300c0110040300000043400000c00401c400c0100f00001c41c54000104c00c0c00401300004015000470c041d0000040c5040101d0513000000110cc4034000051030000404015130740100400c104000010d00403100fc04300400044050405001040d041f1d07c4fc0c0030000c1000c0f00001310000000400014cdc000c03000000cdc04c000c050cf10440c77c110334300100031040004100000dc00000cd0400010c0d0043340000cc1c0134000c4d0c40c4c34d410c000005000d0074030c004d00cc04c11f0543c1040cc0400c0c013c00f11c00c703cff000000c100001450c0c01007140030000c43030014c1ccc4f000005d005c40130003d00030000000c0101077d0070000110c00f311030000004144c000c054f13c00cc100000f03c100015040300f04170000300f3030d4310404c0003c440c001c000003c004730000701c4c733000103030c3400c70000c00434007f1055c04000c104cc70c3d0070370304004004c0000530011050400000c0000070040130c00c7d0c411f540304130003c0004f74004004030c400333c041007040d43103113010000001c1400c00001f0300dc30010031c00401000404000cdf30003f0041d4c10c40000400010d040cc004403354d40c1073cd4c040cd00001400c0d000f000003033d010c41410000140000f00044d1403c01f0c00c430c01c00313000f4100030003c0c00300d1c100040101c0040c00300d000013300400c4300451001c00cd7d0101004c44013c3100000c3011000c01c044314414000004140054340001003c004100400cc0043c00000cc00004001c04403d03c4cc3300000143105d0cc43000400c100cf000000cc0c000000d30000000000cfc00003000300040010d03d3100c0000440000000000000030000014311000000c05000400000040d3400004000040440cc0c40004c00000cc01000443cc050004013f04fc3000c10c003d343141c100c0100000454c04104df00041cc44000044c04011000f10010500000173000303c500c04400c540f00f000303003001000070341ccf1cc004000040f4f00c4007f400c4000000000c0000000d3c0d704004000c10c00000c5700004030c0710cd0040704000041c0c000400000000400001c000300c3403c0c53d00010f000c0ccc0000401c300f001c10000cc3cc010d71c44343000fd000c0000f00000010013033000010c01c0000043f0007c005140000000;
rom_uints[918] = 8192'h350000000c011103003304300f101c1005000001000000c300000f0000371c00000c04fc140f0003304100000000010100c01c140003105c033000703c000c300410150113040005010004030300133300000010500000141f001c1c00c400301013000430300003340cc70000c10401010c11c0c10f001d004100003c000303030030110503001000000331000c101303100000000310010110300c4f0100300300010403305030110c0000cc0300c4013004070001500d33000001300c1100141304000100000301010c000010031c0000d70400c15000010f00000c333c000c000030000f140f000004710034010303001c0c30040000000430004330000c403d0100054c3030004000c301cc000000101040301c3003ff3c01501513003cc03004001003010100301003c300030004000c01000311001c000400330030030f14000001013c000c0700000004c004013500c000cc040f5d0d0f0c300d301030373c00030c001000030034c0000f310c010c00c040c00317040d3c0004100040011303001f105331043000fc300c1c040003000c00000c03c0000300301300010503c0303510000003001030041701101f33100300301300135f10010c300000040034500010000400c0000c0001010103510c30004d3100001100c0110d04c304000714130430035c1043013301310d00000f0003000030000000001c3cfc300300c0c010003000503d3000c404003017004030000d000010003f0c00ff0c3013510100040010000000330c13000000f030001c1010000000000031003010000d010303014d00100130040041000030000c00001303000c31000000430000000001300f0030000001700c04000c0300100c0c0c031005000004000fc10300001c00000c10000330cf033015003d00100f4004000305c03001000734003010004130010f00c00c04000330130d1700000c311010003301000030000000300000001010000000000c000034003c0d31041c0cd030001000004000f0013703000300400400000c000000001c04010000003c3004003410003c0003000c0c7100400110007304004300000cc10303c300470300030011003100030030000c00000100001101c3001033010003000c11003000c014000c30000004001713000103000c300f005d003c0c000007d0000030033000f701c50cf1304300001c03c310010c000100030000030f1003000c030000070701005000010010001031c001105100445c0000030d4f00001c1c00f30004370000000010000000010000000034000003033d0c030000000000c4030303000c001f31000430000014000c1c0330105c0033000031c00433010100340400050cc00000000000033c33330c0f300100010031001000d40003340c0130300000000003001040300c010c0010000000;
rom_uints[919] = 8192'hc00c40000100c01070c3007445c0000c0303c14fc013430100d30103c14331000040c00507c30000000000010404ff0fc0407000000007770cc0cd000344030440c331f3000c00c0010000c1330001c0440300c043000fcc034001000015f000c1010107404040030040c5000c0341000fc0c005c000c0ccc00100c0344000014105c0400003c3cc00c0c0c0130143000000000000030047c0450000c30c410100470c0300003c403c04d0443cc1c0c0004104010040030104c301c10c0340c004c0000040000101100003d330030303000000040001410303c30143030cc0000100000040000040001c00300001000100c4cf440310003401000003010000034304040030011400000031c101000000430340c1000300074040c0000041c04300c10000000000c3000030000700c3c00f4c0050c0444300030100000000c100000cd50ccc030001c304134f100301000c404f30c03543c04fc4300000cdccc74c00c310c3004c0c35473001000410000000f0c040cc0c40007031000100c100d34cc0c000c1000c00c0c000f00143c4400313c34000c1c040400700104001c0c00c4d014053c0000003000001d40000400005c303c300100000c00030005000040000cc01c0003f040cc50343000000c30500030050c143c0000001010303cc0040010d0301040743c0000303000c40030000140175d000030000000405007000010f0005034000400c010041030010c30000c10001030c040001c0040c000100f0c0513c00000004c03500c00010c0000c004c03c0ccc007c00c0170010c300303c04400000001050003c4030440c00c01c3011043c1000000c311dd403001030511014d0001034c0000030000010400f101050100c0030000400000c1050304cc00c003300405c4d10003100004303c034c03314f00440c0c0000340f0405cc0c0100404c4c03000000cfd40c00c34714c0004040400001000000001040000101c00300000c00c3000001000101430005014c11000f00410003030310c000c1000001c7c00cc3c000040c1040c35cd003011c74000100004c0d05d004400cc700c4c00341001005000100004000000340000000000511c0310103000c000140c40040c0c40f110104310300c10d000000031ccf40414341040000c04007000003070040c000c000040000400300000703400400c0000003c00001004c00000300404c033000010103140fcd00c343d300c441000c451503c30001c0030f013000c00f03033054c3000300c300100040c703030101c003010c030304404400d0050000c40000000400000d040101710cf000c7c300400c0300410001c0000000c4014c00337d0500000f403001000d40000400010c0050000000430700000040030000d300c0300000010300c40c03cd00000000010040000c400fc300c000;
rom_uints[920] = 8192'h30040040000400003000000050c034c0300030103000304000cd4000043055c000d4c0341300404040100c0000c04c0004400000300410d04c0100001c0000000c000030044030c000000cf0cc001000001134003300c00cd030004000c000000001c3040000cd00c0010000000f05c000000004004d000cfc0c00c000f00000000c100cc01d0000c0000003cc0010010100000000000410330401cc700013007000c0c00400fc30c0c00000003c000c00f043c0003300c430c0c003cc041000c01c0340000110000000001400c04c033007d100c043444000d000040cf000fc41c0004c3000001030000000344f003c01014000000000100c10000f3000000003400300400c00030010c03000000040000141c4c040c4314030c0004004c3c010010000010001c000300fc0000000005000c004c010000000300001c00000c0000000c00cc03000d0f1044c00c070000cc0000cc500004004c0ccc00000000030000011cc000000f00c330040f00014100000cc00ccc000c0c704400300c0004d004500434c00400000c00043004cf0c00000000000c400c0001000c0404c000300c003000300100010040000c000000040401c0000040010c400301c000c0000041000000000100cc407000503c400010300000000144000000000004c30000000000c000000f000403c11300000400040003000301000304c400000c000400040000c00f040434140000c143c0000003340000500701000411c5034c073540300030c00c0000303003c00f30000000000c000044000c00430473040000c10c140404000000000400c0000c000003014d0033c00503c0000c030f000000400000030000000010c00f0ccd1c000004c0000010c0000003000040000000000c0400310300030c004c03c030f03c10000d0070000007c000000000100c300f003c1f0001003001000c00000c0ccd3000010ccc400000000010000003cc4400050000040000000c0000001c034000001030000305005431d0033010c0000030110d000c040c003001000030000c000d00c0000040c00000000701000f000000100fc4000000000010300000010400d001043000000300001004c00400000000001030c005003030104c00001000070000041c0001000400000050000cc404410040040005070004000000010030f030c000040c00c04f00c1c10340c000d3040000000000000030030100001400c000c4000c00c0400c03c00003000c00000030030000010c00000044c0cc01cc0000c0cc0c3000045030c0033040040007c0070c03c0030000304300000c00103400f4500303c0030004c1004000000400035040000004c0000304f40000c0300ff000000000000040c00f04000c400000040000c301030c010300c0000000001000000c1400000c011c00300cc10300c000000;
rom_uints[921] = 8192'h10003000007cd0010050000ccc00030007400c0c0cd0000000c40000007430c03034c1001d130c000c4410001500100073700f0cf304105140c00070000104000110100d000000400000d0d01000d001400c00714c001001000c00f40010001040fc040dc0401400000c3c030530c0410003007c001100c30004400045040401c3014000dc310100004c003004001300c413070000300400001030303040001040130004000000310430140000070014003ccc0100000010d30000100d001030304000304000d000000f00047030411454030c70004c1330070004f3034400003f130010700300000c040017001c070000040d0000000011000004c001100000730c40700c100d00001040cc10010070300300144010100c0d13000f1000044c00004000ff0c000010031c00010000c000031400040000301000000070c0300014fd100d4030100037101001000100003340c004400c30044f133cc0000704040000140030c031040003000c00101050004044400cc0003003000fc00000040c50c0700f00000430440c0000140c051733000000c300c00c4f000130001000040c1c0030c341100400304000003300070003300500c10c041000c10700c01000dc75300000031401000000001c00c300c40000000313d030000c00403cc0100d0c410c01000001400004c000c03000000d00045004030003000c0000050c400f30000c1c1403c00c0df310010f00001414030000030110070c000000d030103c0c1c010040d30010000000040ccc0c01710c11000404c0100014300353005300040003004cc00000c00000c3001c440300c1100044410000310f000004cf00c010001000170c300100c01354000010100dc0100000001010f330000c0c00fc7000140000040c50c04413044010007000c0f447430430104000003330140010000414000030033c00047010001100c01440c30000000300001350300c000000041400031010001c3003000c13030f0f330c3004033440040003c133740510044407000c001c40000010c015300501003c0430003d001000000330030330303f0434030030300c3133c0000c000030004030cc050000300000040c37374f44030c0004001c100400010050d00c413c3300000005d40370300cc30000103f4000000100c000001400101000301fc7c100001c400013004403c400310000103c00001000f04c4030300004040c001030700041404f4c0000700100d10000100004c000d00dc03000030001030c05030000cd0011c03c3010d0c000001c031430000cc40001c40300043cc00000c100cc10cf04337000000000dc00000c004003f00000004073003c030d4000003c010c00000040100000c0000300c0413000303cf40d3c1100000403031017400030000000040c0f0000010c4573741c503010c000;
rom_uints[922] = 8192'h400700340143000300f100c10000300d03014c0c700510004c300053c00c0100000000400c000d00031110004041c040df0c00005cc741c31004c03d0001405300cc0d10400304000001c071000000c004d04713300011310114710070137000074c144100340040300c313000000c000300100443010100403c00003400100c03c130041000c00003000503430030003004100001404d041030000cdf30000033cc0c400411030c00400513c00c400000050000c00cc0030c000133000000430c03013000540100113040343400711c044dc3103010100c4f1101f0cc414410171000d100300300000c450f44c0c0c000033100000041004003700000100001013000c1c10031300d000305103000003003101030433030c401000000100031000100000070c03cff104c100053301010010cf000130030040c100c0cc0f003004100c0f0401000000033000000c034000000133030000300001c4030c0333010410033400c00cc0400c1430040730000500001000000c03511005d1c3040413f0033043503101405407031000105dc0000cc0300c04d0331400030000c043f00c0000c040004000301100303c1003d000340c04011044040c1001000c0001700300301000000003010011110c030701030110030550500000000043131303001004400d303c303c311000110004011101d4c0000700010000d00303f413134140130000000f300401010c3f3000030040f101c00410040d331c0c00340040000700c1133c1d7400000000000c75330c4cf0030050040000d0005300030001cf5d3370001c010150130110c0c0f00000430000030033014030000100000030030000300040004c0000137c40001c0cc40140001c00c40130000103313330150010300100c00c300003d10c700100051dc000000f100c00000c0000d00000173c100100037d33f03040c0c3431103001300000c0c030c03010010153003001030000300000300141000003300f007531047100033103013d03303c010c0041030003075100311400004004000c3c0014000f0500003300013000d0303c03007000001000100033d000004c10300340000033000300031030c30000110f304000f00000c04f3004c330c00010c53c00f0dccc45000000000070000f03d03503030000000000c40c70400d40070031c4100004f0030000c410100030401040c001c0d003040c00c004d00303c400043100c3300d30001d001101000300014130040007410000c3d03430004000f004340703704010c3300000010c003000c3c0100010303cc00f00001000103000301340cdc073000010000000310003ccd31100310041c10114030003030140c1301c0000040c10000003d000000300303100f03040c04c00f04f0400c33000131c00013010010c1010d000f0300000c00000;
rom_uints[923] = 8192'h5001040cd030400d0304004c10540c10f400040c001c03044d0f001000000400d330030c3f0004133c00010c00004403000434301f3004c0040c0c013c0d00403504c3000c400f000000f170005f004c33d401340c040d1c004000000000030510040c00001c000434cf3403c50cf10d4300304c4000d50cf43c3034dc0c143d30c10401400003003400107c40000f0c0c50c0000030c030c13001f411000c04c0d400000000c4c400041c34c01030400c0d0000010105fc0010331451043140cf0c3f043401c04c04000000cc44400403010304300c017c333c30f0d31040f0000030c0c30504000000fc0100130401c540003c0010000d10030040c000030034330f0404031f003c305f07100dd30043054c3ff41c34cf4c34c4001310c0001300007d0010000cc0c0c0010000c3000c00100000000c300c001303004300010030030004c000c1004030fc041c030040c01f50043700000771040cd0fc004000500c0010100d0c0cf01757c003000000f10c4c0c03c4fc13f400c0014c031c01c00c30030000c40c0300c10037300400330c0000ccc03040000c1c00000cc4003c0030430c000404c44c3d330433000000003ccc00c101000d300500073c3c300400303000043cf45310000cc10045f0001010001d44001101040f00c45400300c3c10073f00407c5c1cc01c13c4401000c00c3c0014c403000003f40003401c00c04c04440704f11c0400d0f00f0c03c304dc4004511c40543304003100f00005010000000000000314c400303f37c00d140c000400104103303c0000c03104f104300d004c14031001fcf40c31100400000044300007f0f040530c4500103c000310030c050c301cff50000cfc0401500003000100d4d30c00043030040d073000033030000c0c40040001c700040054c0541c1d0104011f00fcc0f30c1510500c04414f003c501f4070000c0c0c0ff00404040441403000c30c01007c13013003000013000174c0000c3f003c40301cd01cc0cc30c310d010001f00300c007000c1104540c0f00000441004140c34d05d01030150040000030330300014303003005011d5330030d40c0c0330343d041004003100343cc0cc3007330040c1044430f0c05400040f0c0000c00000000c400c00000c114300043c50430c5430c00015040c0c0000c30c110000001404073010c400001004cd04005414050cc100d0540400f031030104000403003c00c403030310051c0c0033c0070c30f7303011c0303d1000000cc40010534c4c000404000c3010c00000000c0c04030133401cc307404dcc0101000100001300000000f0000c00000c050000000d100000004cf0000ff005c31404c40030030113001410541000043d3004440000333000003c4c30c0c1043cc3300cc0df000003000300410f0034d004c410110000;
rom_uints[924] = 8192'hf4404100030013c0004001000100035003c4001103c010000000c00000c5c00000040cc307f34000334107070740330cf4c01c040d30005710d00c01cc14300c0c004f000000041400000444c300c04310130003c00030401c01110c7cc40c0300cd07070030100003000f000043030347004043300010f00c4f31007073d0c31040340c54c00040c07d0010000010d1d0001000004dc000f0c3300c00040374113100040100100404dcf0110000c003003d53000007000304000033c0000400130c337c341043000051c340001c45033040103040ccc35750300010030030000444000004f34700004c00c574334001c004d30c1c41000070040100c10000000d000c0001d0300104103030cc1401d101f000150101c0c4c0c0f00cc0d000cd000f0100f001003000c0073007004000000d3c000cd030cdc0c3010030c05000c41307c01000c00c3cc000100000300000303001f5c0c4c400c43114030f4c4040350c0073c3c40030100301c13017001c340f031c00c0d0003007030000cc00f00000c0cf0cf000441f30c050004173c4004103300137000c0000100001c03f70030130000003031c00050c4010c0fc030344d000104000010003c04103030014040005d0000700000c0001c4f0470413040300c04055c000c1400010c1003130050c0411f01030013ccc00007f00000444c0c700d0c00c30c01cc00cc04100104c000c40500f00104c10c410f344030003c100c00041101c00ccdcd01c47100030f70000370c03403303003344c10000304400001cc7330004d00000003000c0cf0300000413101330c0510cf451340000000001c100d0c10d000347d030dc50cf0000030c1f0431c000f1400044003043c000c0100cc001004101c003cc0153c4100c0c00304740f30030c003f73c000d41c00101007331c01c00300d033374c341c0000000103c3dc40513001c30c0c0c10d030031000340c0c00000000003000004030000000fc300c370375070400001400431007c031400c04030d0034000000111104d01004007100001300dc04d0c401030d30030000c07f73c110c0430300301c340011100000100c000c100030040310c53000c00000c04700c00131000100430dcd00033d31cf0f00f3cdf07c1d0cc0c30c004c03403c0c00300d1f301430003cd00c0c7ccc003030030400d30330f400c1c700450071000c000103300003d0300c034100710c0003153c1000030300c0c5441000000701331d0c001044c0f00d405f103001c3c0d01031c04dc413010c33033d0030103f0000cc007003004000010000430100000d4dc00c004700700500000c00000000003010013301d330d3004000041000000d40c0401cc00000010700003c03040031c000147f7307404400f00c000104c070c001010c0c001004040cf31000440001000;
rom_uints[925] = 8192'h10300003003cc04004c0000000300003000f003003003030000000300c0c04001030003c33003405400400f4000130100f0c0c000001d010300400530c00300010f03c0001c00300003300c00130d4d01ff4003cc41c303004330400400010371c03004000030000c00f0cc0d070000500cc0c01c50cc00307000013103000c430053014300044000c003304000705000400000000000c00000000031f1030000c41010034c3103c3000103c43103c003030000000010f1331030f0f0003010313303c7000007d30000030c004f0310040010cc04004c404004c03103500170000003100f1d430000c003f00c000c00c00c1c0003404c0100000001000000000c00c0c1030710c4040c004000004013300050403c700310f0030041c1330c001030300010c100703100110000011030303300000301000000400000c0300fcc400400001000f0401000045f4d31300170c35000cc43c33d100303c033c11c4343003013cf41037031005500030331f0013100111c40c30300cc7001c00cc400c00000000c00130100f30c0343313303030030000003000030000001c0413100c0c30000000c00d00403c03cc04c300df000300103000040cf0301c0330d05f10000c717000003001000000000c14014004100c0014f300104100000000d03000f01f0104f40010431400001c13075034000f000f003001000004001c33031fdc0c300f0f300404000100300101040c040440000114d5010340f0c1c43cc001140c0c00303c0c0000c00c3c41033c10000d3300cc0ffc3000333040130000040010014000000400003f1c001c40003000040300c13001003310000430030000c030403000001304100100103400c43430130410003003000130040004503143000033c0000003000010c33004003c000ff1300c301303d400040c0044000c00733434011c033c0300300307300000030003330014300471001370df000301c0c000053400000000370400000c1f0030003c3043470000ccdc00030430f33407010000403033100004030000010fc0403000d070000030000010100000030010d00010000c30c0400300034004cc330d31500400010d040000d03c1004400003100300043010100430110003300c01c000103c0410dcc30330044300400c400030c000300430003300005d010030400030c30044c4f40014030c000000301c00000004400033000031010004f40010003c00000c00c0c3040300003040401405c0407d3cc01010303007103030c00404030030303000c00c7c304f30c4000000430f0f0000030c0300c00070cc300000300c300000001300f0340000c133000c4c400050004c033d0013700c403c401001000000000100300033000014000034400004003001001000c00103104c100003000004003003040110403013340030;
rom_uints[926] = 8192'h4000c00c11c3303c3040000000c301000704040c00000010400500c4c004034001045c100000004440f41000044001d1c40010c30c00df0000cf0c7040c00000475c0c00dc04000300103c340cc0cc7300403303310000c3000103c00d00c000df000304113400000fd300000c7c1100010343401030330001400c40410ccc0000dc0440040001c00000100d000005013100c00000000400000c00c70011c11000004400c0fc030d000100c0c1c3cc400d53100000cc7070000100000000003dccdc00000140000344037443cd130400c30c300004c30f0cdd01040010041100000cc4cd000004000003f003003000c401d4c300c000000cd1c100000500143700000003031000d0010c10140700111073d07c0034c0c3443500003033c001041f4100037101c10140c00f03004c01003030300007000005c0c000330111000013c10010d40040000d0000401000307330c001000300d10cf1c0473301000c0003040d000740400000000101cc0d1c00300050000000003040000134000017477c0331d400043400f03000110d04000000c000000001c0004003434041f30001cf0d1c4c03c0310041010000c004f007c040c40004d00111300300043330034cc14300f0700c0170300000440001040cc44301cc3d70073300404000050030000003c700c1c400070fccf1343074040cc0f40010c334413cdc1003c001c1470000040001701401d34000440c0000c0cc050140310c400030c0c0400110cc470c0cc331400000c0031c40004fc0c00c040301407000030c001111340000c15000c04043100c0300170500003f0301c000f00c0d45040303c000100ccd0033433000cc0131133003307300c0c0000cc1044045033004000000300141000d1001c4c100f03003c070010137003130374334c51d0010030000100071007d00c30cfcf10f0000303005c003d00c00001037003d3000000c04000c0104000c33434401c3140000000c0703c7c003003c00105c10c500000304c3c014c0c103c0c0004d00c034f10340010041c03475400c000c000c03100d0300030004ccf10043000407000005c30cd1c0c000140030c0031301c40104003f0100cf0400030003c304300c44c03c0314c04133030003c1c00000040100d0d1000001400d04004003054f40300c4c04c1043000104000050100d00431c310004000500c004000000311000030000770c0000000d1c0000300001cc0040030d31007140040004430730300d30000001cc0c000030c447001c040cc0440c000c004400301c0c0310f1404c0443503c7c1304c4001c4040004c000000103430010cd0030f400c0003301003100d103110300c330001544f0030000c50001100c403cc0cc0c10000707044440073037c0704044050c0000777d0c004000c031010040003047c00340c004;
rom_uints[927] = 8192'h300f3303014d03010030700c001fc0010300c343011001144000000700000041000145300000000005c00043c4c701c4c140c00543070000014700400001000000c0304100400000001300cff0015c0c00010cc00f4f010f43000c54014dc4c11303044d03003144400f00f0d10000c3c153033f00c30001410043fc14051140c0cf00430000010000004000c0000313c0000300000300101c0007c0c0104340500440c10400000404401030000c0540030003c300c000c003f40000c00100700500000103404dc0004000033f730c0000000101dd0000f04000c0c30c40150cc0000440430140f003d4c333001003030c00110000c31013001000c000f0110130053c00c70f1f00c0ff000000c000c07d07000f0305034000040d00004340c50004c04101000440404774c0007300c000400300000001c404003003f0c400413101000f0103300040010303c1030c4003007000073300c450c0000c001005c33103000d000403000c04700303000130000007c00100c30007000003040c41c0414103400c0c3000000c0003f3d0030000000003c000c50040414000530000f0c430c14301100314000d004100c00304004013340003010340d0000040011d033000d0040f4040100003000000031c4c0000d01f170400c404c4040333000004300041fc01040000c7033000c1000c00c043c0c01f304000004440400c304103040350000000c341010100010fd0c5c4000c4d0000400044c30300c3c10043c00003dc00c00043cd0303000101400500030c0333301003040010000044c00400c5740010000004c04001001700c000071c004400000007543d0fc0c1003000504013000001301c0d440000000d443403c0d0001130010040c441005474c130000000500040c000000d413d01003c3340054f30d000400c0c1000103000000001000ff04077430043000003c301070300370c00c00003d100c301cc0c00c300410300000f0003c000040c07000300000750010d0001000d440000400300000001000f1000030000c0440d0001000003c003000d00004d34c0c000430100030000c003c00003100d000c000073050000c00003c00000040041c0010333040f000000040073005040c100010c0000000013700741000140403003c00003c000010010000f000700010ff00c1003c003c43731cc100303304700400f4c00005c0c040003c03000001341000010000c070c0003c0000c000d330001000033110c04031300030100c7400043470000500c540400053c10c0c003073013000001c3103403100000000011030c04c000c400000000f330000003000040040f0f73400d0d170007c3f04141030733400100c004043000000000000f0000001000000400c00000101000000300004003000003d0c100000003000000130000c00c0c0;
rom_uints[928] = 8192'h10dc3000001313100033000473000034cf3114c000103074000400000370330000144d05000030001c040005043c03f0c3dc1000400c0c1300003033100000410310370000001004040030304c00c00f100000101c07cc3c0c0404700031331c0000d0404d010f70100cc0000d00300003143f01030c3cc00c000001000004007330500007c0000c0c00000c4f00005000300034003030000d40300040d00c34000000110033c40104340400000403000031000000c0001f0c000000000c000003030044000307f00d000100334c3070033334300000540c4100310013c40c0734330000003100000013000f0cc000301d133c440d4c00003004000d001000034c1050100c0030100000000c10d30000000031073c0f00001140101c1c000010000c30000c00d010031f03000031c3000c30300c00111c000040000c3c040c3c000100001051000033304d3c3001430000000c00c03c3404000c3c1c300304000100cc0cc4000003043c00074150f013000300004000d0003cc00110c0c0c300c00c330c0c0c00000000301044040330000000330000004003700003cd003df010470000c05d03300030000c105d530c10000400300f0010f0003000c03c000301050f3000000000000f04001c0010150000001007113703000105073c30030003301c31030c311f0034030734fd100430313000444730330f1170001000c0041f4430030403100c00c300010503040547400400c1000f00503003030c001000500dc40005c4030c0000100c70300d0d10c41000003f30cc003501770c000f1c0310070010030d0300110c0000c3f400000003040d0d00000d007110c5400000c33304010700cc000337400043300340cdc30441003410000130c31d0c00303000140040300300040304000410000000003c171c000f1c0c00313000470c1d00c33300030403c00c33cf70d34d003c000c30330000130c031000301033033007d10450000000003004000c0000d00f000330000101440100141c0c3cfc000100040000034f3f00fc0c00001000013300340000334010300c040c0400343040000c0415100330001c5400c0cc440000330c00300c000730500033300301040c001400000300071301305c0040301c300001c4cc030040400c3015c0070f00414110017c304003330100010041000010034000304300000300404c4001c40d3c330d003f0110f30000310000dd0c0c3c0330c3331000040407003000310007c303000530f03000140130303c00f00cff03410030fc000c100c04041c004000405cf0001100f30c10303f0f303000701034000530001f00101000000c0000c0cc0c30440403310330010430011c000000004010301011110c0100041030013c30400500f000f0000000335c404401030130c000003034c30310303f0c03cc000000;
rom_uints[929] = 8192'hc0010000ccc0c000003000c5c404c100c0000007c301c030040000043000c00000c050c504c0003000401000140cc0300c00c3130400011040c1010c04003000c007340c000000c0000013044101010000c001000040000000303c00c05030100034d5040c00300c000130300303000c4000004400000350010000c00fc4c000300000000330040000c000000000c00004000000000004c340000c0f00403000d0030400007030070004c00300013410000000c0000070c040301000000c0c0001f000000004c00470000400c10000f00c01c0c00c0401000000000300000410004000400000000c0000005000d0000314c03ccc0010001004100400041000041000c30c0000401000700c0003100001430f050000c4100cc0c3000710c040f10c30300d0c00001001f441000000c07400c4440003c000010100c0000c030c0cf4c0100030540001000110400000000c041100c0d07001cd304010c0007100000c004c0300000040303000c411101000c0c00cc0037000c00001000000400004c000c04c0000304c00d00c0040003040000000c000001000010d0c0000cc3404c4c00c03c00100c00000010000c00040c030000000000c0030c103004040c00000c0000c300000d400340001c000c0c4000400000344c1c0004000000030c0c0434c004000104c30313c00100300000100000000004300c000000000c43000f001030000003000003100041013000000c000001001c00001c0340c004001c000f1c4303033000010003c00100040100000000000c0030300000c0011d0034c000300300c5070400cc00004c000440400c00000001000000000c0001000004c00003000030c00cc1000041034104dc00000f5c03c0000001c0c04c00c04000c30100000430f000c004401000c000c003c003d0f00c0010c30000f004c30004c004031010d00c000300c000004010031000c0c000000c00447000010c0000c0c0014000030000310000100041c030000c000c4c001000004100000000c00010004c000010050000000000010000000003000030010d50000000000c0004130000010000000c030013000000331030004000030004cc0c000530c3030c0500000c3c0000004400000c40400c0000c003000043334400c30000001c034c0704000431000000000c00000040f04040410400000100050500c0c0c00c4000340d0000003003c40c00000004040004340000d000c00c0040000cd300300000410004000004000000000400c304c00300c00000040000c004740400300004000430000f000c00000000030003f00030001400100040010031000c00000c0000d0c0030c0c30c00000000c03000004cc000c000300034001000000000c40000000c00c0003000c00040030040001c40440403300410c000400034c00c30100c000000000;
rom_uints[930] = 8192'h3c40000c0030c00dc1300c40d01c1004000c30d0c00400c00000c000c0c0104000100c00c0c000000cc010c0f01000000040f03000c00014f400c044000000000040000300c000000000cc54d000c1003004c010f4303434000cc0100000300000cf100000c0300000300000040130400000403003c0d01000403c00f0000004c0500000304004000000c0c03c3000d0c03010000000c01014000000503040400004f0000c3400104ccc0000400003007040f0000040004c0000c0c0100c5000c430f0f0300000c0c0301000c000c0d00004c00000f430001c004400304011003030000000c0441c000440dc30f0c040003040c100004000300001000000c3540c40cd304d100000000040c0c30030f03000c0000000001c00f00040c0300000000000034000cc0000001400c00004c40000134010c0003c00000c04f0f000c0c400c00040000040c4c110101434044440f010c04c5040c003cc400c0c040000444000001000c40000000030fc30cc00003014000430000044001c00c0001cc01050d0440010000000000000d00c4c004000000000403010040004ccc070300040f300c040c0cc400070c0004144c0000000f01000004110c00040004000c0fc10c4cc0c4000000100100000000351c0401000004050005c00c0003030101cc0003001f03cd03000fc00c0c000c0030c0000110010c000405010cc00fc13003030c0003000c000f0000d401040400000f400d000f0404040c000000010c0c3c0f0001c300010000000000000001010000c5030000310d0000c100050c004303000303000007010300c100004001000400c0001cc500000001040c00f00cc1000000000c0f03000c43000c00400400000c4001100c400000000400030017c004000004000c00c00c00000c07c700040301014100000000cd0000c000cc0441010f0c000c0305300004040dc7010300c10c0f0004c44000c000000d0f004400c00d000001000000004c0000000003000c40010c010c000cc5010c0400000c4000c30000005c000c030000c101000300430c00003d0c0c4300c0041000c10504431000050f0001c0050c000005004c00000147030304c004040c03010c0003030404000003c01c000043030040c1000500ccc441000c0c100cc01fc00c0c0c0d10c1c0000c0100000c00004010030c04030303040001040040c40c0400000035010030000040000d3300400101000000000f00010340000003034100000040440000c00501000000c00c0403010300450540400041c34fcc000300c300030d004004c00f030004033001030400c1000c0c00c1000000000cc0c00003000c0100030c01000f00330c0f00c00000053c000000c0000000000007c400030303000c04000400000000400000400341004000004d010010000000030d04000c04000140;
rom_uints[931] = 8192'hc0004000030000f34c470000000041c03d4303010d4f00005041004400000403000517000c0300c3000003010101043700070400cf4131c0000c3000033103c004c14f00010003000003010000ccc0033c03fc0c010500cf45000444445000d0c7d40300000040cc43c00010c003c3010000030cc0c3000c340c0344c00c00c00c4300400100010003c04ccd00014070000103000000003c03050c00f0054dc0fcc000c0000303400c100371013cc110c3cc030000400503c00030c30000c0404dcc410c01000050030400030cc00001000000cc3c03c400c0000c7ccc04d10303000c007400000c40c07000c03140000f10000003c0000305050c0000000103000300cc430407015044004300034471c04710cfc0d003f0c1004c30f0c140000000000f0001c1cc00000f354000cdd30d00c04103fc0c40c003c040c5c4c04503c043c0131c00450c54df040000000000cd00003040410c054c0c070c000c40c1c4050000010f4cc0434dd400cd0000404100c04c03c0434300c0c3004004140403001ccc051301cc000cc00071110400c0cd00000f000300000c00c00000000740000c0040c0c0410500cc0c0c4c044440000d1c000004000003c100cccf4d0037004c0c0040c004d001004c000cdc40000043410404410f4010c00c31c0004000c1c00400c00cc5c004c4000004c004011400000405000c000344030c37440000f0c100000c037010070300000004c001130000c440004004c700000c70c3c300440044000c00050d0007400f003404c0004000c3c0cc010c0c0000c1c15174400340030c50404400030cfd0c00c400ccc040c3c000000cc300410c040c01c4100544c000c40104100040c000000300400cc04000d303330cc000c044c500410100400c00c3000007000000c4cf4001c100014c0001044f3d00000d0ccf4100c001400c0c010c01045d1c0c0311cc0140cd000d0400c0100107431003003d000040c00000000400000000cc400cc045403000000340434044c00c0047c144000c401c0c00000041050004c041c000ccc30cc0c3000033c001135400cf000401000c044340044c007c0100300043400f4031034303c004cc340100c04003003100d3000040440cc40c0c310c440000000c40c0c1c00044000000040c050000fd0045c0040101400c30c00040450100c3040000c003000d0440050100c0401c40c0c1c03300330500000003c0370c00030470c053c100c0cf0043cd01c1434f400044440000004700040c4140dc4001cc0007c00071003501fc0371074434dc00000ccf0001004000041cc00c030000404130c0cc000000c00f00403f4c000300071c000fc0cfc00cc0430c0700c0f40344010044034c00400c770104003c3c044303150c0400c041000040c000040c00000c4c004cc144c003000000c400;
rom_uints[932] = 8192'h1004000000013040000c0c0070001077fc10001300dc00003c001100000d100000000c7c00030c00110000341c00311fc401000004000011311c00100d000300001c4f0300f007f00000040000000400541c0c1f07010330cc0000710cd3001430000014d130040300003400003f0030000030440d17c051103d017cfc0cc004140c0000c0010030040f01011000340c000c00000000130c03c00c0030434030300c4f1400c00d4303000040000000c3303c0c0100c0f10f00010c003000000000c0000cc0004c0104040014030000001011300c03051300300000dd11d010c0040c0f040c5c0000010300dc4401100d1111054001f0000430100c501411003cd3000040304c47030dd0300401000000010c00c1030013007400000f10030f03001d300000101d13030310d00040c3010c00100403510300000000000004300f0014000c01c0c100013c00c1c3100c0003040040000000d000c003143000003c00c000c3100703c07004011140c0000430033100000010410c00040400050100100f305000004010c0000303710000c01d0004c0300010003cc00300010000010c4c330030400004000304c001cc0c300430005104d000044000000030003c3440c00c0037c004cc0fc003000000f0410c0000043d010004140700000470c03c33000710303001f0000000d001440000c41410c44c400003104d310055000001030101711134c44104340001000005300030000014300c0010400d70301004044c0c4c0013530000000000100f000030004c100000100300000004041000113000c13000000c000134cc13150c0007000700000c1341030011104000c130001c0031004c1d4c0033000003301100050c5700044003017000003c3c05c030000301c004103000000307410401c0d0000c0010101511041003001000003000107cd000000c0003001113d0cc310c00000000700013700310314c3c0000c40003401c00033330000004400c0005007000300c33d400003c44000004000300c03d1074000000dcc004140000d1170443003cc3004cd0030c3410000340117003303001310c10300100301c00030c0040c030c030040033300710010400040410c00c41c1004000340c04d00cc00100004c0100c0100031334044041073037301011411400c3000031c400010c01c500031c0400004c000003c0c0c05dc0000000700001003031044003d4fcd0000013030000010c00503301134f100400011310c30104473030300330704000c0d0000030c01110403000ccd0000000d00010d0050040c1410000404103313c004040000c50043000fcc00c5010000c1000710040003dc01000000034c40043300d003041400147110000c003001c4c0340004053001ff0000100030300010000100004400c00c0c5100041401003c10cc0000c030;
rom_uints[933] = 8192'h4010040c301000000113000000000101001c0010401030013030cd00d0001000000004003c3c000310040000310033400001c01001c00030000330503000000000143530713300300000031300300004000000c74050c00333110cc30100111000d10c43110031303050fc100304000034403710303330d000f500f00010000015000730044c000010040040030001310030000000030000f1000000140001403313f0030130710000130040101c1303d01c370000033017f000333351c0000000003030000001c010300100343130c00137f0030000c00000400000004f000cc3000030000001d00140000114ff3001c1304c1130310000301000cd00003003f100c101c03103003c1f300fc0000030000cc04000d3f00f1c31100310c0c14100310000701c001000000050c00100300300031100cc010c1c11000004c03030c103300c1c10010110350c4c3300c031010c01070cff100c01c04340000000300004100113105003f1000000cc403c400040110c000000010453000000050d31500400010c30141301c50000300011f01000004000003434c11500000c003c00103040013040000000331003300300c0013100d0cf0f1100c0d0000000c43103001303004100000031cc0330000014000004040c0501103001450700c30c30d0001037dc04133c0c004001000f000400f41030010131c0000040310001403301000000c030000c1000300040410530000030cc0101550000110010000011f030f10401041010304300f0000303d0330001104330001003f31730000100000000c03070000c00400000100103003d3750001400000c100000101000303001d400343000c0d5fd000700400000330c410003335f300c0000000010310c01c0000000c0c3300000050003c00103400003300010300d10014001003cc00030c003000fc000f01d33400c131033003000f31c30300003053010000030dd0350004330000c1100010000003000c1000070000000c41000001c00104c000c00000c0503300050d33110100300c00f10000000c00000d000003100001013040301000034331011c030100010030000cc00f00001d414003033000031001d000010440001d00300c4c0fc0f100d3003c05c300101000043c03f41701003c0003000f0f001dd3300c5000103303d1f003101501000c5330010057c00c3c41144000010d0040d0051003000000103530013f300f5d01000000031705001030f000003c0d0c401d030000130111030c004c403010c33000000370130000001001f000001c00130001c1fc0001107000300410c11f001031f10c0330033050000d000500c3301031c000c0013fc3000000410004303103100f11000000377000f155000010c03d0330100111033c0c04100000000010030330001000340103031c03303000001;
rom_uints[934] = 8192'h34f040044374c30c0f300430300054c3c405013015030c0000143c041044430100c305004cfd0004000f00004001003130300c0000300317003343043d0010010c043000fc00004c4400300c0c0c4000001c3000340400000174700130cc040010cf001c000001000744730035700d004003300c100c003030dd00c500041000400403003103000010140330100010030c01000000000730001000cc113341033700c0000f334fc0f043130030f004d00c04100400041004140001700700c00411030c000304000c0430000104c04700040c00c0c003014411130010103f31001030040007f4000c4010303500ff0c30cdfd40440014000c0c0003cc073000c0317740300013d0fd0300c73377cc00c0000d044031040cc0307f3030303d30000043c700001000000000130005000040300c0df0043cc00000450403ccdc03c01000100f73c0c3001f43d40f100301000c00030000fc003000000f0f0040000000000c00f1c40c1d3c000000c07033000371c47301430c345133000f0d4040003501400033c00000c00d0c4004000c113500f0000c0310c4041c000030c3070034053000030c001000cc343d14407c4330003f000fdc300000110cc4000303001f33f00c00070010001c04001f0f04001c7d05000000013000400f0033c103053003000000051f1000105010dc043001030471143c0f0c007407000031c40740700c00300d10fdc0c0dd430400373010430d0c301343344d0d0014050400300040300410400103400040300047003c0f04f4300000450f0301c4c0303400300013c0c1c0041070000100043414c0f00c001c0043c10004000400044c1c5c04d340500000d070000500103dc0003070c0347c401040d0c04000c33d00030000c50100c00013000440cc3005101c000730031c0004030070340000c3005c00f44410030040cc000f0015053000005000033003700004000000040d313c0c000000f04c0c40000000c0040000000400040f440c413530010c043000313401cc1500cc000c00450304f0000100334001140403000447000d00000000330014040c0100f300cc003103044300130c000103c40003040000000744004f040c3003334400c00000000001c730070c0f050005c00030c00d3d3c0c00000d0040d0c01cc000cc0000040704003030c003f1d545000434000400070c0040473400cc03c1040c0c00c0000c0007c0c01cf0dc04c40030344430f00d4000400000140fcf030070d0cc0015000c03000cc01f0d0534c011100304403c13c0041034c000c0140300c03300703400030c00c00c0047430f000d04140c000c000004c40004040f13001557300000301004037dc000300003c03c40c04310c0c000dc0f00c700300d0c04c044041300c1c0cc5100040c03001c1010440310004c00c0000430c01001;
rom_uints[935] = 8192'h130004040310c30cfc001c11000400c310001400030000f0030370c030c4001c044c0103c3004400c3c1011100000d000370050c0050c330004fc03ff0c0cc0f5310050004c00410000115c400c01c30c4030cc0c00303f3043140c0114003110d501300004c30f0040dc0000fc1cc03c03005330070c1c30c1c0d00cfcd3040457100310330030001c004333104c1d5c0000c000f4d001371030403c00c1005df0000007f000144403004003cc000000005c0000c07c331c0040cc003040c00c30000c004000d000030c00cc00d0314510110000371340c0f000037fcc3c0400000c1014dc4100033cc00d03c5f4c00cc537503300000d34c10437c0010000fc30fdccf313050443071c0501003c0033040c10c0400144c57301407d110400c034c000303031c04000444300000fcc040f00c000c000000010c31033c40c000001000003c4f0001310040700010ccc353050403414000037304750c1cc3c0d0000354c1cf0170113ff0c00f51103cf30001400000075c300c50c3cc0004000744dc0c433004443c04000001fc004330c30c0330c004c00fcf5001c5401000030c043f01004034c00000170001c303f0d1c50700c4003f04040400ccc370f1c4f110c0f00c35c3d100715c13000400c30000c343cd30440300300c1000034010c003170001c1cc30003003d30000cc00400004010d000cd00730cc03100073d4000f0fcc000c030004c0000043300f0ccc040350314003030000c1c03300c0c1c3037c0c01103000c30134000001c0000110000034c4d000004c54030003cc0330340c000104f100031100c03000c00c00100174370d4000004c0405100110f0cc100401c001010f0f131040c30071c33c0045370d3c13003300cc307d010c10c41000c13f0c05c00c401c0114f00370003fdc0c50001000010f304c00f430c0000130f031cc3330c07d0030400003cc0c040001d43000cc0c0303100700001441000003000f444f00000d000100c310014004c40403310c110f4c00034000c10000f500cc033340411407000c3003c1100f05f3cc1c030f43c3f103c00cc0c34c4511100103c0fcc000c0c000f0000430003030030501101c73c3c14300f40f113000010ccc00503c1000c30400cc010000055c0c7cc00ccc51c000c10330300f00f440304f4c100003cd040003000c3cd1110c0c0c003373433100530441c3300003300f00c1d430310044000f400340cf000000cd01c000c011030c00400001000740300140370000c40c0403454000030c0c073c000c100c340070f00c4005d30c30cf0070c173454340d10110f401c10300400003f0000300004000300315c33c53000c0030000fdc11c0010f00000044000040010003303000000fc4003000100040c000cc041000330d40f10413000c3cf00f000cc370010374c0000;
rom_uints[936] = 8192'h31100000303001c050f010100300000033000031c010f000000000000504000000044c50011c003300030050104c0c01c303001d130431c0000004c1333400003300700c000000311000331030c004010403c0f4000004c33000030040500001004001d10c303000f30010300031501d3304f011000030f01043004301000100104f000c00f130030c0000300c3010370000000300330100c0030c000d03000000003700310007013000000010331cdc0000010000000113100100103000310c100c300040000000000c001cc00330034007401103fc073c130311133cc500301c530000140000000010000004030403003cfc00334000000030003c000000000c033c000c3c1d100011103015300000013300d01000c40c3333001303443000000f1000103030010000310000010100f40c00141c3030001405c0400110030000030030304c0103c103c00110f0340040c5000310010010d0001c1c0c1013700040d0000c400133540001003000111400001030000003001c441c0010003070c11010300000073001170003004010d03000130000001c005c004c00040f0000000c100170f5000100cc0300000cf7100300007013001f300101300300000000101000000f0000037100140010001000cc0030000c0004f0005010000000c03d1000330000010115001110003c00103f0c01f01d0f103c300f3070003001000373d43303401000000c00c001400003411033534c010003300401300f05300c3c3030310130113130300311300013300c301000000000300004037c0f0c0030030d00000100000110001300301033040000010c0003373c00000700344403001fc03001370430103103003000030010413103c01300001fc00100140000114c0c0d70100100000c1105300c31cd100d3030c0300000030310003c00000c705130c004000000003410130f0411003c000000000000003330003c000c3400000c0030000c03000000300030001000141300004c1300340030100404033030f0010d4c0001004100033000500d000000003014003000000010300d03331011001c00f10c0c00c000001004000c004c3c31003c03330000311041001003001f01001034110130000d33340000000fc007330000310147334c0000d403000000051c113031d00c3430130040010043010100000000331400c003400414000010073300c00007310300000d1c15010130000c000c3441000013001d000040503100f00c03030c0000001004310000301c0030335035113c3000000000001000103c100310110405030000c000c10103041010003030011c3000300133000400111310d00001004f1030c07100134c53300010000f40400014000000300c013003003000330c3c3f011110333104000000000400030c100000c100000000000133004143;
rom_uints[937] = 8192'h11000000300340c303440340000c43c031c300400103000040000004170000000d045c3c00040000031d0c3041000041400c0d030000c030000300400000440403005c4000000f0000000070000441001010030040cf0470303c40440c0100404440300001050000033d53004000003f0400034d0d000400ccff000c070c30000c4c0003c0000d0030500500cc0f05c5c7000c4000040c30440300c000dc40004000004c43c01c00503000cf50350073041100000030c03000100000500000c400cc10000000000030000400300444400c0400100400000410c001c100440c0c0c00004c4c4c000000c040000014c004040f0071c10000000301100000000330400044000c0400c10c40c00700f000c04c340f001110000433000c47004014400070100c0000000000c040003401c04000c1ccd01010001d300011010431000c00010c000100403c0001c0000100000f01400100c5303d0300cc43000f0c000000c101c10d40110c4010f43d4301001c0f004fc0c000000000c0000000300c4c00004001c00c0001c4003000070f000d00000c0000000000d140440403031004c7c014000d04000000010004cc1003040c3033537101053d000530001c07040c304400dc0010410000314003100c40c131000400010c10c40400000c0000c0c007030f00000c0c0d0c3c003400ccd04f7000c00c0004030c0310030414c1000c300c040c0c1c00c0043d0010011c0000100000540004003000110130340d04071000301c1111c130040f4400030510000c1c10000d00405c010d0000104500001140334031f00010400c10300c50100001c30c050cc000004000043cc00c4c0034000044fc100707c3404c000001300310cd00000007c004105c00000c434005050307000000003500300004304f400c0d0f0414030000110f00c003400d000cc4070c100c0010c000004f0c0cd00c4304cc4c00300300040c00f3000130000500044101000004040000004400000304000d4000040c10043304000c01c10c00000c4010c00404000c00c4c00400001c4000d00c0050000000004c040c031005cc0c000cc004000310000c044410f0040000040030cc0400000400c304430d0c0c4000430100cc0000000c0d000000c00c0013000074001403c0000004cc0410d04000030033d4000c000c4440010c0000500400050c00d1c01c30430f00000000c00010030004000c0005040003000c001c100000000c03053000001030040440044101000c001500010c001001c000300100001cd1000000013701000003010c0010cc40100fc004000000004004000140040140010400000f000400400100043f0130011c41004c000000071003040011440000d0010c030f0f400400400c14010000073400f0050100000c40000c7000001c043d01cc300c0c0c0401300;
rom_uints[938] = 8192'h303000000004005c4400003cf4043c03f4cc004110003c100030c000001f30000330cc004430000000500040000c00c40c3c4c0410c04440c0000000104c000000c0003c04400000300c047f00000000040010cc3c130c3000011cf0040000000443c00cd0dc11c11030003c0f0303400000c310000c0f3000c050001030c00014d0104c000000d04c0004401c040c5d00000c0000f030401000004c0c50054130400030000071000c340400cd100730001140000000004c00000c0d401000f0001000c0010000030c0013303300f03037057000cc53c0000030003000300400c00000010cd03000033044f33000103c500330f030c0000c00001430c100003ff10c01130cc0040140037401000c000c340003011c34033000c1400c001000410330000030c010c0000004000000007c00000303d3300010003000c00000c1010000400c05301000d0c00503c000000000000000301100100010c0400c0301c0001000011c0040f0d0510000100100000c0cd0000050000c00c540c00d0031403c0100010000cc340400000c0001050c000000c00000f00cc0c00ccc103140c0013400500c004300c01007100150100c000040004070010c000ccc10070c00000033304d0c1c0d0d10d4100450104040f0000000001f0ccc4c40000c5c00c000301005410000101c0cd010300c10c0030434c000010c3400c05cc00c0c1044701003000c5000130001300500000d4c00511c100c1400000f3103cc0d00c5403000177c0000100c3000007004f4000c0034013c000000001000c0d4f3100151501100c130c00c0003000c0c33004c143040730d10cf00000000c013c100000c314000000dc0303c0000003141000001100000000003ccc0030010f00450004000431050c0100ccc41100cc0c1703470c000110c0030c00d0000031101c4cd5c001c10f00001301f1000c11000c3000c30101440c30000cc5c0410343c0f300030d030004010000033f30000000d003000003300004cc500c0034000c04000c000000c3007301000003c3000500000cf00000c050001010000fc0c000100f0001000010400000400d000007c0001100400003c00103c004010444000101000d033000000001000c30cc04f0000000c000c015100c0c0c0011034c000f000040510011c0031f00d0110000310ccc10cc003c100c00000c00c000000f0001700f0300040c040003c0003c004410000000f00c00103001000f1400c300c000c0300310304300300013441300300d0df0cd0301d0010340c005030300c00005000c0c0cc400cdc30015030300003cd00c00c004df0000070000003c00000003000030000041000fc000110000c03f0c001000000000073000c040c04770100000000104030040400400c001cc05100043c0107f0f01c111040c4ccc0dc41000d0000c;
rom_uints[939] = 8192'hc3300000400f303304000033001004031c040f3000300400040071034c40300005011c4d304310300ff01c340c0031030030000000c001075403440030001403113c5cf000000300000005000070041030050c30441c05541130113030040041433c310033000400140c30040f300f0014501c00003f0c0003030033343500005df00004013000000d3004010033043100100030000c3c00040c003d3c0040440c00000d3d401030340c04400c100333003000c00314000004401cdc300000d0030c031c01044010140004330000010c00011c00107040000000003c330000100050000030153000d4f03130d730043134d0040440100cc010444004340000f0333c3c0f040773000401000c0c1004343d14404300c01cc0c470c074133044700f3c00000450000004701011000014141300030000350001c50f00043010000030030704301c0c0530003010f31414400c7014043c4007010cfc3400000301070c00c4001374305c044000041c0004303c04f300401700001440400f000033000000c0107c0000000030030400010c0100011040000010040f5c04ccd030400300fc300410001030001000001000000030030030701300100c015cc010300c053033030c03c5140c0004001070330c0000c0317300000c01043000000000c3100000c0341d0d0000013c05000300000c01003c100d0000403c303000f040d433300d334c50c0000305100004310000041000f01410340404700004450440040c000d0310001001003c00300d100cc0001c4004040c1010400500103100000000d007d0003451343000000411cc10000000301c00030c0c000000c004400cc1003c0c0c3400370c04003c00000c000c0c03000c1131000c1334043000041070300300c010100c04000c301c000c0c3c0000300c004c0400400c04040d001d1000101030c000001d000c04010c00003c00000430000c001f1c00000f0400103c000331f0000000000c000c0c14030003034000000005c03d003400040003450115000040000003100c0030c3041f0104504010cc400c00400d34403000000004001c3c04000c0c04703000040101000c054000000000000000410400c00370c07003000011c01433404030c00c073000000c01141040004354000c3330c4d10d044c01c41d304000000d000c00f100004c13000110300300f704300000104c0004004c0c0033000c0c000150fd0010c0c33053400315d33007151004000c0f14144cff4010000103010010030010000cc0c41003030c7d000004cc10cd00103340d0003000d034037c0c00040d140c144005d4c03cd007030000075000303047400100530000333c1001000330103010000030003400103c11070303717300340030100c001c00140cc40100040cc3000c70300cc0044d00c4f03f3000c550300;
rom_uints[940] = 8192'h130000000010d01000034510000130c044041004100030000330c4003c01070000000070c50700d040f4040c0000170434d00300003404d40c00404140000c00004004100004f0100000003000000cc410404c30c0fc70044011000100c3010000430000c40030f7ccc04000c0404c1c07403c0c00000c0000344000454c01000c0434003c040004000c0010307c0533c100000000040400400004300100100700740c400f000c000401c10043c030d43c4d5c5000c005003d0000107c00404035400c00000411030043cc000030103400044c03c000301c3004000510130000017d00000cc100c0033c0014cc53300300c0010000300010001004c0400000c000000c0010000cc003000044310c003d033005343700010040fc0034100000340007f4004000c004000c130300001c301004004001100000c4cc0c0044d70004450f0000103004003100c0f031031031330c0004001004d40410040c0000403c4040070004304130001300100c0c00300000710c00f40000014010c0c00000000030cc330704340143140400d11010040400c044000000004c10c01c0c5cc4040ccc015000cf0401000007100c4c01c411001000700004f0c430c00c00040d00cc330c01cc0000100c000c03110cc0400407003004017c1000c4c0000f3000f0340150037c3d40000104c000003c0050040003000410400430130000c0015004dc00004c070cd401c4f400400c04173000001000000040103c0400007d3cc00d3c000100003400c0003404404000000d00000c00c1c3c0433c35001400404000010000100100014001073d00301043000c410c4070000c000000cc0005000cc100c00c00340000000044c334000c10000030d40c0004d0cc007300000c0c00c0100433003000000c00000000c30103430400000403040000000040001cc0c300003c000000c000cc00033030014d0033000dd30700c0c0500100c410c0c443400010c00000000c400000003040003004001434030303340100c03404001c35000500c030d10c0c4c00300040074c015c00000cc00c043400104c070cc4303f334014000004d405710d400070000000000001c04d000d0000070000004000401110000000000000000040100c004400000003451500030d0010c030cc0c0c1440c0300c0110c04010c40700000cc00004010c3040001f003014c0c00000000000041100040c0c0c000000fc0c00004c00003cc4400030130cc0c700310717403c304004300000cc0051033004051400c40ccc114003300434f000000001000103053300c40050c03c000c00004c3c0c0c00041400000010c00000100007403d400c01504400440f4c10000400044c03400103004000044034d4c43304000000004400c14034453c3000000f000400000504040d003134d00cc5703000000004f3;
rom_uints[941] = 8192'h1000400000c10400000003330003c30300c00311d0c1003004007000c3c55040010033f400c001010054070000c410c300c14000cc0300500010c0004000030001400000c000c310c004303051c30040c01004331000130033c300c103c0c0040000c0c0700440013f044013001104004300300000004100c00cc0300040c004c0c14000c4d0000000003c00003050c5c330000000700000c100c0c440100310c040f0000c0f10cc0400000000c003000000c000030044504035c003000100000000000c000003000300330000030000000c403c4140c0030404c001300031d403c0cc00c3f30c00000000cc01110c000070c0017300404730303370c1100c4cc1c3030000400000000d000300030000fc4001c0c300d000c00301011d033c134053c005cc0010d10100300300000c0030007003004010004000000344703341400013c01f04000c04000d0c0440c1c040cc00c0c040c00703c3f14043001fc0000c0037034010304000c0c031030c1000d000440001033074d001f040041000c00000403040430fc003300700030440c00000cc000440f000c443000100c0000cc00c0d01c00100003cc0c00014000100031400c345c04000000001140400c0000043004371c3400cc0c00010030003c0011000310340c1131370030001cf0000c000303c34c04000d4c00004400ccc1000000c10c000403000c0c04400c00d0330c0440040f0300f4cc010400000001070c300400010040007034404c400400403000303000d4001000043430cc30ccc113c000c0044c3050fc40100c0c430001c4c030cc100d000c0c040010c03000040c0d0003c0000001003001400000c040003370400043c1303ccc0403440c01440030000c50003000f030030f0430403305300f04000c07040030d4004050000010400c00100c03c0070030d000c0007ccc000000000004000cc3300000c004f00c030011c0010c000c0414003000400cc0300c000c400000004000010007000003003030001110000c30114d0330340000003003000c000c000130040400000c00040000703003030330f0c4d10000101c411000043f00000400000000cc1000c103040c0000104000001005c0400c0f00000004040ccc00010c0c000f00c04d00300030400c0000000130d04c30103c0c0c00000030c40d0000000004000000c03c0513040d003f000c00000c00040c00304100003c7c0000000000c4003c000d1000345d000004003451400c313703c0003000070030000000300033004c0003c400c400044400530f34040000000c3033300413444013300043000014003c0c74000100040030100003301400003000300000040f000030cf0001400c4c0000010c000000000050104cc4300c040c340c3305344304470330300440f00cc43000014044001304003000000030;
rom_uints[942] = 8192'h3c000c0ff0144ccc303f040cc10001010030d0300d00017c400001153c3001001404003c0004303100000001c4073043003c00000cc00300f00c7d00101040014000000c000c00000030100d33d41c3103004030000010cc0c0000403f0000734d00d01740cc04000c0004013c000114004c0001c03c135500104c0c00003f5030003c04100c431000343f50c0403000000000c0000d053c31003c00300007c15413000c00400010015700000cc00350300000000400000000c43400700c3c030000000c4d4410301c00f1000404030000000700f0f4100000003c0c0011004c300c4300000003c0010dd004301330000404143000c0504030d40000000001400c44040007c300040404003034340001143c00303105131c0030cc3c104400000000c0c400cc0c031c001504000034c03c3003040000000054700c0030033114404c301c1000300054000c0000cc0c510004015000400530003c043400001000013c1015143000003003401004fd00303d0c50000010000031000104f300d500f110003004000c0101000430033c00000000000003053c01000f53000431030000400054050c00c300000c400c3d03300404f0000000070c000130101070053000000cc400d0100041000003300030303100003031010007c0007c0d0447c00010300330403cc3c1303c00013c300037cc000dcc310000041301571701c003001430503c000000330150c310000300004404440c30c00c047001307034c00000040000cc0c000000100c0001000000cf03000004030c0004130d000000073000000f04001030c14010100f0000003000004c00041310001007c000f4c0c0001c00107f000000c0cc0d300000011cc04c3417000303001000001400004100000000300000043c000c10403f3c00000100044434c00030000000000c43400041003030c3300c040310053400dc000104c33cc400cc003000000d003000003c003c3f0000000000c5330000cc4d00f0310d4004fd0001cc0c0444041300000130000d301d00000000400040000404000c1010c030010000703c000c04000d3051000c3001010031000030410050003c300c00000000014c10000400400000000101c000000c3c001c000040100000000040033100105103c141043030f001000114c30510000000c10403400d10c30d00c01500c017004c1c474440040c003dd40c005100330000010000073fc000c053334000000c3c0c33000000000030300004d1401c00f0f0440000c03c1310350400100400100100040004040310001000000310c1001010013000003003007c44d03310cc00101400010000c3cc000400000004c0033154000040070100007f01400c0000000c00000d3c00050c003c0310000000cc00004c133370000c4011000003140c3510000040000000304c00;
rom_uints[943] = 8192'h5c10111000430713f0000c10010c1000fc001003300310040031c130f033cc100003040c040410001f1011000300100dffcd4011f0430004d00014303c033100011040c40c17101c000000d0011031011304003000313c00300d310d0331c1700104374004000c3300c10430000cc03010003cd10403030c0001001003300100100d5000103030140000000730000403003130430030001300c3100cc000144150003000151000003030700400003077013f0434000c0010d0003c4c0d301c030030300333c07430300410400cf003303040141004143114000001c40c730401c07c00100300050000c0340c00030c010300017c0434001001044f10303000300000000014140003c4311c0431000430110c0c3100147c05001f001c1f53400010000c00c0015030101c013440003303000000000004100001010f50cf00040c1043330007304000c03040500030003c0c3113300300310301300104c33033001004000f3100343d3105c0cc013001d0001c0000c10c0c10007c1cc40330300440d0030dd51000c0300300000501110101300c030c300dc4011043300c1100014f033c000000300300003300003101c00000c0401750013c030003030300033c113c33031000000010307010140000043104103c170d05101130000040110c0c000300053c013005c4310c3f30c30c1015017cd01010310000040010000000cc1310300c0004153d34140113004d143c7040104500311410300031d0013050040c403c3000413c331000d4037001030040533f0003033331004c131000000d11f00010110330cc00043c00040f0403000c3c1100031c30100c0000000c3d1100c41c01443c0dc03c0000001004010dc00c010433c001110100030400043d000f103c003030010001300c110c4300130d1ff0101000cd7c100310c0013c0303033c0004f3331d3001433073317010041c101c0310c03300c010000004301103014f00d03050007000010104110c0000004030cc03104f0c1040033d30003030303d00001030300040011000073dc13003300c3300004101000000c030404c10303010414c03403c000c001313d0f000001100000010031300300103f00033000df03c0011000010043c0c101300c33000130103010013000400013000040311001c131000c00400031310f300404001100403013d305c30133c444f00400c00d001331330000100000431d0000d133c1c330c1ccf013d10011400000d00107d041301043033000000340100303c0001010030110f041700003000c00311010c013c0c3c0c3004f00300000d411100100700f410037f00d3000000d0000033d033001001c000341310000030000303100000004010000c30730c303cc301d01010140004300103103c0c0c30043030f0047010030000303130c01cd0000c003300;
rom_uints[944] = 8192'h1110000304007175303000001000000030100014000001000c70d0000f4400000c5400110734100007300104050c0c1317100c340400c4101010300f304030144c00c0c400441041300430330034c45000c1003d0330030c370000301030400104d0114313110370100503103001c5000400010010031c054530f1c0c14000043033c0000d4314d0040400431d331400400c400000030304500cc100c00cc03000300434040403403030404c03741c10357c00000c30d005304034c00000103410300003d004001050f00c710440003000f3007010c31304c0500c030070014d01300034303f00004010004300000030005010004310040130000440101000000c0c114c140f345000303004cc1300100000103003001005040400d300d0041f04c01000051004c00c001030300f003000301000c00040000400351005c0104004100c0030100703300400c030100003f000000433d00d40400000007c303300300c0c0071343330f30000011000011c34cc3401043000407c0d0003030044c57570013ccc4000000c41101c00043cc0030400f03001300473c0f0700cf00d0150100c10071cf0000050d0000430cc03100003f0304004504030300cccf41c0d30301040c0104410300130000300300c5c0030000cfcf311140000000c1354d00f300c700001304d10350010013000743000303c340c003000300100140d0510000001d1300003101c043134000000070300043514301304c0403c1044030c1700330c00f03f10000004300410000007dcfc701c0cc4d1040c4113000010000c00003c00033c3000c4000c133cd10c0cd0cc34001033403d30040443471c030000c0013170010030000010040034c0341004c0001c34141c117c000c00013030030ccc3c7304f000001300300c30140c3070341037c0004000113004000c044c3530000c0001700030404f300c0c373c03003cdc0400703010044010003700f14c730701100cc01cc3000003010000340030dc00c000000017000410007f04333000c0300c15004c00403114711400c0c000004c101100401030110030c7c0004003c0001c30d074f0010c0431000ff04c30c1003001305037f0030000c30310303310c7f0001014331010000100301000fd704055c51000340003000c00017111000c40f00d301430000400000c00000000343001100003755c010030300c1000303d001f00070000310c00c00f000c1c0000100c00c0103000003c14cc00440004c010000040c43040003c30300404034000000100c00030001003f000040030440433cc044100c0404000040415100cf03c33100100430c3000000c010010403330d03f04d100001010cc407040000014001000000c0000040c0104100c300c03403070003100041c00300c053000d01430f03d04070c317000500030040;
rom_uints[945] = 8192'h4c70c0030000037701001011c0303000d0300400000c1c01d30010c000d1c03004004470400400003103f0070000170cd30000100001003000100001c0700000c1045070000070d040035003110ccc0c41c0c0403011000005c0d0d030d000710000f140c010c43010c3000034c30030104040c04050c0c004c0011400f00000c0511030004000400030034000100000003010300003003c11f00000000c0010001030701310f300303000003300c0c013334030000033d00000000c7030f0c00df040c030030000000000013035001001d0f01003103130113300c0003c0300000003140430300000000c004050c03d3cc000c0310000400100f3004030000f03c0c30004001300500033101071400440f500040130c0cf70101003000301c00010f001d0c0000000033000cc10030c0043f3010043000000c0007000001c000040d000000c3005c0000310c05070300003fc7000500500c0c0103100300000f00c113030c441d40010030370cc00c100040000001cf001fc10c00000010000703df3035c1000d00cc003c300101cd43000d0000000d0110010040310d300d03100c04030500001c000f050044010c03033301c103050c0401300301001700c0114305cd00000f700100000100030401110303030f0c0731000001010c3f011300340500d00401c70d0c0300004c004500334c00004c10333433030400003005001000fd0f3104107c00000707030000051340f30c03000000030ccf10000c0007005f0c14000700103000000c334100d0310013130001040533030500cd015c114330010000010d0c07040330730d0d040c70030004301c31000c03031f01100101044c01c0040c000000040cc100040300c30c040400300003043d30001c07030000400c41337c010c053403000100000100000c3001007300015c00040f014000431c0cf0300310010000000500000d100c10000104040d1c07300003003000310004000c000d000c31003f000100404d03c10c00030704000f01341c03430033000f000c0101300000000013031d004331040c01000dc0040c0f03100c0401d3050010030f00030c30003300031300000003000c001030004401400707031c000005430c10070100000400430c3040301c350c10300c310043000c01040403303f011101030005c30c030000c31d10010310030c3010d0330030300303c0070c00010003430003000001100d301400030001430c4101000310011c301c1001013000004011040010500d03303731043c030c3414004d0c040001031000011005300f1f04c33f00001df30001f00047001c04000704000c00000003f0c3130c0d3100000d04000040000f0f000000040103004017c310011c3300010100000c1300301d000c0d00cc030011f30ccc030f4003313047400d011007000000;
rom_uints[946] = 8192'h100000000000000405030c0c10111340f0000050400c000000413000110c00003000001030000400c3050c40511004033300004003300000000000000434003030c01d0c00000010000000500300c300041300003011001034011cf00c10000000300110000001003013f3000030c1400010004c005330c003f10000110010001c0010000110003300000003100000101030000000c0001013f000000f30040000000105000030440000001033103050000004c000004030010000c00c004000000c30003010400c04c00040013030c01033303003040030331c000c10000330000001040070c000000000c304d3003400103403000000000000003400100004ff003c30000d400000030cc0300004000011511010003f0003100000d0c030403014300000001000100000330330300034401c0000340000f00000104003030010001c00100103000010001000000010c004c00000f01013300cd01030000c30c050131c00f003c000140c0070005040003000000000000000c0030000401c0000d1303103000000000000000c00c3071000030000000000334000000c040000007033300430000000500004c0000330c003100310c0f003000c10003010300f51000000f0000030000c000040000005100c00003000000c00340100c0f1001133103310303033303410cc1000c100cc3400000c0410000003f400c0004000134000033000d0f303003f3030030c103010303300c5000c0000000000001013003403400cc10c0c00001000040000330030431c0010000050001c30000f000303413510300000000030000030000000300010301d0c30000033ff30001f00301050f000301d30000000003c000501000d100010301c10003000400304003000000c00000c110000104003303000501034100f54300004000000000000400050004000003030000000c01033000c003000330310100010c01500400c0030350000d000c30f0000c0103300300031703004030134330000540cc0040f11044c1300000030300030010000001000103100000f3030000d3c0000300c00004000f0000100c31c5033004c0300010000c00000c004300010300c0000000000035300000410000004f040300001003c1c0030000050005c30f000001c300010443000000004f0403040c3103100300101c0c000003000003c1c000100040000000000501301010004100040100040c010003000700010030040f040000000001c13040030305100cc00400040300030400100c03003103cf4343300031003c300000000430cc73000300c01003000500000300000310000c000000400c00000300c0105010010c030043005000c7030040010000000000000011000c05300404344330004303030c100000100103c001040303450000030000000335101045000000000;
rom_uints[947] = 8192'h37c003000ccc0001030000003101dc00300000101d0c333000031c0104c0331c000305000400400110040000000004030330001430000000013010c3000003000410030300010003000040c3000001100401cc343000d300041c33c00005000500100000100003dc0000130c0c0307030f0100350c0c000000000300104c30010730400010cf000c0001000014000050340100000000d0000044034030001c0c00c04000030f3c104d0f110400070305300117330000003730010134130f00100400040c0c00003000300000c00030000004100000100400c403000001cc0400074400333c3010030000000410300300430311000071000030004f340030000f0100001014700300000c00403c3100c033100040030d0040c00c300037030c10103010000001100f031cc00011d4141301030100000000003f40130000010c000c3404000003000c0004110cc444010003170f000d0005fd13040f0c10300040000005cd40001430030000c00507c413d303130307000f0000130cc0043300000d00dc0010000d0d000003000003cf010c0000000c0030000c57c4000ccc10043c1000110004001000303c0000c00000c010310c070d1000010003100030010500010104030000013410010000000d110403001f001031000400003000000c0040043031400c1703cccc10040cf330000f0c3c0d04030000030d00000430000c000c0104050010013000000d1c1300101000c13033400f10040005013c0510100014dc3c0300000000010c00000131033d0003000101310014340003340c031030000dc430003c04004c0404003c30c00000010030cdc0000104c401003c10003300043003000f3410100403000c1004fc000d0c3c340c00000c0c000000141c14313034000c0700370001c0c33f030011040cc0cc00331c0000330013000000303300101c300cc4c0003c73c1104033000300c0c00c0004000703c3103d00100000100c040000030500000003130c100000310100010100c3310f000030000004000301300c00000013100c30014c31440011c401050400c100c000113c400000d30c07c01c0070c4103cc0000f001041000000331033004013001000000c3c1033000004103001030c04030100cc3000101335030547040f0000c0111111103003000d0030c00033041c03130100000000004030010003700c0000013c033070000004000300100001003c7000003c010fdc030030dc00303000000003001f00040400140013c30d30103c0400004c030300c0000c010001040c01030c00440c0004010c1c00000300000d33330407013100303c0001000103310040300f3f0011040400000300000c000c0c04000010c3000100003c403330034c04000c1303301010341c000000030000c1340310c00c01333700cc3fc4331c3c00000030;
rom_uints[948] = 8192'h330040000c1144030cc00003500c004000000000000d0c0000c0300c0cc040000000c04c007c000030c0400c000300cc4030310000004d0c00c0000000004000000c0c10c0000d00000000c43040cc000040400054040c4000c00000000030400f040044100003c000c03000c4c0d040430404440440040400001fc04c0c0000400134c4000000003c00100c000c4c0047c00000000c00003000004c103000c000000000c003ccc0001c4c00f04c030000001000000c000400c00000c000400000c00c1c100000c00300000000000c30000c0c1000cc00440000c0313503004040400000100000000c000f000044000001003000304000000000c00400000cc0003000000c030cf100c00000c00040c000f00004f03c0c040440c430c0000040000cd00014400000414000300000000004000c00c00c000000dc00c030c040c0003c03c000c40004c0700d0040700007cc0000000133c000000534003000c010040000c0044430000c400c10453c1c000401000c0400f000c0c470400010c0c0f0000001300000000c0044000004044df00cc0000000c00000404000000c000000001c0cd000005003000000001034004c030c0010c0000c0000400004054000000400c00410450000d0100000004c000070000f1001100000000000c0000c00fc000400000004000c000c500000c0000c0cc0400000400000cc0000000040c00000c43000000000004001c001d04c100000000c40c4000010cc033c300c0c00404c00433cc000000000c0005300000c00013403000030400d4310000001f070000300004003000c34cc00400000000c00400c0000000cc0c030001310000c004000000000d00430c401510000400c1c3000000c0c00c0040000c000005004004000001c00000f0000f00ccc040000f0304c4000c0c030c000c0c0010000cc50005c140001fccc00300000dc0c1040c010300000000030c00040001000003000000c0000000cc03030c0000c00000050000300c00004300000003c00004c1c00000000001004c4300000000004fcc400000000004c1040c00000c40c0030c04040001c440c440d40c000000c4c0c000040003000000000000c0034054404300050c00000040d000c0410400400fcc00000c003c00c40000040c000000c00c4c000c0004c044c00000000c03500300001000001cc404000c04700000c0400300000000000000000c030000034000cc0100c0cc000c30c000000400000000000344000c0000c00004c3000004c300000cc000004001000000030c440003cc0000000c4c000c4000400000000000014c050400c0c30f0000000000040000c0030400c10030004c01c00000000004400040000c004300000c30c040004f004403f14000c000000400004000140c00400001c0000300000000500000000003000004;
rom_uints[949] = 8192'h40d00c0040304010003100031f10110cf700300400070c0040103f0001fcdc00000d0f05401c000000150000301434013f00c07040c0dc05c000ccc0c7100c070404107c004c0041c00054410c000c3c003f0c000000003070171c0300f110003f03100010c43c0010003f00000433100000c0cc00c0103304000400d004cc0cf3041334400d00c000000c4c0000100cc0301c0000030110003c15c4cf050f00c00000511c30304100cc1c001000334404340cc0000701d704c00004050c0400000f0c0c3000030305c000101c0c0100000c0c01f00f30cc013d344300001734c004000c30d0000400040005c00c0404f40ccc000003000c34403400001000541c00103cc330c034040c03030c0404c0c0cc004c30cc00003307040104000000007f0c000cc34110cc0440000000050004015c04c410043c140f10c0c030000c0010000000300030d00030300100040c000030c000c0003c000100c000c3001000cc0101000c0003c00040001c034d041344c00033c0700400c3cc0d0000cc0311040d0003d0c0c004300c000c00035f0c000100000c00000317c030c40c3f0c171c03404400405c3000001070101301300440cf000300000007000014001007014100000c00001d04070400cc0000140d000000444000000c001400330000401000000000040f000c500c004004040010001d4c003c0010104000003c0400000d040c330000300c31d1340c1410003000cc0000300c000400300cc7f430500d0310130cc0d4cc5d000003c03304110003d704041cc40d00c0c000000700340ccc0301040430040000c304f0d040410304400000c1c304000c13000d4d301700040f3404c50034040000040c0c0040000430313c010700000c3110000330dcd00c300400053c10747003041c50013c00c40c15300c0000c00000300c4c00050004f10c010c0000110005300050000c000c00000c0001c3010400134c0704300041010c1d00000000cfc0004c04400000c0100004df00111004003003050c1c100c0000000c000300001404d4000403070c0c004d044c0c1cd0001c3c4004c7040417030c410c00000000000f000134155d000f000d00040430000700c33134043c030113014ccc1f0c44000f313010030013c001c03c0330040c000c0c0c4c001010001c10c4034004003403c70000c003cc0004143030f40c010c000131c451310000001000100c10030c003d00003c010041c000050700043100c00303030fc0004000c0000c004d0000c30c34350413004d303c041000c0c0c400003c00333f37033cc00f4c000cc4044c07c030ff003c0410c40001100300300041310d070170770400300c0000340403100c00c400001004003004010c000030c0c0033300701070c4103430000cc00000003700315c001c000c573001c0103104000d0c;
rom_uints[950] = 8192'h1c04c01000300c701300000300003343001000000030030707300000010f0c0f4c0300010010501034403133141030000d0440040000010000000d040c30400c300300000d030030000000100000100100c10030001130374c00430f34131c000100040f01300d30c4371011101000001305030d00037430d30f310044400d30f0000c03000c110000dc7334000300000400001340000030d00001304310103104130c03000000c000000c04104340000000c001c04013310000000c1000430000300d3d30001400014c400100000c30030c00f031300c041c00101000000333000010400007001c11104c01030d71031000140101041070000003c30f3100140d33101400015d0300013031030004333000010710003103000000140000000030000000030313000500dc333000c0041d000000040c000130340c3400030c01040c00000301400000500c0330c00f004d333c1000d330005c004d003030c0001310031100041f0000005100010401f40cc3000c301c0000304333400c041c01300301030dc00000010574000c0c0010000030030104041010017011040130100c1d0004000400000004000001503117d00100340030003403110300000000c00c131c04c00000131010000003400000c0330d0000100130000000010c103100301311c003013130c00c040007300c3c40000414000001330c0003041000c300c3c300013c010c10f00101100c001c10010000040f3c0c00004c07401310100c04d4300400340034000d0000001000033030130010d31000003dc40100030001003c0f00000100c00000013000000303300007000300431300703c0c03001114010110cc00004030041004310c300c030f001400c31003310030010004001300000005441000f1dc0700000010300007000dd0000d0030000030400010441000c4010d0713500051013c0c0033000003100c10c10000000030010040003c0c00000101300300f10c11c100000040103c40330c001007010313000110000c07d30011301c040000c400003f0cc103300c01301031000f010f3011010000304303001005030000c044cd007170100d0100040100345000c01000030430300c0c4d000330010cc1f3041301040c3101000100000000000300c441110011cc000744000010033c000c400c03100500c104100001c50c40000440101f304000070700000400000000000004000330030c0000144c3114c00d013031330c403c433330000c0031100035000d0ccc000cc0c033f0300000000000140000105004010000301400c01004100001000001103310400010d00d0f00000314d300000441001440000001000c00c3000100703030330004011301004c0c103cc0000000000330011d10010c30000030d00f5303170010f70013010c03040c00031;
rom_uints[951] = 8192'h43000001000000004000470c00c0000000c05f0000c3000fcc0300c5c0000000030c00104000430400000000c44c100f404010034004500440c0c0c000010000004000431000100000c00400c5c0004403c0c1300c00400141c0c301010000c0000001404000100030c04000c0c0004d0101004035c0c040c00100c3c00000344500c0c0000000440100c04000040040c000000000d0004530c003004000430013c04000c1001003c0c00001c304000c40c1c000040000700c010000cc004000000301400cc1c040c00fc3c001c04101c0c0004141f30c0000030001c04010c300004140030001030000410050000030c0c0004130040c00400040400300030000c0014400c341400000c0c300430000c0c030c300c30c413003c040c0431301f30000c04340400c000040c000c30c014c00c04400400040c150000100c04c0040005400c000cc340000c3c000c0000c40434040c0407d00c04173c140c0c000000303cc0000f04000c1cf400c0000c00000c000400300c00000040004c0440340c0410c000100710000040001010010004c00400c040cc004c4cc4c00dc0343c101104d40c0c000c0410000c4c1c00000070300010000000044c04500cc0c4004c003003004070c00404001c00050c44001000c0100000000400000c000c34000c05c00c00030c000fc01000003c40000c0c043c0c04c3453040000400c00110103c0050000000341c300310000c0030c40017003010000c1c30cc00400c0cdc0d3d000400400010000c10403c0004000000401040040c04d40400000004000f0c000400000c0004f0000044740400001004000004000c0410001c004c0c01c010041c04000c0000000000001c0c040c04cc000c000c0cc0700444dc04040c0c040c0030000c30f01000c00c4010100044100404000c00dc07040004100c303c00040033000c00044000fc100c04000004040040007014000c0c00000c00140c05003000d410c4003004000000040c00c00c1c0400000c100c3c00044c0c1c000400100c0c0414300000000000001c00c004003c0c0cd4300000013073000c0430103c500c300000300c000c000c0400000c400c0c000c15003c04000c101000000000cd300cc000140c3000003000000c3c10040f040c0cc00cc011000c0437c0001000004400401030c00000c44000043040003c0c1004d0040cc0000c0404300404c0003c000c0cc430300c0000007d00000c143c5c0000c004100030000441304c0cf0003c000c00c0c400343004041c10300000000410004400000c00f0d4c00c000030041c104c300400030c10703004000000cc0000000c030c330c3c5014c00000040c000400043000001404000c5000440c0030d33500000040043c50c00000c0c004340000007017000c30000030cc00030c3c0c0c043c0130;
rom_uints[952] = 8192'h1310c4044730000c40003330300c0d073c0d040000c104c4004c0100003dc70000434400104c00000c1c00c04000c10030100704c001001cf40010c00300c70c0cc550040100000040000070d7440d4300c0f0d004404747134000f00040004c40000c110000000c44011c0300dc0440107040f31c0040c44333c000040cc10045d45410000c00c1043500040f00c07c54100000000400030cc4c1f0c003004c450d0c4c00405c0c00000330c0000c330c33004000034000c34300400c073030004c04cc00000fc1fc0c000030c031044041030001c54004c1003c0c1453ccccc00f3004c01c40004c0f00c0000050c1f4000d300140000410100001500c0000c0c1c3f03400310c4c0c0051c0ccc0000543403300004031f05740340fc5007004500c0044300c0c740403400c300043000000cc404000000301040f0041004c010c034c4000df00c310c000c0134340500c0c5011140cc0fc0f0100007c73130100004ff004300000004c4001043c3f0000c41c00401c3c4f7c340403100ccd000c4401113100013f3c000040c041504000000c040043004304c70000053cc10f550c001001030000003041000dd400f7f0f01073030070c434144c03d017cff34043f00c0004000c010100c3cc30c0f3040d400c00c001c0401d40c003304c0c3444504000c01054c05fc74010000010001cc100000000c0cd000011003013101000c7001001005cf43cc0037d000c4f50c34300000c00030473f03003003540443000c03c401400107103c1c134c3300344000300030440740100c4003041f000400d3000cc00f170040743c000c00050000001f10100ccc3300c4003c0cc051004c00f100040c04000c000004004000c44cc003d34440c030000c0003c44c30f30c300404030c4c000404407040000c1004c00310477000100013c0040404340011340041001434000000010113003fc44003c41c04cc0f0f0dc040000003044c43300000c44035000c00c0fc3104c01c0f0003400f051403cc1c000000f40003700535340c00100000f000c0c07f00000000040004007000003c0c330c010f40fc0f0013cf5d00003c0c0c000f005040c00000000004c00400cf7070c0000440005003004c1c04f000700050c00c04c003000c003404c3c0010000c30cc0cdd4c00150000040f0140c0f00040700040014c004304f0400c4c40003104410010c0031004004c00000004d000ccc3c07030344fc4c1f3017700000400000000c001f30000440003c0fcc1c0400000014c001000100cc044c0400410c0c041033c0c304c0040d300003351000000040030fdc04300141c000340003503010043fc4015f05004d1040cd3000000304cc04cc10050c0cc43030307010401c3c1100301c000c00c301040c0c013140c3004004010f0005050c0c0004701000000;
rom_uints[953] = 8192'h4c00c0000cc10c0cdc000013c400100070104c03014133f005003007c00c0d0040030cc44000000011c0031004fc0003003f0351c1010070013100c1004303c10007c0410101c0c000001dc03000c37100d1c000050c00000000f00001c3c1034fdcd311030000c0003710000c431303c03007134000000034700f1101300003c41d104c00300700000000040c000041000c0c0000c0f30c000f00343000400d0c03004003c00d0300c4000c10000cf100cd510000004d4c0c0c001f440000c73cc0c040000000d70d00c00f0c0c0400000700313c740047f074030c01100003d410c30f10c0000000c30c100c400c3c010130fc34000340330300304140c1010f31c3cf103031cd07004000000000cf05333750cc0404403ff00f0150530cf34003000cf0010f03010010000c0100400000c00cc041030104430013004300440103000c40010005c00404f5010430030440c01007110014ff1f001c1c0004110000c004034005041c3d03430f1430c00c0d40c4400131c00dd05d00010dfc100170133c404340001c000c04030c0031700447000000170003500cc00c4100c130c00014044401700103d030d0d17300004501313400000030c7c4000f4430d0045d01c300c343001443100050001171331140000004110c0f0cf00313014000000d4d000307011c454100c14c100033c00305401dc400000c73000c0000fd4d0330cc0000c344430530c040c1534400013310f3d140400330f54c010cfc01003d00700cc010300003414c01d0c000013c1c00000c33430051030000000340070c04014f00c000d0137000343353030010030011300054300403010500000cc03404033013331040c14340000303000d300c00000401704c33c0030014400300407300c000300110c7f4010141ff133d140d0f0c0030d000010fc004100c0c04070cc033455000303d000500010000330fcc1dc0034dc0c1740fcd00004c044101057400000c0c303540c44c045300f0031330c000f1c00d41c0030cc77544014003010410003000c1010c0701000000000cc10f014430000cf043d414000007735f0150000d01c01000d330003000010c0031004000cdc0030cf003100000440000040070503011cc454d000c0300000cd004000f0307000530dd003010433c7f30040044c0c0000c103700c100400401510400000c00030f1d0010300c01104000c30ccd010043000010000040f303cc0c1c47043100c0000000010340000c03ccf0c0003100dcf4300000c0c731040443430cd330400cc0c000044330000400dfc3000c010c0fc00403000cc110d00730503d010041330000400c33ccc0130000c3033c001300001c0f010c3400000d000c00c0003013040f10700003050c330440c4c000044010433700f30310001340140003cc0700c1cc40c00000037;
rom_uints[954] = 8192'h1000c033d0135703030014000010003410103300040000000c0003d3401000001c3c14d300003050040c0000003130331013003000c40c0300305c000000000041c00c0004031000055c00003314000030100c311031300401043000070414d30013003c70000011451014104c04010001531010000c0001c017000c330003150300000000000100000100001000510000000030000400000410c410100010300d341031c000013000000c303010003034340030d5100010000434100403040030303040030400c00010170034100033300c00003314c0033004003d10000033003c33000c0c030401333c1000000053000040cc0014004030010c0030100010140c10101c00c034331d3103100c30c0043003003c10003c03300303000400000000c0054000000c00130000100031100030001030000c00c0003300001304043133003f4000300000c10c30300c0c033c00f0005001c5001010000450003cf010001c4d003000000003f0000030003c031c400c3c0033100c001005fc303530704010100100030400040504000c1000343c00000000c030143431000d000c1c0c04300304000000fc103403300c303000f510110000011001001000c330100f00300c3c30c4000c0c0010001c0415101030003c30cc000004404c3000040300005c03050430104c07000c10330c00003c104c0400003c01050010004550030c0c30453300040001000030030030c3000c3141330000030000003c0c00000300300033000011000c0400cf000000f330400010c010140040313300300c000430001000311c0004000045000c4400000404403011130000130c04300000001400000c40044001301c0f031000040300400d00003f14c0030f00003040100015330c00030010704440300000001c100000113c3c0c000000fc0000330000011104373f000000040700c10100c0111c0030130d0c00003003103303300103037000031100000f000c100030000300c0044c3c30300000f00001000000f00c0100000f3d030000310000001003c7c40400143011000300001000130004400c30341030303000000d3c000000004140c0000035f0103c0c30017000000c000010001000100c3300c1003f03100001303000403c10300040c0100400141c3050011c170031000000000010c3300c01500300001c031070000003f310500400301c000c3051000c0300043400003c00f0043000003010303f10005530005003333000000400000010c0f13f00010c0030010005dcc03001c0001c11170dc040033010000030001c00100010301c403400400130041d0f0000100030340000304c000300c00c3031031404303030010c00003c003000000030300004030f1310403cd03010303350304030403c00100340000001101410543330001010c000301000;
rom_uints[955] = 8192'h4d01f01000cf0300c0410010f3c0000000050114010701004030754000410303c0c3c4000c04000100000007f00400140333000c00070f0cc00000000c0cd50c00c100010300010c4000000d00cc0000cf007d0cc014440f000000c5100104c73101000c030051000005c030000000c001041034000037104700c300c0d30000510000cd400000410310c00403000000000030040004401303c101040c0300040450c003034034c00334000300cc400000c04c13c310000f4010400300c003040000071400c000c3c00cf0330003741000000300037000c300054001c0c000c0c050000003000c0040010300c4007c4f010d0003c300010c00040000c000110c1d1c01d000c0030d40040300040c4000c3033100c300000c04c00000400d04000d3cd4430100c0c003000d4c010000c40c000c0000d00c030c000140010005c50435c000400300010300000000c033c03301043000400fcc4033034300300700000300400101004534000041000c4300d00c000000010cc103007cc0430c03000c01700001f303004003c070c3030000000000030cc3031300000c0700404d04000300000040030001cf30000040404300cc0d057113000000c00c010004030000030103c0030400c133cf00000000000100c30c5044d305c000c0000005c0c00104000000450cc3000c000035000070ccd4400103cc110000000f0c01000707c40c00010140c307005100100c0337430c00c000dc00400c0c00004000000440c44400030c40dc01c3030310005cc400030340000000c003c000c40340040f1300000c303004034403cc030400c7f3d40040000c4f450000400d4000c050000043c00c030103c000030040040c0d004d000f000300c34000c540517100740c040003001003070003c30300004d4f0c0c010f0c0000000400000c00410313003401c04c030300044003000d000000030c000d01440003c7c001c0000c050301430000310c0f000000c0100c0cc101070f034c0f030431000003000d504000030000010300000c0101c3010fccc30300dc00000000030001c544501004000f07000140004f00010c0c03000040040d0100cf01cc04440104c3c3000000cf074000c7400131000110000000040040074037010110fc011000004f0010030cd30c40c0410007c00001c003030001034000c403c5c00001300f0040000303000100000100001047040d4000010001340111010033311501c0000f05030341730341000300033c03000c044300c0cc0c0340c3f00141000303c70303500c0137010040f30001c003300003011003104003500030000100000c0d0043030cf0014700c5000000c700000301030000c000c044400340030301130100c000c00300004d00030000130001c30300000c0031010310044cc00340c001f000000000;
rom_uints[956] = 8192'h1000f00107010f070003110001030f0100400103000000000010c10c030c10005300434000c0000000f40310000003050303c001303001000000100003000d00030400040001000000300f0400405000013041000331000003000000c40433d5700000050c300030010000001000000000000000101f000f0030c0113011030103400c010044000100050300030104000000000340443c0c00000110c00000401000010c0c050000340040000073005114000003000f0000113c3c0030000cc0000104001000000000033030410000000000010001005130031300000c33030400013301000001cc000c00401c11007001030100000003070400100000c0403004010300000c0c030c0f000c00000100003000500000c1c000103041004100300100005100430000c00000041400040000013000000c00003c05c00000301001000000c53f00030001003000400dd0700000150000c0400f0c00000c3c0000100000c00300000f0000030103000004030001fc01010103000f3303000d040100010c704cc010030040313001134003000400010007000015000001033c0103000300334540000cc0004011310c030000100dc4d30000040f0c00d03f10c0304000c30001303001d045000000033040040030105c50c5030000c0c000000000040133300d000004300070c0030000043000000740000300000100007000330030c0000011c040000000000005000030000140100000c00f01101430130000014070001000001000000003130f5c3041010c00000100401074050000001000300400c1010c0113003400c4005000000300000041cd00010f007100000000fd007c0000030000c001000030000c41000004010003d1000004001000c00703000340c03300000010000070303000c03000000100040d00000000000003030400c00d0100003c01300001c00c0011000011000030000100c070034331100000030000150000004c0303000000003f03c40151400300001300740d0000c0400001300000000f000014000cc0c040000000000540100004000073d003004d11c01000000003c01030510c0300100000010414c7000000000301c00c00c0100705000d0300c70000000410344300000c0d000030040c003400000f313001000d0000d17410040c00100001330405004c000000c0cc0003041000c0014000400000010000d007003d0100470f00040400013015003000330003000340004c00373001030000000000c00011330400001010030010000000100300030040000f003011003300034c00003f0003301c003000170070010c0400140000c0c00000400c10050f03c400c40001010c0010000100c00000011300dc0050303337f100000000100c3003303400c00003000c0003000000100003000000fc0c0d000000000000;
rom_uints[957] = 8192'h3c1000003c4d1c00150031030000000010c00cc103005c10001c700c500034301c43c00dfc0c0003c03c3000c00000013c0001000c003c14cc00000004000103004041007c0c70411300005c040030c000000000fc0700400c00710700031c701071000000410010dc4001100000001000300c0dcc01000400c00330c011f00cd0144050000000400cd3004000004030c1c300c3001000c340003c31744c0f70cc300410c0c050c001000000c33f01d0c054100d00000040c00010000400c0000c010c03014400030d0f30110000d30400004030003f0457c0f1c3c0001400001000103300300400000000370f0c331000c00c3440510000100c1c0310410000004073003000104400c0005c7430003d0cf304fc00c04300000741f344f0c000004000000030303f0d3cc01c1c0c00c0cc1430f03100c00030043c3d0c001000c000c0035041f000d00000330401d004340007000041040dfc0007000f3010300000017104030c004030d0cff00c34300c00144c10440000047dc00ccc0d3c000700cf10f401413401003140000310c41c0000400000cc0000c0c0000400300000dc40000030000700000011000c433c4001174410d1043540004000001040000f1c0000303000f100040000dc000c00f004040c0044c7c3301103003030f3cc0043000000000fcc1174c3c000000000100000c30000005300130003410001cf70100030c00030c05104c0c403c0c4007d0030441c0405143740c0c000100100400c03404030000000000410c404700c01700000000444d000cdc00300000100000000004c0000103000030c003301003133103401c000030070c0540000400c04710010f410001003c7003c130000041040043370474d13100011c0c0cc304c1045dc7074013c040101301f1c50130c04cc00001f333cf000c3013071c00041cc4400100000133000030c1c1010503cc570c03d0010403c0300d03c001000403cd0003400000000430000f00000100f0040f0c337000074405040c000d000f000000000030010cc000c0c010110011c01300ddcc0f00c10330c00003c00440100c07070f01f04003f0000f000500c0044103000000c004014040710540130101300001037000d4c040dc010007000043004f0000c310000750d00c1d0c310100c3c04001040cc01007000000044300110dc0004f0d0101110c3d000c05003f0400014fc0c4000034700007037003d30500c0050c005430c1011001fc300c440103040cc30010c0003000c000004c437130431003000300ccc3ccd00f0130047000010400003305c401000107130000000ccf0100001101c0c30100004004f0c00c4410d0300300010000c400013000000004c10000104c1030c0c4000010000000c3003350000c00000013000d30c0001101043010cd00440000c0000000013;
rom_uints[958] = 8192'h3005010d40c103400cc0050014103c100040c101040400cc0d0100003d104103300c00010000c11700010c40300c0f00f030c700c4cc0403040033030cc004001d0d3000c041c70001d03140c50c300d040303d0000040100ccc04d300034113c00c000004c0000001004003c303c00003cc00714100100000000100000001040c4004310445000400750c0100310103c00000030000140140000003310004030000300500c0400dc0304403000315003103000040c3d00c010c030c000f000f000c01000c001c5403004000010f1c004c0400c4114100c30010103003040d4d00070dd0cc0000d30307073300040cc311f000400000d00001c400000c33001101c0c005c4c0000d0301040003000034000510070c00c0c10300c0701440400dc30000500070004417003c010040010000040331370004110311400c000041400c100110cf00003cd0004000f40010c330000cddc0010f0c0700c1dcf0040503001f00004000000c010c00000c0c3030000000cc0003100c40cc4c00c310c57003d00131000001000304000cf0030c004100300003000071c30000040c00004cc4c0004000dd00031030400c0014c000c00530c00103000c001040000001c40047c710030000041f10000c000c003c4004300c010cc0000010000c000310410134c4000c000c30c01d0c00030000d100c1c140150c0304000000030700c040c0c30cc103cd0c0003153050040cc01ccc03000c013300c1d300444003cc040174030740000000000c77000f1c1003004000000010004c7030d113c0000c0c00c000c00040000c0d001c4c0000000040000300000000040403c0010440440c0310d014cc0c3003000010cf000001030000c40dd0f4c05104440000100c3c000110c003030010c1c3c0004f100740c000000c0001c4000c00c00000c0011041c41100dc000034c00fc30c0541000100000c0003cc403004c400503000040030c400050c01000330303100001030000000014003c1000300c00003cfc0007030000000c41c000010070001405003004010000015030100000f004c00043070004303000000c10040000c00000430000c740010400000001004c0c4030d003001710700001301301100003300d40400130501f000331140c000c1d300040001074400c4000101c003540000d000000c410000030343704004c011c000c0c0000475300c170030000140010404c000030001cc01000003f10001400040030c0c0043d04c000000100c70000c03c00000c07044110300440d0003cf1000003000c00fc4000003100c040300000001011001000435cc03000503000040000040073000000c3dc04c000000d0434003070001000000031005404000030c00004c1005000403000f0c030c00010c0d0003f010043000000000340dc043c10000000000;
rom_uints[959] = 8192'hc01000000300000030040000131073003000000cdc10003000300001003340030000000fc3100c00103c0001c004301c005000c0000000300040c004c004c01000000cd01000000000001040f000d1d3c0110100f0d1c000c00000c00034101000f140001c00f1330010050010f0440c00030305001c010400c0003c30033100404450c0c044010c00100000f144301010c000c00030100010144070c0300c4003c330000c00310000c0400170c00000003017c0000c000f100010f330304300c11003131010030430c0f0c03070c4c00007007000c0001030400000d01000007104000040300030c00c00c01f14040404001000c4100003c040044030103003004c0033303030cc00110c04c0c0000000c30c0001d1c440701310d01c40c0cc00403000001010030000c04000700003c14010300c43310410100000301100001030f100c01d04c0003000403010c040c0004010d33350c0730c7041000303330050101040f030d0c03300c000c010003000000000d01000c1404000cc000040103dc30300c00010431000300030101440001dc003000000000c31c0f000013400d044c000c4c04000001cc4000000c00034001000400011c0013300c00500054c003004c0c001c030043400c700401c3f1040100040c45000f000c00500033040000003000173cc400cc0d01731c11310d000f00f00000040000000d000100fc0d044f0133513100100c043404010f1130c1000340013001030c0f0100410000f000c31c15c000030c31030000044301c70c400000f0001100f0150cc000000f01c300003c000050d00000000c03433c111000000000030330300134303000cc0300003c00304c000000350000000c00000dc0000000cc0c00000001c34704c04d1710035400c100000c0f01d00000370c010f01043c070001144004400100030c000c0000c7401c0041300000101030003cc4c4cc0cc5c03004050c10f00c00073d0c0000030050000003100300103030010031000704053d1003c0101000301000010c0400000000010c1300340300000d01c00d03000000c1707004370f00033101001405040101041f410344044100010003030401000d4003000300000003700001cc000c040df00f01000cc003111145d043000003000430000c4400440533000000c001000500034c0130000000000100c00f0c440dc30400104000c10101033c030000040c4001101000c0401007000c0c000c00470003010d0c0c100d00f003000001000000000f0c00700301030c01cc3c030700cd000c0043014404d340000c0d04130c00040001c30c500c000001c004040003000000400700010010c00004000000000c03c0c00000000103010001d00344c300c0c0030c00000403030000030f00010f5c00030340030030c000074c4003c7010cf03000000;
rom_uints[960] = 8192'h4101000004040450000d000400400c0040000000000000000c0400500100000003c0040400000c0000000030000cc05c0000000100010f30c0004130000000100007000004000000000400c4040004000004000000003cc30400c001340004010010530100000c0300540000c0104400003f000404003300000000000c00001c0c010000300030000f0000004000fc00c400500001000000100100000003000f000c0300000c000040000000f000c300001f040000001040000000c00000000014000d0400000f000c0004400040300000c3f0000014030000c00004c010004401040000000000005c000010f440c1000400000014000030000030f000000c04041044003000c0000400000040000000000000000000310000003c000007c0000000000003000000040300100400000004005c0000100000001010000c000c0304000000130c0c0d003104003030000f0000c030030011000101400c0f0004000c00000100400c00030400000cc054000000c00cc00000105040c40003000030c05300000400000003000030000cfc0100000c0c00140c040000c003010001000c10141c00000300fc00000003000c00000431000440340000f3000001d003c4030c0000000000f00040005c000000c0000000000400310000030c10000c3cc00000300001451400c0030000400c0c13044030000000300004000100040040c40c01000004030000004034140000001050000c440005030000340c34003000003300000c04000000000401cc000041001004000c00000c00003301000000000c00000000000c04400400f00000c00000000000000c003000000000040c5000000000404c004000000cf3103c0000c0050074000d0c0300044000040000000000c0000030011303f0440cc307000c4003400c04000d000c00000000000c04040c401c3400400c000100000034000040c0000c0000cc4000000c410c00000003c300000c03000400f3000000034000cc0000000040f0fd00c300c0000000c00004000000030017f00010000003070000400400c300c030000cc0005000004000f0300000f140040c0110440000000004fc0000040c000010000004c0034000400cfcc000c105000c000100000110030000400437030000004c00000c001c004540040c000c000c040000000003000101000f4cc01d00000c00500400000000000000104f0000003141000400f00cc04000000501000004040c0c0c100030330c0c0453300c000550f100500000030040004000c05003c0000c00000100040c00c0c000300f00400000330030030c00100c43c00c0000000401000000000f5443000410c300c04c0300400000005100000014040450000c040c04100130110c40000100000c0c00300000010000fc5000030c00c0000000000001040c00c00000;
rom_uints[961] = 8192'hfc000000000003c30300000040000000000003004400000441cc0000003700030000000cc000004300330300040141000c03330000c0005c000000c001000000000000c000003cc40400c00100000110041d00400000100041000401f007d00001001000104000030f130001001000000000540003000c0000000031400000000f00000000001000000000000300000000c0001300040403030000007000400000004000001400000530300040d000000000c0000000000000000000c110000000031100c000c0c0c01401003000300700004403014004014c0000010000c04330000000c00030033003011000000000c1000000040000030000000300030003000400c00000014000000c00000c0030c007040004040001113300000c000001400000001000300100cd030001100c3000c0003c400000c04100404000c000030410000000000000000d030c0301000040000c0001000100110c4401000000404343004030010104cc300000030301000cc30101004030003100000f000c040d100045003400004303ff00030030000040c1000071007100004000c0c3cc0000010000030000d0000010003110003030c1000040000c01300c0000f040003000000003004000000c0000000700c44000410040010cc0000c3300c00030c1c704000071003c0cd0400003f01f037000003c0433400c4000f1004041f1000040100000000000c04070010004f4340030110003010000313101f00004410004000f00010700014c003004d5003000c000c000000010000c3430000400400100400000000003034000003100101001c0000041510000000d04400001c3c00100000c0100100003c7c330000000000100000075c0070001440001c000000000000c010000100014000300007c000d4041410010c010404403000000010c005000000d000fc1004100000340001000030c10400000300000400000030000000300000000000000000410c0000000000300001104000000c340000003000004000014f1000c0000c000c7000100c00010003f000340000000c0000040500040000000004500150000c0000040c00443300000010000340001300000040c004d000000303000000031000c0000c00000300003000341000400000000103000040000000000c00010307c000c0000c030500100c0000050000000010300300003c3010d3d0000300410000001003c030030403c00010c40000000001040000001c0070130000c0070000d130040000000c00f0004c100000000000030040001333000000c0001d00001000000000c0000003ff013000000c3000000000c00100c40300000701f000000c300010000004000000400d0001400010040000000403000000003010000000c01000001104000000c0004043f001000c00000000000;
rom_uints[962] = 8192'h310100140010040400c00c00000011730000003040007000c0030000004400000c00000000400040110000000043f0540400f03040307c00041040004c0030004000cc40c000400000013410000cc01030000000c0001070300100000003003c100040003044c011007000f0447010c0c003700fc04000001000043003f0c04000050000c040c001000000004000c714300000000000000040c00000c0c0f040330004c10000000c0000700000004400000c000030003040d30010c300000000c100c4c0000000133000004000404000303144000c003000c000000000007c703000100c00c1cc07d0007c104440001050c000400000117000c300000300c00010cc04400010741003000c00301030003030003370c0000c1404c04400c03340c4d70000c0c00000034100c4c0c0100000c04c00100d0000c000f45070c00300c011010c00300000043000004000d0c0304003c01300043ccc000400d03000003401c100000000000cc0040450c034c0030000c0c0000000c050004070103040300000530000003070440000c0303fc0000000d000d43030004000440c000000100000f00000c00000041050c00c000300010000000310d10000014c03330030000010000000004003000000c000c444400c0000c0000d10000034000400103c00101040c0d03400703000005000100cc0c30040404130000030c0141001000d403004774001c0300d10c010030003c414c140440000707000c00101001000c0d0fc00000010d0000030400030004004c0130000c010000054f4700000100f70704003100000000cc71051c04000100000004300000040f0003014d00400c10c41040077037010030040d0000d00400300ddc0c0003051c004c404000000c000303000104004401004040050004000c0cc50c4000010400000730003c000d0000f3000c30030c30040c0c3003c40c330004400c00000400c00000400414000104010c0000000004030c000003400c00410140030000000041500cc4054c0000100103014303010000000004440c000c40050d0c000000010c4dc0300701000401000000c0cc010030040dd0c00000c0000004400007004417001c00003c030cf70c001100340000007500040c0d000000000c503300001003044d301300300d01000014c00400000000003000010cc00300d000c43000f0341c000f00040d000000010034000c40030010030000470c000001000000000001000000300307000303c05030010000100c010c00040010010c04030033c0014c0d3000c400010017000000cc3d3030c700000010d1704005c3c740000500000300000003040400070000000403000004000d04000404040010000c000001c00004cf00f14d0000000000004c0407030140000004343c0c00433c0100100c40010c01350040c00;
rom_uints[963] = 8192'h3300000000000114000433040400c00000000300000100f000010000000004000c00004000010004000c1001c1000000307000c00000000f00010040000c0000000000000000005c00004000410303004c3301030000000014010440c454001000c00000030000000003000000c00001c000010013030f000000010d000c00000000c000000001400000c0010000000010000f0c4d1000000000cc00c00000000000000000440c010000030000410000000000000000100000010000000000040003c5000000330000030d0000000300000441000d1051011001c40104030003100000000300100033c000c1050300000000000004000700000000101000300c0003c0400000f110000300000510030000440030100004000dc40340300300010000000000000c41003000000c10000000c300010000000f4d44004d030103301403000000444000000c000c300000330c0fc501014f00c0040100000034000100000000000000c03000300c4c00c0034c031003400c01000000000413000031c00001000400c001034d0003000000000001400300300000400001103300000f00004000000500c003110000000011c04001110403000000000040044100000d010000031f33003000c14300100001000401340000030000000c040c003c070003400100000000000c000f03400004c000000400000000014c0000040000f0000c00010000040400030010004104043101030000030404010000450000040004000c3000010c00441000000030000000000100000c07040000010101c0c003040000000004000000000000000140030401300000000004c0400003010100030130c0030c001403000000030000040003c000040000000001000700304400000000000f00c000034000c1300c41000000c00000001c034040000000004001010100000010004000000c4004000000000000000300001000cc0000300300500100000001000000000030c00300000400c00400010400001007030000000000000000000000030310000000000001033c030300004000310005050000004004000004001c4100c00341c10c04310040c000000000003000010c0c0000000000001000000000c03000000000000c1c50430d04c1000000003f00310c00100d0300000000c100c0000300100000000004100500000030040400000001c0000000330c000044130400001100c0f304000001000043000043000f03010000040003c00000330101c000c01000c107000c000301000d00cc0000000d0003d00000300c000030000d000001000c40c100141000c000004303000000c000000000130cc300010003000000c4000700000100000000000010000000c00400004c000c0110030000c001110000000030000000000c000111010cc0000300000000;
rom_uints[964] = 8192'hc0c00ccc0c00040000004c000040c4000040c00000c0000100c0c0000700003cc4f01c4c40000040000003004000040000400000c00000444000000000c000004000004010c00000c3c00400fc4041c5000000000000004100c3000031033004c0013000000003c0c300000003c04000400400500500000000300000c000030cc0000c0000400c00000000000000040040000000f300000000c0d7400140c00043000030030040c00000c04000040040000000d00c000400005cc300f00004030c40000040004040c44010c030403000000000c003c01000001400f00010c440004010f00100000c10701c0f0000c0040cc0c170000000003001c4040044400000c00000704040340030c3c000c0fd047000c4c000040c04c0531310005000c0000000c000700c001004c040401000004000300000000000000100f044c0301c100104000000c000c00c00c0c0030011d0700c0000047000c1043140400c00c0015c03044000003050f0c04040000040c004004000c00000c01c00104000300100000000300040100000c00000000c00000000000000000000c000400000034000c00000504c0070003c00c00400030000f00044001770c0000000000c30c04000c00400300300c300000c00c00c0000000c000fc03100413c00000000400000400c03400d0500f4000400143003c0c0003000300030c000000c000100f031c0000304340300000040d00000000300c44000c40000000400f430000000040030700030730c100000c444cc00000000300000007040c001403070040013c00000000040004000000000d4400330001000400040300000c4c001004c70400401000000c0c004100000c000000010c303005001c3c000c41100c00004404030d0000400c3000000505000c000400000000040c0c0000030000004c04300014000c0cc000000c3040000300171f000003030447000000000000000f0104000c04300000040000000c00000004f0004000040cc0000c00033c04010c0000cc4304c00003000013430003040440000c0700000c0c0000000000330c00007f00040c000000070cc30c0040000c0f0c43040c030000000c0c40004010040100040c0f00000304c0c0040000c00000010000000000030c043c0c0104c00434003000100c00c40000030004000400f7100004000c000400030043000011140000000004000d050303000000103d0000c3044007c03000c0003c40cc010000000f70c044030030c00000000300010300000000c00c00410c0414000c3004c0000c4000004f4003000004014001400004cc00cd7000c0300500000000f0010000000040000030c0c0030c7400033000040000003004000000c0000400010c040700007304000c0100003c0014500000030000400003000c4001000c004c000300000c030;
rom_uints[965] = 8192'hcf17c0000030f00340c0004140010400cc010c0f0c00cc04040f100104004cc000004000340101000003000cc3000041c0034000000040c3c4000040c3000004c0000140040000c0000000c00000cc00030001c43c000000cc0100410c040340c341010f400c04000010500000c001000300c000434c300000c404f500000000c0000100d00003c400c1004300041041000c0000000c014100c140000000c300000000c004000f0404c400100004000400030c0000c000050000040000000c0000100000000001c00c0000000cc00c30000041000331c0000000004dc003300000000000c40f000c0003000004cd0c0f040f7000003000000c0000300000000305c0f0000037c3034040000001c10044004c01001000c04f000000000044c100000300000f0001c001c0c0004030004300c00c01000004000c010041f001040001c0c0001031c00050000070400d00010c000100000000c000410013040140000000040000000c0c3000cc0c300f410040004500004ccc01004103c00c00000c00c0300033c0000000c1000041c00c410500410103000041010c03000c0001000014000405030000000c0dc0c005040000400040101000004c000c4000c0300cc00000000000c1400541010140001044cf40000cf005014c0400c00c010c0000c0c003400041440cc0000c010110011001000050c3c000001007010043000000000440000c000034003cf303004cc000000000000000040c010074004500004000034401dcc103040000000000013500000403000034c03100c001000000c40c104030c000c000c040c40001003c400000000005000010c003c130000300011c1f3000001c00100c00c000400404004500c0304000c14100f003c00340c1000010011000c0c0000500000c00c0c0c0000c00c1000040c00c00014130000c04000c01f400030040400000400f440100000c0c10c1c10c000030000100000c03000000010001000004000d0000004c0cc0c04404340d050040001c104500004700c000c00d00000c00030134010000040034030104c100000340100400400c41301000010003000cc5400110010000000040004000000010000070010f01000300030f00cc040100400030034100f400000011010100100000000c0404cc0c00000034c000c0c00000000000000030c403400c00400c0c0004d700c00440030cc0001000030c000041000000453c0103004300003003000c104c4d000c000cc00030044ccc4300000040004000c0000143440044ccc0c37c0d300c4000740400c150cc000c00c000130010003000014000000501f0cc00c0030c400100000013030001030c00000044000000000c40000000034300000c000000000100000010c300dc3300010c10c100400045000c130040000035c0000c0030c400c000010000;
rom_uints[966] = 8192'hc330000030dc03100003330300001300c00300700000301000100110c10400c0000110cd004000004400011000034107c400000000000c7303000000c0003000001101000000000130003303100003030410d0c30011040000c000000cc003100dc01010000010010c01000f00331000400430010100d7c3000130040000000000100030c100010001000000100000440000000000d100c0300f070004010d00f03400000000000001300700070003c000000000030033330110000030401000c3000070000000c0130010d000004040000010000010000c00000010007003000c0010300040d010033030341000000007001c001cc0c330000000000000000000710510010103000030010100d0000000300001c300d3040050000070c30004000000001000003100000000101350000440c1004010000000000143c3c100011010000000c3000150430c00c40700003000007c000f007050001000100430d00043c034501c000043040400000300000011100c130001000cc404403440f00cc00103010100330000003030003003010000003000001300140000400011100370d0000c000101d003074150340000340113304300d004c010004000003010c30100001000400f3010d000000c00040c003030030404c00000000000f000c0000c0030000000105000104030d4001001001100007073000d304000074000c000c45004003411000000003301fc10400300000304d000c340c01010c1c00c00c100000301d0100010001c0000000013100d00100000003011000053300000c3000100400400104001033c10c000343004f0000000004100100000500100300c0000414000104004000000c0c030d04000130030f0001c0010000100400150300000303010100000c30100001000307100d0007011030034500000c003301c100140000d000010101c000040cd40d00030300000001030000000700001ff000000f000c030000100c1000101d0001030000004400110c040c0010401c3030040010000130070140303300000000400c3000031c1f0100000000031000c0401c003d000000301d0011000c000c0011000c100003110311730000040000500000d10300000c47010010c0000000f00301300033000f000f030003c3010301073105004c000104000107000c03100003001000030c30030000000444110000000003c0014103000000013003003030000310c4030000053010030000001004300dc033310030000030000030000705000d0310030030471000001500030100000000300345c11c0004070001000000030003000100000000000001000c00001000000000000034031004400303110000004000000000000730000401003004000001040000010103000000400000000100c00c1001043c0000040100001130010001;
rom_uints[967] = 8192'h100000000000004400043011001041000400000cc000000040030000040c0000700404000000000034000010007031100000000000000c000000000000000000000c05000000400400000000001cc00000c005140000c0300c4d310c0400000000053c040000000c10000000401000c300000003d000000040c00c70000000f000000030f000c010040000000000100c0000000000300000000000000003300c0c00001d0c00040000040000000010000000000000000010c40010000000c000300000040000000c000000000c0c300000003000c0d01100000004300c003000000010d001c0000040000cd0400c0000300030004000400000000400000000000000000400000c00400c3c4100300400ccc0000010103030cc000100100c10040c00003004000c00c00000040000000030000cc1000000001040103004040000000cc0001004003100001030000000c040d0cc0000000ffcc010c000410401001003007400000d000cf0001000004cc00001000c000cc11010d40c30000d00013c301033c00c00000010000140004c00001005c000c0140c030430c0000010004500000c0030000030000000d000000c0000413c00004c0004300400c403003f01400000000030003014000000040044000000001010c0000040c000300040400000000000000000000c4004c4000c4c000c00000c00300c000114000000500000040440300c00000c000000000c400414100117000000c000040001004001040c00410ccf00040000c0000400170000000000403000004040cc0c000030003010000c0000c0000000000000004c000000000000c000c0c000000000001000000000d350c0c0000000300000c0003c0400400000004c0100000000c000d000000030000c000000000000001040f0000400300400000c0c001400044000d04000101030001ccc00000c000000040400c04033000c0004013000c044000400000d0000000000000000000000000000000000000000407000400c04c0000000c00c0000010c00070010cc043040c00cc00000340000000000000000040000d40c40400000f00001113000140000043c04300c000c0400c01c00c0000c000030003c00000000003000c00c00000000010000000d00000c001040000000001000003000301000000000040000000031c00030000000000c000c0c00000001000c000000cc000c00001510010c110400300000300400004c004000c0000c4030004000100000000000000000100c70c00300101000d4100c000030040400001400c0440c300000c04000001c00000c00100000010cf000004004000400000000c000000003000030d0000000000000c000000010070000000004000000000f10000000c000000c40c000c04cc0050000130000000004400000c0700000c0000c4000;
rom_uints[968] = 8192'hcf00000001040c04300000c000000004000000000304f000031c00c50c000000040003010f000400005003030000040000000000000c01100000000c0041000000051100c00001000000000000000100000c000000000300000001c00300000000430001000030040c07000004030400044400000c3040000000043004010c00070300000000000040000040000001014000000000000c0300000000040103000c00404d00000c11004c000400300040000000000c0000000100000400000000030000000000040c0c000003000000000307c0000000000004000000040000100c0000010000000003004c00033000000000040103000100000300000000000f30000004040140000400030403c04000000000000c000000c0000c00c0000000071000000103000100000003000000000c100c000040000c05000c0000c0000000030304000c00000c0c00000300000cc0401000001003000c0c0030010300000000400100034c05000300000000030d00000400000004400cc40000000700c0000500010001000f0000000700000c010000000004000c04000000000000000404c000010c000c00000f0000000c00000000000000000040c00000400c010000040000010c0000040000000c000000000300000400300001040000100100c00034000040c400000c00100d0000000000100f000100000010c000c00d00000000000004c0300c3030004000000d00000401000301001fc00000010000000000000000143301000100000000070000000000c1000000034000000c0000000300000000000300000000000004000c400000000004000000000000000050000000000004000704000000040001000001140000001004c401c00444000c0c050000000c03c00030000f0004000400000005000c0100000000000000000000000c000311040400010000c300030f0c00000140000300000005000000030000000000c000000000c0000003c001000000000000000000030300003003000100000000030001000c0003000000000c00070000300004c00001000001c00000000000000010000000000301c000000000040000000000000c04000000001000000403000040c0000c00000c00000000c0000400000c0c0004001440051f000400030c0004040000000001c000000000004000000004000100030000350c10000403000003000d00300000000d040000000000400c00000400000444000400000c00c000000000030000010003000000000f000000000c0000004c0004c00c000c050000000303003400000000000c0300c10000000100040c0000400000000000000000000004000000000004000440001040000000010400000000c0000100000400040010000000000001300000000000000003000001000000000101000c000c00000;
rom_uints[969] = 8192'h331000000105000000000000140000300000041000043000000000000000001005c00000000100300000305031000000c0100000000000010430000000001400000000cc000000000f000000001000000000003000001540000000000000001100001303003c1000000040000000000c133c00300013000c00c00000311000030000000000000000000000c0300000300000000030000c000300000c00003300301000c0001000c00003001100000500000030000c0000003130000000c00000000010000000000100000004000100101000040500100000000000100000000c000000000000000c0000000004003300d0c00000030000100000000004000000001000c40000000000300004001c0010cc00000010030003003000c3000010000030003c0000001400000000300000000000000000000c00100000031400000000000010000001300000000c3c010000c1100000300c04001000110000000130100031301000000101000001000010000703001000300100300000300df0011000000330000400000000003310000c0000000c01001000030000000000150c1000000000000001003010400030340000300000004000000000000000000400000330330010104100000000000100000040040000000000001c000000330030c000000c10000030000000000010000010000c001000000000301c0005001000000000330000040100310003000000003000000000000000340000004000000c000000000000004000101110000010000000003000041000003000033000400010000300003c000030000000000000001000000000000000043000040000430010c410000c00000000000304000330010000000301000000000000300000700c0000000004c0000c000c00400c0031100000000c300000000000000c103c01101000000000100000003000000031000010000000c01c00010041000000300070000000000000000000000003000000000000003c0030000c100000000003000000051100000003003000c0000001000000010000001000101c00004000f0000014000000445000000000d30c0000004303000030000000000000000000004000000c0004300010001000300000000001000000400070000000004100000c000c000000000000000000cc1100000000000000f30010103100000000000033000000000c000000010000430030003c00100010301000000300000000000004001010000000013c330000000000040000103000000300100003000310000000003000000000000300000030004000000000003000300000000000030c0030001010000000011000000c00000c00001000000000003c00030130000000000000300000000000000030000100000c003000000010000000101703c100003000;
rom_uints[970] = 8192'h10400000101000000010100053001300d00c10003030005000033100c44034000013000113c000503400003c10000400074000000c0c00c400100000000000000000c1c00013300000000000341c1030000413c1f3003310000011000047030000410070040001c0c00000000010000000001030333c000540000d00c00040004413f0000000004300d0000000c0300000300010003000000401403410004030000000c00051004c0c30000043000010100300d00000500030cc003411000000000000000000c004300000000000d4000040d010100100004c0c00000000000430000000000001004000007430003000014400010100000000000000410000c040300000010040300030003004c0003000370040001000400c0050000400000c0400000043c00000c00000c00c00dfc010000000000010003000c400d03030004c03004000000c000300000100000001700030c010c000c3f0403040000000000000000000f0c0000000000000000010000000000000033c0044000c000010001000030040f00000100400001100003300000c0000100f00c030d30000300c40f00c3030003030000010000000003500003000c5000003401c3403f0003000000000d0003c00000400000010c300000410300400003010130000003047300043004000000000000c004030040000100c00307000000700103000010000000003300000c0030030003c0140104000c00004000010c04000000000003430000c000c0c0401000c00000003000050003000100373000000000003000c00000045000000310000004000000700140c0700001010000400d00040c030001000c010703000000070000001000000cc0000300004004030000c0c0000101000010030c301000000c030c10100340000c1401000c3c0000004000000000c000000c040000030010c0c3003cc00330c43000000001030030001c3c0003000001001101000c40001300c003c0400000040000f4000000000c0404000000040403000c010c00000000007000313000000001000000031c0c0c40000004040103c0073003000000001000340000c040000100000400000000000001344000000700030000c00130000004003c040100000030000004000004300000c00000510c0d000000040c1c0000c00000000000000003000000003c03040400000c004700100100030003000c0f0c0001040300043300100000013100f100c004050400c0040030110000010c000300000001000c010000044403cc00000040030000c000000300400001c043330130000000000044001000100000000d000000c00c000f00004f003c000400000001000c0c4340000c0c04000000000000040110c030c0030000000100000100000000000007400053000004000c0000000103000f000000300000000;
rom_uints[971] = 8192'h4040000000c0c000000000400003400c000000004c00040003c00000c1440000c0f0c4c00c0000104400000000010305c0000000d0000100404000c00000400341050000cc00000000c00034000040000000c4030040007d400440000c000001c00000c0003000c0010000000000d045c01400c10cc0050003034000400000440100000301c000004000c000000000040100400030c003100000c0400000004001c0000000d00000d0000000c30043000000000000004000000000000100400000c043c0004310034c00000c0040000000000cc4c000c00040003000100000c030000000c000000040000100c0c0000004d00004100005c000000d00400040300000030070c00001000c0000000000c000004000000000c00700c00003d00000400300c0c10000000040c00cc000300000430c00c541000000004300400050c0c0c0cc00004f0004000c0000c00000000003000005400000c0c00000004c0000000000400013f0c00003410000c041000c0000c0c000c0400000c00000c000104077c0c100001000cc040000c00c00300000400000430043000000c0c005000033c0c070c000000000c010000c00c030c0c04c0000000740010000000004fc0000000000000000000100001010000104c001c00000000c00000040000040004f00100c0000c0c0004000000044000004100000044000000001000030000040c00000000040000000034f0010104000400000c000400c0140c0000c0040300000140000004000c000000c004000cc00000cc4004040041c000103004000c0c0000c030000c00cc0000f0004000000f4000100000000000000000000d000000341c40000000040001040000004c04000c0000000000103041000040000c0404000cc40000000004000c4050030000401000001c700010040000000400000c30000c00000000010404011c000000000c4000c404000000040000040400000000010000000000000000040000c000000000040c0c000000400c011c04000d00000040000cc00c00001010040cc00000000c000001d00000000400040100004300000c1000c00c00003c00040000000000000c040c000040003400000c0c000c000300c004000000000c0030400000000000040000cc00404010040000000100310c40f030000004c000700000040000000004c300f000c04004110c000c000c041000000d000400000400003ccc00004004c4000000004014000000040003003400c0001c30000c00000000000c00cc0000000c00c04340cc00040c0dc00c0400000401c4000000000001000c000400044003300440300000000400000c00004c000510000000004c000400400304000000000c40000400000000001000d070000010004000000000300c0cc0000001000c0440000c00000c000c00040c0000000;
rom_uints[972] = 8192'h300000004c040c0000d000c00000d033300c000000cc0000f10004403300300010f040003000c0000040044000ccd0403400000040000033400040400004004c001010000000100400c00010015000000070001701400c0000001c000000000010104003030fcc0cc04c0c101c031040c0404c00300053004c050c041004004f043001c4000040000000000000000000100000000010001c70fc00c004c030f00ff50000c01003c1000c301003000c400c00400030c400330000c4001000001c0000cc0000c0400030340003d0c0cc0c00054000000010cd340cc030110000400004f30000c10000cd103fc0fc50000c7004000d700c00440c00c00030000000c41c00c0500cc0000000700c00c1000100300000400000000000c50040000040100000044000000000000c000c00040041000000007000140014f04100000005000304030010004070000700040300c1d044400c00003f0003004000000504003010c300000104000c4400c00310cc00cc000000040c0440700c00404000f0030c170043400000000cc3c1ccdc0c00000000100000040001f000705000430000c000000010c00000000344000c0c000053303000000000cc1c040400000c0003004000000004c004110c004000000c1cc000040000000000c010c00c000000040000340001500c0414105c50700c010c0c530000030070100300c4400c00010700c0045c4c030c001c0030c40f04c3ccc00000700000000000030044003000015404cc7144c0c40004000000000030000000cc00cc00505c0c40c00c0000314000c0c0007504004cd3000c004400000c005000000040000c0d000000004001000010c04f000300000100c30c0050000c30000000400c000110040000ccc00000c30f0040300070040004c000040000005100700c04003400000330040000c0300000001000040c0c00034d000d0c0d040c00000000c001040000031c00000033c00cd04000000c00000000c0000010000f0cc03c301100030004040c000430c0000400300c0000c0c0c040000000c10001000000000000d000c30cc000010001c0017cc000c40074001001004c00000001c30c01010000c0030000c400454001000000c300004040000c00030000c0000040c04c303030cc000030c043104400c400000000000001004440c4ccfc30404000c00301000c00403400000004400c340005000c3000045040000300001c10003014405043cc0000000c0c00400014c0c0050000f040c01040000c0450c4101000c00000c40010004000c4000040107c004c00010000c04040400400000f00d0004001000400000010000c1440000003011404441000c00cc04334c000300000c00000000000000000c00cfc0c3c30c000c000054001300000000c0040004cc04004c00c1000d31c000004040000;
rom_uints[973] = 8192'h10c0000000304003001000300000c00100000040000013000004101f000010000000140030100030350000c00000337030103d000000103000c00004c00103000330c030000040000001f0001000030110c0111c00c000004000000000f01c000140c40400000403404c01c00303007000040030c031050000c00cf0041c000c15000000000000d00000010010010000030000000000330004000000040000000010101f00c30f0500000c1c10c0010c0003301000010000c00401c033000003c11000400000300000000000300000000400000000305107004000001050000100000003c01140000c0041000cc00110c0d400000100000000c000000000000701033ccc31000c00004000c0c0003c040030400300000113d11000010307040000f3000400000170000000c000000043040700f011133700001004c0100000001000f00000000000000030331010000003400000000000c03c0c00100001303000503101c00043c000700000034c000000000033031401000c000cf1300000040000001c0c1000c0f10000504303c0100000030000010000413040000000000000300000d00100000400d40c4030d330014110007f0004cd3104000001c000001400041dc0d0050000003010000c0030c000300000000503004340c03000103f0040104010040cc0030303000c000000001033000000010c5030400c101000cc4cd000000c000001c1c000010c100000c00003001c035100030000000000c007000041c01131c00000cc750001c401c00d3100003770000400031000100111c40000001c0000000300c30500000000100100c030041c00000000c1010000300300100111c4000c3040030004c00030301000c00300c3000050001000003000003010c31000000004001c40704000000100004001f700000007000000c0000001c01000000c030033131004030100100443c01340100100003000001003c30040013000c0000004000c000300000004400000004031001c0c0000033030000101100c300104000400030133300c4000130000133333000000000c0001001003c01c3000c001c011c00000143000c1003100013001010c00c03007001031000011010000cc3f00cc00000000030003043000c0000000d00c010300330033000301003cc04030330000000000000000100010000000004010f000c01100000000003c000100400001100000001003001030004001040010f03000000000ccc4003030304700000c0100100c04030410100003403011010d300000010000000003100110000000000050000010034300000000c000130000c0010031d0000c3c0500404030030c0300c0410070300030003000c4dc400000001010003004000001c000410003d0000c0000d000f0000000044c100000000005c030c300003010400;
rom_uints[974] = 8192'hc04000000010c00140c0400350004000c0444040c000000000c1000000004000000000400c100000003000430c043d40d00043400d00044000040000010c00000000400300000000000000000000c00000f0003003c0000001004030c0001c40c01050030000000000000c00030040c000000007000000330000004044010000c00c040000c00000000000001300000000400040000000c030000000030001004000010000334c0000000401c040400000010c0000040000000c000000000000030300011000004040010004000001300010c0c1004011c0000000000000004000430000404100003040000001030000401040c0000300400000000100d00010031000414330c001000000c01000004001c00100400f10000c0000c0c00000400c4740000003000040003000400c00000100000c00000340c0000000000c00400c4003030c40400000c0400000040000c010010000100c410100c107c04000c00000040040030000010000c00110c043000000c000000c000043000003c0c000c0c10c400003000000000000c0000c0000000000000013000000000100000000100301500000000440005100004400000004000400030014000030000030040030c0003100000003043c40000000034003300000000003000340004000000000030000c1001000014c0d0113403000005000c000003100c0c000000000030001000000c000f0000000300030c04400f003004040000000004330c000c00300044103c0000000000300000c00000c037004430000000007030c1300010040c300000001004001c10000500000030000c403c00040000000000000011000000300c00500010d010000000000000400000000c040000330030001c00c004000000000000400c00040000003c300100000000043c1400000140c000000000f004000c00040c0000040000f0cc0c0001300010000000000000000000000010000000000000300000000c33000000000400400001c50c0c0c001300100000400c3010000000300044000000000040000c00000101300034010000033004040c400004004c000cc00010000000004000001000030000730000004100001c00003000000300400000100404000410043000000000004103000400400000040100000300c0000000030c300000000c000040000000000000100c0000000054000400000040f430101000000400440000034000440404010030041000000000000000000000100000000000cc0030101500000c0300000000041000000c000000000000000c00001c0c00001c000c000004000000000000000004000000303000000003000000000010040000c000000100000000001000100404000000004000100400000000300c0000000030114000300000000000cc040400000310004004f00000000;
rom_uints[975] = 8192'hc030c000cfd00500cc03cc011000044000000003c000030003003004c4010100c0c7050400c00100c1400040030030030033004300000f7040c0c00540034000c0044001c00101100001000c0000c040000004c04000f34003000300034000000d47030000000043cc13000d400307000c031000000331030040010301c705c00304ccc30300010007c300004100470f10300c000000c300010030131340cf310f404300410c44414307004000000003010104000000557003c00133cf030303400103c0c000cc41010000030001004000c000c00030004043c000003330000f0dc0c0030341000001c00134000c43cc00c0f1000100000f40c0040301c001c3000cc1034110100043003000c400040330c100d0000301000cc0030131733040000000040300000441ccc0c70000c300044c03050400000003030000040100c440434dd0004004001000c0434041c110030300030304000041440000c0c0c0cc0500410400030f040040c404000c00004037000c0c0cc403c1c30703000fc004c0f000403030000000404033000f07040000031103030000000000004007000101d1c00d004040c30301404007007c00000000304c034040010340030100004103000740000c0c4043c1000100c3000f11410300000f1043000100000001c3000c0101c40003044003133c030040000047c303414103401cc1030007030000c040c0c0030300c4000041c4004440c3030400c30043c13144000000010100000300c3004001d1c3100073f1000500440303c043000000000043000003000c4343000005c00300c00000030c0003000c000000400005d40103000440000300cc4c440301c54331430f03c30000c00073000040c50307c10013cc001401431000c0003300c3000071000c400300300c0000c34dd403000d00030400400300c0431000040043c143d400030000d540410000430c010000034000c04cc0c30440003400000100000c0c004000003044000c00c10301f000c0c0000403000040031343000011c1400303400001000003c3c0030000c300c000030c000c04c040c1000300010000c0d001d34000004001cd01004003000001110300010500030000c0c1050000004001440003000000010700044003c1000c400741000100d000c004030400c0444000000144000103040000040001003c00300105410000000cf00f00004400c3c1040704030001ccc0cf0004031403010300c00301030000000003c1004303470041d00340c40040010004330000004501010003c0c530000000000f0100000040050c4044c3300000040c000045c1cd4003000c41013003000100400043c340c3400430010040004cc10300000011000003400c00400301400f10c00c44400000010c0dccccc04c0004404340c0000000030303004000400000030;
rom_uints[976] = 8192'h30000000004c01000400000f0300400004000000c401050000000000030005400c004000000007000470000f000004c004000003300400070c0f0133010000000f01104f0000000001000401300c030c0c0c4c01c301c10300001f000c04000c000c0c0000000000030003000c00000305c00003400c0c00000000044c0103000001000101c00010000f0000040004c3000100030000000000010c0404c40c031004010001000300000035000103000100050f030005000104000c0131000c430304000000000d0305c000010c000f000000010400010c0007000400c404010100000c030000000d000000c005050400000c0103000c000004040005000004030000004001130400c000c0100000300330cc000c0f000c000d310303010c010100400c000000010c000100040c000c0c00c4000001000000c000000000c00301c1000404030000000000000000010505c00000030003000c05c405c000010f000c0000004c00000400c000070c000000c005000c0004000c0000010103000c0c50c00f04000003000300010c0000000c00000000000000300c00003001000000004d0000c10c400003000100000300000501c1400f0c0d00030100000005000401c00001c00d0005000d070100000003030000010005030c00300400030001030000cc4000000c010c0305000000000c0001cf00040000000c0000000c000000c100000c0003c000001f0c0d00000004000c000f01000d00030c010400030c0f010100000001000000c0000c4f000140000c0000000000000014cc4c0000000500040c0c030031000340000f00040c010404340300050000c004000f03000303000000050140000dc40000030004030000031000000f00430d04410000400f000c3514010000000003410003030110000c0c004c0301010000030000000c030c0c010f0300c0030c00040000000000400001000d0cc4000300033000430703c001000f00c1000000000000000000040400030000014f000d0000030f0304030f00000f0001010140000c0303040500040f0001030000000003000f034000040005050100000001010000004c030c040c00000001134004300330c00001000c400f0400000403010f0000000c000001030003010004004400040c000c00030c000040000000040000050004000100001000c3cc010103000fc00040000001000000000401c500004c00000000010300030f001f0100c04000040300040400000303040304000300010004001d0004000000030001030cc1000004c000040000000304010400000114000101000100000300030000c1000c01010301000c041000000507000c040f000007030f0101000700010001000100500305040005410c4f00050c00050304000000000c0404000001000000030000050011010004000000;
rom_uints[977] = 8192'hf0000000d0004000103010303031400300101030400000004040000110100030140070007000001040000000303000001000000010000050004001500c000000014100005000c000045010c000c00000105033d0504100000000c000d0000000c0f00000000000c0103000d0c4c010104000c000000140105004c000700000f03430c001100040000000300000f010010000000000403014003000d000400000d070300000100070003010041003c000400000000000100000000000100004000030000010010030000030c00000000000c010000000000000c03010c03030c000003000000000100000d033c00000005000d004000000d000107010000030100010700000003100c0d000300040000040000000d4c01070001050c4003c1030103000401010100000031c40701000104000004000100000003300400040014054c0d0c300400c04c000d030400010000030000100c040301031003070003010000004003030105000100030c0000000000000101000000034f003c0d0f030f00000405040f000000000401000c0005003c0c00000c00040401000400010000030504000010030c0000040c4101000c000001040c004003401d0300103000000101030001000c00170300330001033c4300000c540fcf04cc030f1003cc01000c0504004c050307cf050d01000104000c0d000403000c00100000040c0107010101110c0f0004000003004f10000c0000070c040105100c0101300c03010305c000030000000100040d000c00450000000d000f040c000100300000004c07000003000701000400c0010c040303030c0f000003000f0000370500070340050d0001030000010301030cc70c03114d0c010f0101000301c4010c000001300300000f010c030107000701000f0000010300070400050005000c0000030001000000030d000401010003c0c10401000700030f07000f0003070c030300000001010f1d0000000004010000000304000300000003010d0000330c1103000d000400000d000104000f030c00003103000000000050000101003d040003010300000f0f0003030f000c000c0cd10000000f010c0d00030000030111030440000400000d00000d0401000100010430000300010404000000000d0f0103000101040400070010000300040001000307000000000c03000c00000501310300000303010d0000c7030300d1000c010010000001030c00000100010001010c000101310301031300030000030c000100010401030003070f00070003000c0501000000010101050100000510030c0001030000000000030035000003010000000c0f110030010301040c030301000c40000300004000070000030003000c010707030303040c04000703040107004100000f040c0003010107000f0fc404040000010c00;
rom_uints[978] = 8192'hcc0c01300c30030401fc0c011300300c000000010c0000c0000000344050300000043430030000000010140100000000370c00000f70100130100000000000040c04041c000d0000300000001000001c0c0000430034040c001000000003000104400c00100030040f0000101303304304073c0000340700000100403c004000f000030710000c000400001400000400000300000c003011100c00330f000c000000303000370c001403100f371007c0003d004003001f10040c0304000303301d0001000c04c0100f0031f0300400100001ccc000c4010030000100300000000c000300300010000c041c7050c40c07140405330d1004100000000030000011fc00000001010c03111c00000000000403503d0400043c0c0070003c0003041400fcc000303310030031310030000500034003040400000c0404004dc004000000040c04041c00037c10004c30fd003c010f000cc4001c4f00031d1d031c01f00301d000110010330010c004003104000c044007f000043310103300000131053cf4030314000c0cc0110104040c0dc40000030c05000c000030340000000003143004101034000000000370034010000c0c04010c1004040d000c0f0c00040c0100000010300c100c0c000c0c0c07100030001c0c0c0c0300001300030300000100401400100f003c1f3040c330030040033f100000003dfc04300700000c101343040cdc1004040c010d0103101c0c1c0c10030100300133330130f303c0000000101c30000700000c000c3c0c00000c00100c10040c0133003c000001f710040c11c0000c300010070431001500000c400000000000000c000001000c000f01000c03740c00030c01c01c003000004c004310007304300df1300300301300041ccf0030004000043c3000103c000f1d540330430010c00000c0031000000700070400001f300cc0310030000000410c010c0030030043100c000400000c1015001010000000003c0004000ccc0104001034c005140c140007040000300000f0010000400000100c10141c300130340000c4140010000000000c01000003003c000000c00000030000001003011d0000000000140c37030004300d3400043c0100000f000000400f34010004170000001401d40105030c10c0430000000c3000303c000130003c0000341c00130300040c11cc04040303004030000c013000001f00000030030c1110301c000100c100c000000000700034000003100030c010101030000003000c070000013d0c0104000c010f0c1300f007400c100304010110011503005c0010000130c004050004010c05100003000014000c003c700101000000340500140c00000030000001040010000300041f00cc04100000030304c30030300c073c0510c100003f000110cc031000303f43030300370000103;
rom_uints[979] = 8192'h340000300c0010000400300000040c00000504f0043c000000033d040c3000044c7dcc03d004c00050000000005004330c0100400d4530044c040c501c30300001c100000004143000040ffc10cc0040001c353000100705f0010004300003003c4c7140000000c40cc004300000040340347c00400c340d00d43d0c100010c000400c000000100130000730053d00400c300000700c0430000c0d0c10144000301c101710340100343010c0003070c01c100004040c043c3c0c0700003000700c1010043c140000100c4304040017340400000cd0100003040004044030034c0c041504000c1407340c40100c030d030004f003400d043030040030041c0d001000003000104034700c000c00000003f40003003d340f1cc000140300700c10301003c1000c3c10d0c00c03041c00d41c01071410300c0000300303000c04c0cc07000140c000000014c00c0000000c0100030cd00f4174300cc0004000103700044c50305c10140004040033500c0c0d0000f037100000fcf300300034000315000cc030500000003000c0000c40c004310d0003000cc3c0000c1c14003f303000040000011030051c100d3cc4330c040030007d0d00040034000c00003030f0c4100011047c13500000400d000107000c3430010030040000040d40c4f030cf13000c3c0c100d0c0d3c040c1c15c03c004044100c0430c00c0003c030c000000f0c0004dc1005401c147c401c047000100c00cc150034013300c03cc0001c10f00c0c500d300300000d00000c000c7c43003000dd0c003010000000000c01000013401c0440353000f40004000c003cc0c01013001c044010004304c4040054000d0cc003543d1c00043001000000040d7030105000100c000411000c00341140700300031c0003c03c04000c0c1f3400144440040100cc3010fc010c040d100400110c300337300f1c10301d701c04c41410000400f00734d1300404c0043d100010003033341000004f030001040040040434007010c00c3003ccfc500004c5073c1000c00040003013003300000fc4f10100100030013d044c143c1c300c000c0010304cf03041300c1404003004310c0d04314400030340c0031cd300340004140c40140100000400d00404004c440c3570340540000c0000fc5c033c101c44c4d043505074000c0f0400001300151c370c017004504005170431070d3d1cc070dc043004403003000410001c00430410043033003004013300340447000c00040400073c0c014c50100400000004440c54100cf40cc0010100040004301030440003004c0003301000043001300f10000c0000043cc004003000000000001007fc3c10c00470341f100c001000100004100c000400341033d00c14070d000c00770c070f303c04703c044130040000400c3c444d0c03000015300;
rom_uints[980] = 8192'hc3f000000c0c0010c4000cc000c000c331040000000001000030100000000400004c0000000c0000001004004000c01344000001010010050000c01040040000001000000000000c0000100013003000004400100350c0740010700000d001c000c4c0c4d30040000050340100000000000100050000c3040000f00104fc00000303000c104c00000000004030400c000400000000130c0000040c0300003d0000053000040c440300000000003000c30000040000000cc100c000000f401000040100000040130400c000100000103000c0030000c00004c310c0000c340000c0140c00c070000c000c0000300c040001400d0300c000100000000c400c300000100c03c40400c100143c3503000001147104310000001c0c0f000f004030c100000000000000f000c00030330000004400c047300c000000000000000300013010301c00c00430303410144304400031c003c10030010c01c0cc3401cc00c00c04000553d03440c0350c30010000000000440c400c4c000000000000340c00003100100034000030040400000300000c0000000000301000cc144000c0001400d00c00c000000300000c7000c0140c00004c100004f00050407003c0100c000100030040000040040310000000001c0300c00100000cc0000000013400c01000000110c010000100040054c000000001004030f001000c0010000c010000003100c00c441400000004001400c10cc400000c00d4400001045001040030300400011000000c3c1f000000500f0000000cc0000030c0100000000303c10000400000000c00000000000c0004300000d00010c00000010000040c00000c3003300500300cf10100000000030f000030c010010c10003000530c40000000000000740045000000003004c300000c0004110000c10300000000000300000f0c04004501004030cc4030300000000700440000340c0000000004cc000c0c0300000d0000000330000005040000c30004400c0030000000030003cc00000717004f300000131070004005001c00444000000000000010000c44000000c0cc1400100004000c000c000ccf100000000450001300000400001040c04435044000000c103110000003440003400044000000c0000004304c00000000000010004030c00410130000c0000000000030c0c4c00001300000d0c100101031000c00003cf1c00030f001cc04000c0c00000c500004000000c73c0000000001430030300000043000003000000000540c04000040101030040f0000cc00003f01c0400010003c0301040c00010c05000000300000c0c40003c0003000401000100c00443041010000cc410030140010000030000000c004c00000000c03f03000000000d0000c00c0000000000000004c0000340000004c000003004034000300000000300400;
rom_uints[981] = 8192'h43c04000c0c4700c4040000c0400cf0c000000000004000c03c001000cc0404400c1cd10047004000441404000c0010300400110c0410150010001010000c000004c01004040005040030000c001cc3040c5040003407000400311c0000d001c0d0c0407c001000500c0004cf00314050c040d41c0030c000c10101150c0010044000304430001c000000000004000c30000c00004c00044cc0c0043000c0100300400c0041000040100c047c4d0f0000000d0000c400c00000d004303000000c03000c0000040100000000040c10000000010c00003c4000c00cc0101c0074c400003c050c040c1c350000301c403cc00f0c100000004004000c0c000000000f30dc00001cc030003000000104040c5dcc4000041000003c4440300430cc00d010cc0000cccc00004404140000040000373000104c0000cc0c34401404d010c0000c471c1104000010cc1c04040000c3c0300f5cc1cc1f000c3334000000110040305010001c30c00c043030000f0100041000003c3000c000003c00000cc0400010c0cc104c00dc0000c01c1c40cf10000c0c0c00c4300030050c300c00000054f0000c301000ccf0000350153000300000010404c0cc41354134000000f0cc00c400f0000000043c400c030cc0403d370400003c3000100000c0001c001000c0405030400cc000cfc004c004000000001c000c13301c100c010c3c00000300040014100400d00000401c100c14fc0c0d0c41103040030050000f40140000c07340f000100c01000047040cc00c0000104c000cdf00000030004400001033040000dccc00400000011c00140000300473c400000010300ccc000c00001c0004001000c70c00740000c000040414411c000c000c0c00140414000c000c000c00300004c00011000004000004041000000c0c101000000400001c000c04000c40100114cc00040013300c3d100000dc00cf3400003c00114c0c00404430000045400000000000000030001400000070001ccc140c400c001c4000100470c3cc000004404000047c000014040c030cc0c00c1011c4c000000000d0111ccc00007070300030103c4040000010400000c010c030000c00000c4400040034cc04044000cc003c40000c00c00044300c500c0c04403400dc0400c0cc0c000040d300700c00c01c0c0c000001001c443c0c000074cccc40100010d4000000004c00005c0004340c07003c10001000f4103c140010100010c000f00010001000044440000c0c300c0c004c4030d070cc00000010cccf000030fc00d0c0040fcc0100003010000f1000c070000400000000000000100c1c040000000000040000400400504c00f400401404500010d000340040100c0c0000004400007400c4c3000c0000003c00300004d400c0d00c00400000041c0cc000000000d000300c40004410;
rom_uints[982] = 8192'h53003000401001033003d0003000f01000001000c0c3d000c000003000c031000040304000000003303171c0000300001040c0301000c0d0400310033000c030400110000000005040003000f000300000c0410311030100000100c0001370400030d0c0d000c010411030c013104053000050030373c030401000101011003030c010000000c04040000100f0011131c0d0004000f000100100c101c01000c040c040003000307010300000d3003070004000400041001001000130100001000000304000030030c050103000130000003050003111403041000130401000c0003000100000300041100300030300c0001100000030000001c103000000c100c0c0c00071004000f0c3000000401003100001f300c03100003011434010000073c0000170c0030003004030304001000050100040000000000010005043f00000300140c040500030c001300001311000c003c0c04100003000301000d3003000403000f0c1013000d04050000000000300001100f011700c115000300000f0431030c0000010c0013000c143000310000030000001300340100030010010000013000010410010111000417001c01010334030014000300000000010c0103000430001f00000d00110f000300030c1400000c00330c300003000500000500000101030000033f141f0000003c0105010f0010000300150c3c040003001031000000000c1f000000000303000c010f30030f003400340000001f03033f00003c000d11000410130000340c04133003000c1001000c1c0000100000000033100d040003000403300c3005113001050100000000000403010f30000030000014010000003f3030000100010c0000000030000f030c1011040000000000040301040f0000030330140303050104000d30030f010400010c04000400000000001000033000001033100000000003000000310001001400000700043005001504003014110100000c0c0f0100070103000c03030c3f0104010035040d3f0004031003000c00000f330c00301300003000040c040300003700000c0001030c030c00100d35041d041c100c000101033c00000c10000c00000003100f03030d000010110000100003010034340300000c110000111c0000000001100500010007000301300000301c000001000000300c050100050c070f05000034030300000003010c10000000000010030304130004300000000005050f0c30000700073110111004000000030003000f00300000000f0330070c31333c0c00100037300c0100311c04030c0001030d3f07000f070300030014000005000101010000003c0030000003000000010330300c0000013000030000003004010000010700300c03001c00011000000d010000033f13000030000c0000000000070f100d0c0100040003;
rom_uints[983] = 8192'h4c4000400d40000000030000c000004000000f0000000000000400000000c401000c000000c500034c00000400000004c30004400fc1100403000300000001d4001c00030100c101040000040003000000030000030001000301c400c0000104000000000c07c1000304104140c00005000000c1000100c1004c000c304d0040000000030000000c01014003c04000000000004300010000c40c0c004fc30f00004c0c000100000000c100010000000000000305c000010003040700c0c00000c0004131400f000000c0030400010c00040000c300000000000c004001000000500c0040004c0000010c0000010000c4030000040c0000430000000c00c00000000cc00104000103000000c003c40000000701041040000c000c00000001000000040000004c00000000c000030000000000400c0000410003000404c001000cccc00c0003030403140344030c040300004103f003c4000000c100c300001000d4000303c1070f040000c3010340000000000c0c3003010c000000030c40c00000000c0004c00000000000cf0000c7d3400004000f4034034040000000c100010000d0000043000000000001000301c0cc04040310040f0000004000000100c10cc300030000010c000031000000040400c0010f0004000000004304030340050004040103c4c00700c1000044c400030130000300000000c03400000040000001074f0003030100c1030c0404000000010004000000043000000000000300000c0000d00000c0040401d00140d104000003000100400f400000000c0300c04000000301c4000c0c00004c00000000014000c003c0000401c103004003000141c0010000000000000400000504c00005000000000001000040010003000300c00000011d00c0c00001c1000040100fc0444301400000040031000100000301000000c00700000303c40400c1400300000f030000c000000001034040000000c0400000000300000003c0301300000000000000c00100c01300410000000000000c00000000000403000d0003c100000040c0c00004000001c0c0310c000000000f0000c005000114c0050304c00004000001300003000303100000004c00030000c4430000000003000100000004d04f000f000c0403c1c003000400410400000000000000000cc050c40040000c0000044001c000304c01000c000000030001030c000004c001c00000000003000400000c4501400300010003400040c100030000000004000001d0000100000403c000010000040003000330000c00c000040000000000010000000301c000c00f040c0000000004000004cc000000c4010300c0001500c0000000000000000c0000010000000000000000000000004300004c000000000000c40c00c1c0f1000000000003000000000003000003;
rom_uints[984] = 8192'h400000044000000000000d0000470300000103000400000000c004000010000003034000300001001000000004000100000000100003000000000100000000050000010c00000000000300c00300000050000000000000cc070100000c0401030c00140000000403000c0c000300000003051000000000030000000000000000c7000030000000000000000000000000000000000400000004000c100000000d0000400400000000000000030003c003000c00030c0303c0000000c005000c0300010c00000000000000400fc50400070000000400000000000003cc000404000300000c00000c0401030744000304100000000c000100c0000c0000000d0000000000030c0010000300000000000001010010c0034001000003000d400c00000000000004030000000000000c000400000043000000000c00000001000000000000030f040000000000cc040000000000000400000d01000c000c00000100000000010400040000130000000c03400000000003000c00047700040000000000000c0000000000000000040000000300000000000300000001010300000c00040c040000040000000100000001000000030107c000000530000000000400c30c00000c0c000050c0440000400300000000000c03000003000c00040401000000000004000001400000010c4010050000004000c00000040000000000000143000004000000000003030c0310310d0011c004000304000000010003040400000f004000070c30300000010f0000040c044304000440040004000001000301000000cc0004000000400305c000000c0001000000010300000c000303000c07040c0001000d00000000000000000003000000000003000400000100001000c104013000000c000400030000000c041000030c0300000000000003000d3400000000000300000004030c0c00400400000100000c0000040003000c0100000000000004c00700070004010c030000000100000001000000000004000000070000030000000000000400000000000000010000000c040000000400000c00010004000500000000400400000304000100010003000401000310010040000000000c000c0000000030044000040000000000030100040000000000450000000003000000000f00000400000700000300000000000000c10000010c07030000000c00000001010c053000000c030000000c04050300000c000301030c0003c00000000000010400000c0041c00040000c0000c00000000000c00003c00c3c000000000000000000000103000000c0000000001000000004000000000301000000030040000001000000010000000404000000300d000003000003000000010000c000000300000000070f00031000000cc31000000c00000004000c000d03030000040;
rom_uints[985] = 8192'hd03c0000000cc0c00300000c0003c403401000c00004100000434000c0300c000000000c0004000001000040400100000400000000cc5d00330000000000000000000410000000c0000101c040010c000c0000d440410007000030004100003c103c000f3c440040c003300344c000d00000000000000044000004000010430070000c1c14000c30040000000003003003004000000000040140040004000053000000000000303000001000c04000000dcc300000c101c0030c01000400100400000300000140041040040000000c4000300400c000000004000c3134c000c0001000000340030004000140c00070004000f00c00000044400000c0000000054010ccc0000001004000004000c0000043004cc000044000400040340000010c34000003000004010cc01000c0c04c300c00100c0007004c00000000c000000040050101010000003000001000000fc0440000040c0300000000400cc40040000c15410050000040c0013cf00000440004c000c400700040003c0c0100000300c0c410041000400340000001f000434000000440000c00000000000d0004004014d0300c4011000000400c30040d03010370000000000104000431400f030c0d00040000400000401330000c000c00cc0c00000030304004040dcc000c010410000d0310041010d40010004c0300004cd00300100004004403000004001000c44030470000000c00007c0c0540000000300d0400000404000740d0000000030000000140400c04000c00001c1c000c00040c1003000c0010010c4000c4000c000000000400000000000040c0430440000c1000044003100c70c00000000000440110000003000c1400000404000000d00001000703010cc000f00003030003400d0c04100c010c37404000000017001ccc30c0300440003000000001400404cc5000000c0c440100003053c000c003000004003c00000000000300d00100000501010040000000100f0001c004400000000403c0000400410100044000c3004000040005000000000c000000000000000c0004d1000000000000000443000000100100000c000c0000000400030c0404100004000003004300cc4004000c00d000000c00000040000400cc00000000040c0c300034000000030004c030fc0c100c0c000033c3000c00103000404cc00000030d0004000040000400000f3400d00000f00440c000000d4fcc0c000404000000000c0433d0103000000400001c00010f00000000f00453000c100c0000010cd00c00034040030001000d4300040410cc0c100000100040100040010d0000014000d100000c00040000044003c00400c0f00004000004000003c0000000400000010000000c004cc0c00003c003c0300c03000440005c05400c300c07000040cc000000d40c40400004100001000;
rom_uints[986] = 8192'h100000001400010c3010000405131000001440040f500000303000c10c001000130100133010000510003c1000103f0c30000001300010300c0000001c10001003000004c000000000003f0001030c003c70030f300013000000100001040000340d40100303031f00000003d0010100001010053014000010005440007c3f100000130c3000000c000000c0040000040000000014000011030300003f03001104000031dc0cf70d0400003c0004000133000000000041301144033c04500000c03400000400500000310000001010d10c00001300000300c0010000000001000003014000300c03c0000044d00c00411000c0400014100013300c000004c0510011001003004300000cc014300030100430000d05100c3c0010301030540010300000300410133c41000d000030000d04101c00300000330c010003f0300030001cf03437c0000001053000c0000f300030000c0fc13400303000341007034034100000043330304c00100c1000c00310700f300010300311110500001034c000003c0000003015101000101c1410d0000000300c000040004c30041c004747003c33300011000300017133305000130d40c0300c1050d00cc00014c10000001005033000001030c000110001040010300503013000000000000000001000000040000451414c0f313010c1030330c00cc00000000310003300300001141000003cc0011300000000010c33031100003000050c0040000000000c70c0000004000003040c0330004c300000300100000c1c0313100410401000000000000000403c3000000100011330100c04000010c04010043c03013410000100003003403000043000300c00071300003c3110300c0033103004c00c0001003003001004001c0dc300033c0000fc00003000410d3c0d300c00500000000030d300700400100000003073000c070300031000001f4c0010000011033000d40014000000001010100000001000003003103003101cc0100040100134100000001010341300030730100000100044033cc003c0310000fd04070031001003010333000000101000d30530004010007013013303000034c000c40000040c3030000400030000000001cc0300013000000100030000001c040010d0003414010f0000000030013030301000100704c000003003000c040404400010400c0100f00430f00000100034330000000031013035300c00ccc01000c0300c0000d0c00c001ff00000000c000300003100000034404033003c030330040334300010c4703445000c04101100000031000c01000c03030030000c100004000104400000000c000c3100100c0040301400000010000300cc3000000030310340103004310c045000100c00000c30030003040000300001c13034100100300000d13f3f10000000000c0;
rom_uints[987] = 8192'hcd4000300d0444000d040004000000000041000000100c04000c01c00c3f000403000000000000c04000003000003044c100000ccd0c0000000043f0000c003c0000000000000c000c1010043000001cdc1c000000000000000c003000000cc00734c30030040004000010404000041000000c0c0401010000041104000000000004000040000011104400000000c000001100100004043434cc00c1000000000400000c3000000000003c0400000000300400300700000000c0030c00003000044000003c0c444400010400000000003c0000003fc400400000000010003400010304cc000f0f00101017000000000000400c1000000c000130000004044c100c00000000100000101fc00130000000dc0004000cc300010000000000001000000000300000000300000010040000c000100400c000040400033f303010c400000c00000000000c0c4100000033000c1c030cc40c000c00000010000500000c000d3040000c0c000000100c0ccc00010004040c3000000c00040000004004000c101c03c4000300000000014000001000d0000c0001001004f70c0030400c0004100000300400000cdc1cd00c004c1144100d000403070f3c3034103c0c00000c0004000c000004000c0d100010110003c040040c00040000000c0030000c1007000000100000304000000c0c0c0001330310001004000c0000000000c40000000040000000000c0c000004dc000000000310400004000000c10c0c010400000000c0040cc0000c04414c0300413000000404000000401c00130c00000c0003004000043c0000c000cc00000404000000700c000c000430004f0003100c0c000001000000000c0c040c170000c10004c043000c04000000000000c00c0000000c030c040000370f040c400004c0000100c41000fc003000100c050003340cc00000c00c0000000c0c1c00000000000040000f000000000004040004000000000c000000000c000000401c00c00003001c0400000c3300c000003404030010450c0000004014000400030304010c00000000040000000c00000000100d011015f00000010cc00000030000100400c010000c100f00040c04050000040300d4040c01300433030d300040c1400f0001000c00cf30004000cc04c000000034000010000c0001c00040000000000c07000000000000040000350000001300c005c030000000000400003000001434030040000000004004010003003c110c0030000303000400004040030000004040000430000c00c0000000310c0f4c3004003000000000000000000000000004000000000004000c003f000010000c00003cc00400040004f00000001000c40000010503c3400000000030003004005c00000000c00c0070000c0000000000000c0cc00010000400000000;
rom_uints[988] = 8192'h304010000100ccc100010c0f5037030053000004000fc0000000300003000303000cc0f7c3004110001000c00105000c1000000000300014100c000003001300001047c3110110000c00303413030310030c000000cf304010000c1c010003031003370f0c00d01c1130030030003001000440c300041333c03031d014000f0c10400d00000c0c00030000d0001000000c000000000000400003f04340470030110010300100400000003000c1000c0000f1d001000001c0400c0007c000c00300f0c00d00000300c01000414000110c3000300c10d03000010c01130331001c000100001030000000cd00477003300c3330030c00d0000000000031103000013040300131000c011301f10301000010c13450000041c3000cc0303d0004300101003c00031430303000131000c4000000000404c001100000300001cdc007d007000100100704000000c0040343011114000711d004cc1c13c3300313341f43410530001f03c400c0000c30043140c103010c100031000000c0030c030000000001cc3403c01003435000011501300c34000000000103010130000f313c003000cf0034c4c00030030130c00104130013004c04100000730111401341000000303000400303c0035031c00114c304c570710334103313c330000003003000010000c010c131000000130503000000004000340313000003310100000c00010000000000111f000004001000c7f011c030041101340001f0130c1340110307403003030000070c03000000000300300300f3000f10c1d3c0000101000000ccc310310000300013300731004c00000130435000100115030000cd33f3300004cc5040000033301330010f03305400430c73000003001f040d1c110c300000000100340d00000c00030d30000d3100c000001031c00031000100c4300130c134300003130000000c033c31cd011410100301300034000003100300f73010300100031001010000030310040015300310cc000301113400000300400007400103030c001c310401100c3031135001410011f0010c000030d0030000000030000400733000030c0f301c1303340000c300330c00030100034000501340cc000000005301300031000c040030c01c010003010000130103701000001d011000001303043301030010c10000c30304370301001001c441037d001300100000c030c700010310043c1d003034100710c3003d00d10c000030000303000c0131700350d301f5c040030000041d1c07400011010011103000110004000fc0f4010040000030001c0d0300d040104000f00010000f00c3000000005304c10004003100031000533110c0410301010041100000100300050070340300070c04000103130c1f017103000003100fcc300313300000001300f030000d0c000c003710000110c1;
rom_uints[989] = 8192'h100000001c100000300c101010070000c000040000f04000c0000014c0c00c5000333c0030500000304000530000f050c100000000c04030001000053030000000000000000000000000000d0000000001c000000040400c003014000030003000f0310f000000c00000c0000c070010300040000c000130070010c10000000c304700104010003070000000000000000030000003000000c00010000001000004f4040430100000d0003000c031000003040000000c00000000003c1300400001c000c0000030030000000010070000000003c0011000033c00301433100030cfc0c3004000000000d0300000003c103000100000003330000003f10000000c000000300300001000000000001000000100100000000c000000000430330100000010001001010000004d00100340400000700000003000c004c004100000cc0000010000303000003000000000301010100400c030c0c0c000301003c10043004000001c40c00430c01100000000d040500000000c1010d030c0004000d00031113001003000c000f03000403040f000000010001c000000c04000000100000d503000c07000000000340004300001cc0000010000004000014000003d300130000000c0000000300700000000000000004000f13c10100000700030c0030c001000000f1015000c000c30100000c300000000f0f0c010103300013c00010130304c00c040300000300010f10000f0d0000000300000c0c0000c3000000000004c40c3d00c0040010110135030f030ccc00030c3c040c00c3040000000001010000000030000303001034530c0c000000000000010014000000400000cc010004000003310305000100c03700044004000403c1310000400c00000c703000000000004c0004000f07000505000cc000413c000100340000c4c0014000000100000044000301c0000300010000003000705000000c100003000101000000000300100003000004c400004400dc03c0000c4c0c000030000300000104000000040000304f30140000000040010001004001c0700000000000010100f400000000000010c00000030000300000300000010000730000000000030010004c10040100003000000000304000000000c00000500004000000103c0100010470040000c030c34330000000c11d730000c0040001c07004c0000000030000004000010003004f0c00000000410003000001c40101000d000c301100340003070000000300010100000300c50000300100003300030400400000000401030c03f0000c0ccc43c000010f0000000004400000030000000d430010003c040300000000000000011001110400030c000c0100004000400000000500c000030c001f00013101010000001100070004004c000000000c000c000c01030431c3400100300000;
rom_uints[990] = 8192'h4711130303001300d1030007dc000005307054100041cc0000443401c14004040330c011c010c00015c710101000110c00c10011004000dc0c11001030403c100000c0c10103007300000c403000001c004343df0c330100000c0000c000310010d13103040045d0d3d01300c030040fc000000404400401103543000300700007010034013f0c0c000c0000010000010000000000c00034d0c300000c30041113c0004c00c000000013c100c4c10c13400050100030fd0344d00000330c00030011000000100400105034030300d3c4c0cccd340c540c100f3c300140cf00d403103c010c30000470d4c0c030d4333400400c0300c0000000cd00001000000000100f0410150001310dc010c04330110404130344030003740440330000f4d0040c4500030040c000030003100030043040303413300c00740cc004145400c0301001400cc1000005004003005403c0000f0005d01101551040017000f10003301301c10c014073310d00053dc031050000010f00300733001000440000c310f0071330000004000110c013d00004000030cc00000001c00043100070340401c1d43c1c014f134000010143c03000c000c1700053410001050f03300104343044304040f40000cc00700400100c3001c0044030003d701000100004544400c00100101000c0007710413000410430030000070101140040c300d000cd04c04001400000c0473400d0c014731c0500f0cc31040001030300d1c0c0cd0411c70c0133ff310004003000041c070c00c000004000000003300030c044440f00007100d100431100030000017c100003c430004c04010137c10443004000cdc03317107033c035c000044c430034d0000301330740003070440333037000050001000300000031000003000103300cc0c3031400c3000400c004000000107104030004c1030000053c310cccf074710000004770410d00f0040c300000031130004f00030004000001101003000cc003001010d1010004130401d1c0010c07003c30d1000000cc004104000000dc004003011000d1dc000c43010040d0000141100040003310053031cc000000341300010c0c3103c010c0c3c1001c40430300403333f0004040100004007305000013c500000030010cd0c033cc034400001040400043440cc0403330040040cd74004141c34001300300000073140001400c3d0410003000f10440c4000c03c00100400044131101430c000000000010004473000000c0000000010310700d30004034c130df0400dc343004330030303040000070c0410404000103014300c0050001d100cd0c17400340f01000c00000cc0300030c0f01000113c1dc01c01004000401103131300040301001013f010c0400441430003c310000014001c330c03340c0d000443400000003300c340030000c04;
rom_uints[991] = 8192'h10000c30000010c0000000000400c00400000000300000c000000000040000005000010c0c00040404300d013c4470000000000c003000000c040300001000041c0100000400000040000400000000341400c41000f1300000040000000001001f000000000000041000c4031c10000cc000101f0004001c00040033014c010103c003070000000014c0cc100c44003000010000000300000004041c4c00c00001010001000000014004300c004f00000030000000130010000300c00400001c034000000304000c0000d4c30030c00c0c0c10100001000400040f0000c0c0000c0c013c040000c000f31c50000000330005000000000c0c0c0cc00300000004000000f1000000300c000000014c400004004000c000030100cc0c001c40000140000000004c5c00c40040400000300c03400c0c040000000040c0000000045030000c4c000c000c0040c03001000c34103cc411004304034010000000140010000034040000013c0000403c300003130400034c03040c43003c003cc140000c0404c4003c0000300000c100000c010007000000000000000400000730001340cc4c0c040000000043000c10040c300003440000000c400404000c001c00fc1000000000c0000400000c000000700c0000000c10c034004001037c00004000003004000040570000400440c000030c0000300c33c0000000001040001037000003003000000330c0010001330c301c40400101000001c400440104000f00403004010d000010000c31040c00000000003300000000c0000c00300400300003430000000c0000f0400000000000c000300000c00c300c300000c00c305004c0410000300403000000c413001304c00c0003000400401414c0040c13004400014c0000c0004000000100c01c05c0040c0000400000004c000f0004d0000400000110c00003c744cfc1400c07000500c0300000403c1015000c100010000000c00430000000c0040400100010000030000c4000470000004000001010c0c300c000f403c000000c00440400c000100d00300000030000001400d00000300000300040000000000d0700000000073c40040c0070cd00c0000444400004000014cd000000407033430110000000c0007000043340001000000040400c000c4c000010c4000101040c0c00004c0404030c00000440000c00030043000000c0040030001c00000000401030000001000000400c440c000304001c040040000030000000000000000c0c0400100c07040000000040d040000c00c40c00000010000c403407c0000000c0000000c140000100001500040c00000000000000040c043000050001c03c00000000000c0014000c044c40000c00010c0c00040300100407400c0c00000100c043000500cc3cc0003400001000000003c00000f00c000000;
rom_uints[992] = 8192'h100040000010000d050000400000c1f4300000c0400c0000007000000c437300001000d10c00000000440017c000033000000000000000d000100030300043000000c410030000000000000143000000104c10cc0000000300000040000000100000051100000000d0d0150c0400050000040001004c003000040c0070004000330000c0030f001c0c00001050c000000c300004000000000040434000c0c004d00000010004400000000400c010000300310700000000000010000033000c400445000400000403cdc000003030c0000001c40c0015000cf440000000cc00000003000430c003000004001cc01300030000000310000000000000c100540400000714110000000000400000140000000c043040000c0000410000011004c0100030010000001000000c00004100004400cc000c000000004040000140000003000000c00005000073000c4040000c400070000c00f404004040000d00004440010300c004000043000000140c000400400c000000401c00f4d00010040000c0000000000c0c000000000000130000300100004c000044000c40000000000c0010040015050000c10cc0000000c0400c000000540c140c00c1000344000100301104c0004c4c03c40000c1c00040001104040000000040000000c000014c1330030000340000400c0d4c000700300104c0000003f0003000000c000400000c100c0004010340030c0000003c0413c00000430004cd000cc0400030000004100000cc0404300000000001c30c0100014000104000040c00000c00c0410000000003f0040c000300c400c0001000c0000100000000000c00000c00000045400004000030c0f500003000000303c001030000300100003c00400000c3004000040010033000000000150000000014000c00004000c00000000000003100400c0000300010000000004000c004000000000030403700000c00340030000044040000030000400000000004c0000000000c000c00000c10000010c011104c00000c0044000cc0000000c00000001100000000000014c00003300044000001330c0400000400000cc0440c5004000040000000000004cc000c33003030004000000300000300000104000c000c00000000000000004cc00cc00c0c040001030000400047400000cc00030c001000003340010000000033400000300c0000000000033f00000005000300c0000031000000c00040000010003000040007000000000004000134004000100100000000000c03f4000c00000011000043040c304000000004c0410000c0003c000c0000004010440000c00000000c000034000000030c0c000000cc000040c50000100000040304001100000000000000040c3000004400000c00000044004000030000013c010004000043000100407300c00000000000;
rom_uints[993] = 8192'h100c000000001000000000004040001c0c003000000c00000000100040c040000000000110040000001000000000003030040c0c0000000000000030c000000000403c14340000000000040400000000000c001030c4c000f07004f00000040000004c104000000c0000300c30000010000010040040001000001c300c1000003000c010000000040000300000000c00000100000000000000100000001000000000000000000470000c40003c00005004d0000000000010000000043c000000300400000000400c40c0000430000000000400f01000000030000000c000100004000c00000c0000000c000010c0003010000c000000000000003000000400000c000000001000010010000030001030300c3000000c0d0010400000000c000000000000c00c0c1000000004000000000000000000100c0010300000303000000cc00000000010000000300400500000c03000003003000c0000d0000000000000400504000000341000000c300000000000000c0000000400007000000000000400000000100000000c00c00030340000003400100014343440c0000c10c0004004c000c010000000000410300040c00cd00030100000044c00040000cccc0000000004f0000000000c30000c0030345040004c00000c300000000c30001c0000040c1400001000000000700000c0004000300010000000c0003030000004401000c000000010000014300004000c0000000000000000000000000000000c003010703c00c000040000f0000044000010c014000c0000101c00c00400000400000000c0000000000c000044c00000005000100000000000001000001000100c701000005030000400004000740400004400010c00000040040400000c0000c000043c00300000140004000004003c00c000000030c4100c000000f4000004000c3000000000000c04c04400500000001c0c3404000c00440000740000000000d100000010000c10000000000000300000000cc00000000c700030001410001c00000400100000000000040400400000003000c03040000000000000043c0004300040003000001030400010000c003000000c000c00000000000000403010401c0010000400c00c00c0000030000c000c00001000cc0000003c400004000c0004000000000c00001c00c00050000400c00004040010000c0004040000000000c000c0100030004040000000c0003000300030c040303c0c140000040c04100000040000000000503410004000c000040000c0c04000000000000c0010000cc00c0000000000000000740004040000000040003014001000000000000000400c00000410003c3034000000c00000000004000004000c4010000000000030000030040000000400000010300c10f00000000c0000000004040010000000000000;
rom_uints[994] = 8192'h4000004040300000c00c0c00d000001010d000c0d014000004400000cc00004000000cc0c5f00000c0d003c03000cc00400400f010c0c000000000c000040000000030c004000000000ccc1000000000dc100010c434301400000c00000430c0000c101c100c00004c40000050000c400000013000c000c000400000c0400034300000000c000400003000c0000000000c000000000c00101400000040300000004400000c00300000c000c0400004000400f000004000c00c4004d04c0010000430c000000cc00000000000003000000000700000000000001000003c40c000f00300000000000000000010c0000040004030000000000040403400000000400c4c00c00c004010c043440040000cf03c100010305c100cc0305070000000003000c00001300c400004000cc000cc00300010500000000c00004000043000300400003000003000f010c4c01504100040401000400000c000c00000000010004400c00010000400f0103030fc400000c00000007070440070000001c00000c11050c003c040000010000000000c400000001010000030003400043c0000c00c40d0000000c0c0000030c0107c000c044000300000000010000400d0400000cc00300030c0030c10c000004010000cc14004d010000cd0d00000000000104000000000c0400004c004d0000000100300300010d004d0004040000000c043441010c0c03000000c00000000500404000004000041c04040001074300300040000f340d0000000003004040050c00c00c00c1000000010000000000000000034c0000000000430000000c0400000000040001400100004c00000041000001c0010100c30c1f10000000040dc047000c0000400c00c00c0400030403000000c000000004000c400040c00c0407c310440c0c00000c0000c401000001000d030100c04c00004c000000040001070c00430c000003010000000c000000000000000000000400000000000c04000c01004300400003000c0103010000000100004441000003c0000c0c0000300c034000040400c400c00c004000c104000f0d0c00000001040c004c0001c0000001000c00c00c030000040000c0004c404100030c44050000010d4c000c03000f0000000d040c010104000000000c00000fc0034d00c000cc0c0003010001c0400c000c01000303000d01040001404c00000c00410000000000400000f000000000400000c00c00010400000003070004030400040400c04d400c01400000074c00004010004004c0010000cc0000004f000000000000010cc00c004f1400000c0000000c03004d0400400000cc00010000000000000000c4430c03010c0f00c700400c00000000000000000004304f0300014c000000c00100010c40404000000000401000000c000303004c010c00000d05030000;
rom_uints[995] = 8192'h40c00003000000000040f14000040c34c000000003d4000144c000043034000cc00c3c00301400000404f00000140040dc00540c0c141cc074c00ccc00000034000400cc0004000000140c00040c000404ff3011000010c10c34000400cc1000344fc450040000c4c0000000100c30100c04001c001c440c00c00030344400c40400c000c00cc004000000103c00100c3c040004000c03dc0000000c10100c00d0c0000000040040344c04d0d00c040cf0000000340004300c3cdc340400001c0004000000500d34000c70c7ccc4000c040000300c4000004014440cc001300130040100400000040c00c00c0c147c100040f00030000c001010000010000c000000301400004000400cc40030040050f43530300c343c010c0cc01cd01c00004c400400000c100000ccc47c00c0cc00040004000400c00040341f04001400400c10c00440c404001000000cc0f40400040c00001410701010d4043010407430c0401470000000c014c40c0000000c00343c0ccc00c03404000010c0041001040cc00cdcc01000101000c0ccd40440100c30100004340c3c00ccc0f034d01000400c04dc00000000000c00c0c0c010100cc400c4301c144030140014f01c04dd0c0c440cc00014003c301cd0c0000c00d00c000c3044700c4004000c0030400c0001303c100c3040500000400000c10040040c00c040c4c0ccc03c0000c400100410c000000cc000c0700000000444400000330000c004003150043010000c0cc4300c3c043cd0004c00307400001c304c04040000100000001ccc000dd0d040303cc4000000101c0c00ccc4cc0c0c343004043400c00000003000000004300000300440340c70c0404044dcc104004ccc0004040cc0303c30000000000c0cd40c040414cc303c00c0304030d0c0c00004000010fc3c100404000c14000030000440c000003440c0cc317c34000c00000000c4c0c000f44c0c0033c030c4300c0000000000c004740000040000c00000003cc414f40403000c004c0004700000000040d0c00c4000010c1d0c00000c0cc0c0300c00104030040030404c10000c5c000c3074340000070000007404303c00500400370c5430000c00300030313000343414004400fc00040400c440000400151c000c1000c04000004fc040000c00000005100c000410c0140004440434340050ccc00ccc000c0c003403c40c14040cf010c000444000c704440074c04004404cfc3000041cc00000c000344010000000040cc00400005c0000f104040c3000001c005000f40c10f41040441444c0040004c003c00cc0401c000003100014003cc0003010000c000000070000c4404000f003000004fc0c04c030001000041c4000400000d000f05c0030040303c0003c30400010f410000000f000040400cc003010004040c0040c04cc300;
rom_uints[996] = 8192'h400100300c3c410001004070031070000000d000100c03000401000140104000c1000030300000014000040000107c10cd00000f0000c1f00003010000000000403c3000000000000040001400103015410c0040400301000c0f40001000400007f3540000513000103110000c0000103f304505031111003070c000030f0414c30000000000c3003300c11411d00003000004001000031010400100030000c001c300c303304000050011d000003000c030000000300f00000003030000000031033000003001030000000c03111010013000004033003300c10110c3000015000300c0030000000c041043d1000010100101000000030103000011500030100103451004000003c0c01411000000003c030003000310041010331033000001007000031000000300c01100001000000000001f001000030c03030c0100030001000031000f00000000110d00c0300300000013000c300f00100000133100000300c40000f30700c001110000c30c030c010041131000001340040310000cd003310031c000100c010000f1000313100000000000100030004044100000d10c7c33300f000033000f30000030d00c00000111400100034c110100000000300415001003c0000100cc0000c003c000300040d3010000000040000001030301c00cc30100000034c30003c14341000f0c0000c00000000010000c0001d0001000000041c005000000c03110c0cc000c0000000015000c15104f1140c010000400033c300c0010000000c01030014c4003034000010300000303034400005000000030004000030100000c01000040030000300d1300d00001003010f0c04300010000101c0000400000004c010001c14000100000000300041d30040040017001d0004c0c000000001000000000c04001c43f0401000010000010304c001000c3c340010000731000d0f03100011c010340050c0003400103300c0001000100d0000000c3000011000000011000000000000000000100000f05000370c300000100000cdf000010000c010000030c0033043c31003f000040000041010000000000001000000cc00500100040150040c0000100333000100111000500000401d4c3030043010000c0030103c10040000010c00004305000000300000000000410430030000040004c000000030c4100003000c3030400100105030033d0c00c010303cf100000001030000c1400300133003c0010331140000100c010400000007030030000c040010000d30f00110000c0030d01033400c00003000001431304d105d1301004000414c015400cc001000000000000c50c000d000000c0001c0010030003000c400101f340d00c100000003001030f003000101030004141400000100000000031c4d00c00c4c04000c03000403f40040473c0d0cc00000000;
rom_uints[997] = 8192'h3003110010000000100003003031030100303d01010400100030d000000c000000000010113300000c10001310000300040000300100030000300003030000030010030000000000000301100003130000100000f1100000000f101001100100000130010300000001031100000010000013300303000000300030c00030000000100000033000300000100100000030000003100000000303000003013013000400300001031010000100010300013001030000010000310010300030000300000000100000133130310030000f30003004003103103030001100100300000000300000133000000000030000f00033000400000430000000100000000000300033031030000030000000010031030000030010010000301c000101401000000f00000001000000010001030010000000003011000000010000411c001003000007310010003013000000043101300104030000000000030101001001030000000001130300010000310000030004100010000301000000000000100030100104301000003300333030003300001331100000000000000300131301300104000c1000100000140000310300001000000000030000300000110000330000103010000005003000000000000000000010010000000001003000100003000030103000013001000030100000000000000c10101030030000000000000300003330000003003301000000000304100000040c00000011100100001130000013f000073010000030000000001003000030000500000000110030003000000000310000000000300000310000000000300100010030033100303000030013000000000030000333100040000031130100001000300300033c3300100000001010103300300100003010003000000101030313000000100000300000000000103000010000100030030000000000033003001100000000030103300001003110000301000000000001030330000000000000000c001001300c04010113000301303003300001000000010300030000003000001000100000000010100f0000003113003100000031003130000033030f10300000000000001030000300000000133000003031001300003003000000003010000030000000000001003c100030030310001000000000000000000004000000000333033000300f0000001000000030030000000003000d11000001310004303033000000030000001f000010300003000013100000000100000000033031000700001103000000030000003003100030303001300100140001000030000013100000304c3003100100013004000000000004300c31030010000000000000000300000d000000030001000030001300100100000130000001040000000c0310000000000000040110300001000000001;
rom_uints[998] = 8192'h4300004101410c03f3300d0ccc130003c0100003100000400000c0004401f014410300343f43000434300d030003314030500130d301c3700004043000004403034c74500140010040010c11c00400000dc000315100030050350000400540057d30dd030dc000077100700044400144403700514103034003d10f00004d10033001000001700c0000510400000c11f004c10000000f001f03000d1c00414c0307c3000003000dc01130000047c00c30c0c0cc00000443100100133071404404010030c1c00c04c00c000c01300373071430404333f00140c0440110c50f0f00003000c03011000000304fd00300301004c40c0001340000040c0c00400000d310c04000400051d10100337403c000044fd00000000001c0d03000d3d30303f0003cc0013700770040300370400045337000075c4010100dc010cc00703030304131c135710f300134c000001c0304c0c1401c0353310cc10011c10400500100000011013730fcd0300531030501007103010000400300c401c350000c0450f3501450007030d0c0030344074000d0103000014100013001011030c0cc10404004503030000004004cc300c5004000030100c0540130410000310c1100c34cccc440070c0000000000d0330301c00005c000001040005300034030c000d007010100f3303c0100f04c0c0001004000533000d51003f31014543f00030c4043cf00010340c01cc04c00d031344033001041c0d0d040030303130d4000000050c00c00101300410140000440014c004c0c0140000304407001004c03d340004004004cd003300103000000540400d310040000430c0004704cc3000004c01001c300c100cc10000004410351434001000c0440f0c40d0c40c40070100d0c40f0d00cc0c000100003ccc00015410c034030c1c1040004100c70010c0030d0004543c4400100c00000004700c40cc04c07141c4300d1401400f5001713d0000300000001000c400033004f100070403000c400f0c0035403000314031140c00d0010000040d3c030034000000030440004010004453c40034004000041000c10c003004000011000d510000107100c30003400400047100000103cf000c05030c03110d0c14f13004cc00141f0c304f0500003dd5004341040000cc0074d00314dc31c00001353300c001075000c0314410003d30c000470100433300000ccc350400d1003c00000001101c00ccdc04f00300140413033c00140010000000c0000c00cc0f01c1003330000cc003003c00cc01131f000c00d00c144043c0d00105351030cf404401704300000010031003030075000403000000c01403000304130444c01400000404300430410000303000c00cc0000000010000c3030f3400000000041051f000003500c0141001000040cc0000d00004000c1044004401c04c00;
rom_uints[999] = 8192'hc00000000000100f0000000011fc000004003030003000c0ffc040033304c0300c153c01000000000000000030100133cc10000d03740c0000100f0000000000104000000030000000503000000070000040d0000030000010033014000d000c4174000403f0c0041000f000110000300000040000103000c014013010000c104030000f34000010000040104010300000100000c04000110c000000f00300003300040000d0401004040010c01d10044d0000003040000c1010cc0000000c0c000000001110040000c0c00030044400300000001000000000c03f4c00000f10000014c00000003000004000c030333434000040000000340f3400000005300400c0c000004400001030100000d0c0440050c0005130c00c0110010c0304c0c0f000c0010004000014400cc003000000001c00000000000000103c0000000000001300c10100100000041c00000c403010003015003cc30c004c00000001000030400000000010700c1100c0f01c4c0c1100000034000cc11131000040303001d0003300340000003000040000370000001001004dc0fc01000c0474000001300c0140c00033003c34300cd1000c30000000fc0001000040304c000c3ff00313000340300070003014f040005000400400300c0010304300000100003000cc00700000000cd000d0170030030040d0000f40000000300007100030000000341000ccc34c3000300313004000c04040d00000c300103400c0040000310101c0400040000c430000c010301c001c0000004000303000400004c0c04000303000040030000c3000000440f040030c04003303100c00040000040001c0300d0000000010001400403000000c0304c0003000f004001300000f030000f01f00050c000000000000100c0000004100c00303c0f0001000000010d00000000c0000701010300c401f000047000c000033500033c0040003c01f5000013110400000001001000000003000000010301c0c040000c030001030cc3130f40c000430013000030070000c30000000000f3700031c00300440013030000c30103c000000040001013c300c10cc0d404000033000300000000030000000c00c3010000004301000400030c0010300000c04030000104000003030000001c500100c103c0040000c0c00c00c0c00003000034040000f010510400410100000031000003400f0c0004440c0000040c010000300f000300001c00c0010000c0c00040430000003040000c0000c003400000500000010dc310400c100f4000c00000007000003334433330c0400430010040000101000001000300400f043004000000010330000401030f000f004000000c00000040000043000100000c10000400033000030c4000400c00300c03341001c30c300000c0000d00000c34400303f0003000400;
rom_uints[1000] = 8192'hc3000000333000050c0000c04000400010503000000f33030f00100403011100005300030100013140c10104030000d0000000010400133130000000300000300003d010403d000000000d00c0004f1003000370d111033f0c4000030000070004110000c033010033101000101011000c0c311000000010c030307000000003f30000300300000104f000000000035000c001000000001330400100d4103c0033007033100400000000100000f10001004013000000100100c00147041300c4110c03001303004000c0001300330c30003c030400030300010c00100c1000010700030003000000000003040f3350030300030031000000003c003300010033000304000300301011100040010000000f300300100010140000c000334007000c03000000130000003301000000c1000000007000040000004404003000100c1000003005110000000041131000403c0310000303400031100100113001cc0004401100d103103003010003400c1040000000330f03f000c4310031c00033030f000310110030030300033330000000300000000001d0000074000010003051c0c50010301000030c00010304003c3330110300311001130000010000000111300004010001000003033001310104000000000000040003c30030040c00301c00c0310c030410510001011000000fc4100300100030033f03033013001000330140c53300000000cc00341307103110d0003000500300044300503c000f30330c070043001103100001430400030503000000003010114000340001000031000001c3300131300010300f0000033000700003000031103011044000100013c300010c415c0010c0340300d0000014c300030003000001f000000000c01010300401011000000d0000100001d005f0010143f00000003030000300000100103300730310011001030c3d5043100300000f1000000030000103000040c0000100000000000001000000001133001000300000410040337113704000100140000f000100034011031003000404030c000000000f300c01f011003c050c000300000c30003000100000000110003300031330000330f301000001410000001c0143000000040c03130010000330030000000400110003c033000335000000410000d300000000c033000301000c131331003c0000003c300301000000001d0000c03400003d3130000d11100000000c00000030c03d000311d000d00c00000000c1c430c000100d3043110004001000000103c003133000130dc00030000300330111000c50010103110000000d30000000000030f10000701000104003000100100041c1400000c300013003304001000003031c0403000300c0000000000300330000f004403000000000100000000000000101d003000401d30010c03300000;
rom_uints[1001] = 8192'h3c5333004001007d00000030c330040003003101000000000040c0404030004300d05413d471000000300003001c0030000c30c01100f0f7000000c000010000003034340cc0100c00000770404014000030410043400000000cc7331003d0400430330313c300000001000300304cc1c000003c000310400d403130314000003011030000c000d04030001000c0f0104f0003c00000030c13000040300d0100c4c310000000c0310007000d00500030010100000000c33000000003c4400043043c00c0c000033410010040f000c50400c44100030040000000004000d000c3300303000000400000c0000f00cc00434003c7331d0000000003c14000000003330403310000001cd303ccc0004c304000d303c031001003000100f771c4100140334100004400c00041130070400c4401000000000103c00004001001000730030100030050100000c04040004000c00f004cd0010500c0c000540f30003007000044101303c10000004003110c0c30003003003100d3000010301000403400c03d031000c400000c0300001700c0c01000100000000c104100000000cc01003104000410000404000000010d15070000030041304c00530130300001c30003030000410000c0dc0c41d400d00000003003331340100300410000000310000303300143c0004100004f0c0f400c0001f400030c000c4003c000c00041300f0310000001000c0010070300000010000c7000000151000003000103430040030341c00030d01100100000300040004000003710000304c0001000d1000c00744000000c304040000004c0010001000010031330c040010000340d004010d0c1c0334431c05f001000003000013310c4010c100407c3700d000000010001c103030000f30040403113001500004000c03000043441000003c100100000c0001400c00030f07000004000030034c0000000000c03130003300040001300000000c011c00100c000044340300040100000000400d50300034100000140030000300000003000c3100c4000000100000c30000400413000003100000000010c0005001003010003410013370000c0000003330000001003000c000c300000300001f0d00c0000317c0004c1404010000400003000000001c700013301100040000001407471c330303001004000104004100030011310001cc000c001000000000330c00000c00000001000c0c010713040c001430300f000370300c00031c03000000040001c4000cd00000300c0010000000017170f14c040003000c00d00000051cd00010c00100000030000d001030040005100010000c1000000d000c000001000434001010104010000c000000030000005014100c001500d30f00013004003010010000000404c0050003700c01000034030310140c0003000000013410000;
rom_uints[1002] = 8192'h30c000005c0000c0c000f01300300014300403c003000003314c00000000000000340030031031140000000050101100cc00044000c000c05001000033340040000300000000130100040000143c00300000004c30000003000c4000005000000000100000001001030103c4041000100c00404c1f0000cc3030000014c0004010000000033000000030001000000100000000000000c010031000003000c000000000010034c0000f1300001fc100000000000100400040c0000000004000c100000040000001000033c400c0150300000000701300014010c0005001c0300100c0000010c00003000010305000003300300000000000000000103000000f1c0304040100000300000301000401333c0c30000cf00000004c4400500403d00300000cc01030000c003000000c0c4000d3100c100000000c030000300030411c01100000f0c0c54400030000c030000000000c04101c3040000001000030100c1000000000100440cc0c10000030f00000000000303030c00000f000f00c01100000300401700c00300003c3000000000000000cf010000c00f000004100c00300000400001100000003000cf1001c0f00003310d0700100007cc013c000001010010510003000040000000010004000014031000c000000000c3410000000404030000c03300000001003c30030010000100330f000001c100000300000000000cc000004003010c0000010000c0000000cf1010c1300c0300c010000f04103fc100c1000000070c04c0000010010100000400003d001c000005003001010f1d000104000100000044003000000404c00003000330000f0100c30d00313000014300c300030f0010300001000000070000c0000304033000000013000004000000cdc430040000000140000000c0c13000000c000000003100c100400003c0030000c100030030031304300000001003000101000000030000000000000000000000001100000010d104400300c000000000c03f031500000033000000f3000000000000130500000003000003d015000000000c03f0001130000000000000110010030000000400c40303330c04100000000c040100000000103330000003010000000030010c030400000140c300004c0300000c0c000104000c01c0004003003300003001000003333000000411000f0101000000001140d000000000040003000003003cc041000000300010d1311033300101000000000000010043010000c033040000cc0110004100000103030050000100040000000000010331000000004001330000c1000004000f0c030100c0000004000000000400000443140c00c001001400300003000040004100000cc040300000004ff700000103000c0c1000010000100400000000000000c0003000010c04003c01cc0000;
rom_uints[1003] = 8192'hf0340000431c300000440131000c004300100300000f3030030000000c05400000010c00330010030c3501000100301400400104000c03001000050f00000000003140c40c100300000d00c10345c00031c4030fd5173054111000c00000103000710100300034c30d05cc01cc701000415745004c400c04007c1c40c031c000403000c30000007000001000003301400c40000000003c00000005000c3f440000050100303550100003000c03100c300004040000c01c0001030c00f0001013c0040010000750cc040000000003300c304510100400100334100500003030010004000003040000d4f004c00700443c001340d030000004004000000104000c300c0c30000c00010100040010c000c001300500d0040d00c0500c03000c0004030c00004000c00000441001c0001404730010000c4f300001133c00c7c040003300041001d7f0c400000011c010c1000004c0300c0134c4403d35c40c7400010000c005c404041301041010400400300c0400010010c01000000100001000003000000c43037000430033010344030000000010000051030010f3c00c3c004c43073c00103000000000c00000151304041000d0c050014000c41400c1f33000cc1310340000013000000000000c0c000100cc400004c0300300700000400d400303340140400000051001010300000c000500c0c01000103c0000000c000007730137004414000c00140d304d03c03104000000140000f004041705444000000f41000007401c000304300101000030007100040c00400070401410300335d7c4101004441003000010401300000c00c40404000000070400000c0000030dcc0000000040400030000c0011c500140000000c0107c30c0400000001004003000000c007040004c0004c130c0c0cc000c400000010c00c04000d0000000c0014014000100330000300c0010040110c50003703000003000000040f0000000000400000c03004000400000110000004000c00033000c33007003401000740c00040000003c0040f70030004011300005003041c300c0300010400400110000004000003c400000001c0010c000001000c00000000c000c40514044001330010030310000c0000c040000d0300c03700010100c0c400434000c300030014c1000040340140300000000c34004750f03044c404010c34000000001f0000070040f00000040304d00c0104cc10c0100300000010040c0c00000c00400c4c04c0d4074f0f040400000001d000030010003104400c03000040c000100c4c11c043000115d70c000000003000c00100440c15000000f03000074f03000000000001104001100000000c4f03050f3000043104000c0000000001c3400c03c300330004000003c00004040400c100010433077030fc30ccd000040100104000000400000;
rom_uints[1004] = 8192'h4300004004010c00cc0010c141c00c00000100001100c300034fc00041cc0dc0044c0f00dd000704c4cc04010000d70d01c00c0c0430f0d0310c000040000000040004cc0140000500000c05cc00000c00014004cc0c4f00430c0c0104140cc00070c00d040030c0d4c47d000450004cc04040010c31030f004047004c70c10004040004314100440c100000c000040f01c00cc000040f441700000c000004000700474c00c40070001c000043c300cc0c41014c000001c0000100c7430f00001c5c014000c401500300000c3037501400404444c0cc400c300d1100004f000cc04040c000033000000700c3cf44c307fcc000110c4000c040044003000004044fc0c00cc00031400c115700104c03c00044000001300d04410401400704001f040f40000c1c00030000c3000c400c01400300040400cc000000000040040400014f0040000c040c0cc000f1000c0105370c0004404304300c01000c0000010c40001c0301cc4000c33044050000040c004c4d004444050c050400c40104000c5500cc0c0004030c0700c0001500c444100cd501004001014c000c0c000000010ccd0c0cc4ccc004000010c0404ccc000400000c000100cc4000000400c0c710c500530cf40c0004000440071000001c0104fc00400041000c0cf4c0000010000404043f00414c3c00f1400000000000c0ccc501f400041404134000cf004504c30c0c0c00003400f0c44040000004c0c00c041c0c0c430001310dc444c0c1004fc41100140d000c0000004031c40c004c00cd00c40134000011440040000c040040f4010004410cc413004040073300014000007000c00001000004000400c4c03c0c033d1cf4434040000cc37c0c000d003cc01c0040c14f404000f001c00000030404050100300c0c044c0074100c100004030040c10040c0000cc000005004f0000000c30cc00104314f4000000c0430000704c4c0c0cc004404c0c40004045140000000040cc300000100f0004400007c4c0011430003c30c000c074c0000000100d7010f4c00040c3040434c434c0000c000403000d100cc0c003007f0400740c00c300c01d0000110000c044007c0cc43c40104cc00fc000040014c4c04000001df000000004cf000c003000000040d040c044c0dc000cd0c310001010f00010500c4004d0403040343c000c01443004cc044c0f3004c0c0000070700d0c1303040d400c100003100c00043004c0c145c0030110dc0c00000100400013003040c3000f0c050003c0c4c4340c703d0c044c0333003c1000000c0000c0711050c000004cc04030005004101c03c00d00000000004cc0034040004443c00000153430054c00310044000140300000d0c034c00cc0cc3c40c0c00000c00010044010040000433310f0c0dc40000044004400c0000c0c0fd00000500000c03;
rom_uints[1005] = 8192'h10c0000040130004300000300c003030300c400c000410000000000000000400000033300000000010300400dd000100430c00300000300c000000000000104040010004001c00010000004414003000140430104c000100130c030000000000c00c00000f0000300c000000000d3010004100000c0c0000000300000004040034c00000001c000000c000000000010000c0000000000c0000000c00030004300000001000300d1000007011d040007030003000000000043410001c3c00000000014000000000000c30000000000c00003cc014000000003c000c00000000c00000000000f00000000d00c0c00c00c040140010043000300c0000040000000430100040040400c000000c00034030000004f00030300c00d453040d110c041d00000000000411000c00c010400000000300400330000000040010003300000000100000000f00004000003000300000040000000c0000003d0000c50470013c0010c00c0330c137343040010310000d000000c4000040c0300000000c000000dc00000400300000c0000000007c04000c003000000000000304300000040000004d040c30000000000400001040040000f00000040400400c00003400041040041110003434000c00303c000004001c00c401000f010000004140003000400c000000000003400400050000003400000000c0013c04030400c0000c00040c00dc0040000004300300f00c1000000030013700007010c00000404300000c000000010c300070001c0000c0103000c00000301000003000000001300005001c04c00c00043400000c70100c00000000000000000000000004000404000c000c4d110400303100300c0000003c00000033000010000004307004100400004300001003007d00000000000000001c00140c00c040440004100c30003000340400000040000c04000c00300c3007300000340030c30000010c3cc40330c41c3000000c4c004400000000000400300031000440400c00000000f000c000700c010404000000000000000c000c001dc03000c000000c1000400400730000003304000000c000000030000f140030000004300f0000000004003c0000000400000004100000000011000000cc1351000010000000301000400c00103000000003303404000404000c0400000000000000000000000030400100043000000000000c00040040340000700040000c00000000c700000300100000c000000c007011300c00100c30003000430030004c30030003c00c10c30070c030007001100007040000030004033c040001300000034030434c0030000450001000003c0000000001000c00000c44000f000c300c100000000c00000c100c0000300400101000043000000c000030003040041400007d0004000d040400304c01000400f00000000000;
rom_uints[1006] = 8192'h500000003c0000000003c050005000c104000d3040000010c4003030000050040174004000000000100030000001430030003000c40c30000000030010000300040404003000000003c00c0000005ccc1000000033030c300403c03000001003311cc010010000003010000c100000004004d0000c04000030001001c31000c10030003c0004c0003000100000000c303030000c00031c03c30000c00000330014000000104000007400303030041030301000000030c000001313003c0c00000004040c141300031004001c0001c0c0003000040010010c30011303c10010040300d40000100030000cdc003000c000304ccc40300c000030014c000000000000040c05000cc0000000300040004034d400140c000011310004001cc03000000100000040000004f000310004000450041010300030000033300000003c0000700030000000037040000c01350000f000100140000044100f7cc007001010c00000014100330030003004100000000c047000300030000c000000000f340143105100303000001050000000000c01000000000000c05000103000000030000c1c000000001000004400c0c4000c030300000300003404400000103c00070007000400000000040010003110300140400010100400c14000030000000301003c03c000c00035004054cc000c1030c0000c00001550003c3000400100f0031000000001001000000f00100030000000015c040100300130010073100c0f000000c140c004f030300c0cdc11000c00000f30c000011000000031410c3000070000000100700c00000400004400c0000c0010440400013100000100000010c0001100c10431001000c0001001400005c00000000c0000000000c03000c4001010040010003044001000310333100c00000300c40d0d30f014004c104000300004000c000003c00000003010301c4103dc0cc00003300000113400d000010c0003001310040000004c0010000000d000000044000300000c3000003c001400400030000040d4001c00001010043000303000300003041030000c00140000101300301000030110000040000010000003100c300000000c0004044050000403c07310d000000003000000001000000000000010000000003130d41143001c000000c1000c000000c0005c000003010c00003014041000000110c3703004101000c0000005100000015f00100043000000003c310330c000040031000030001030071d0c0000000303c0700403c034714000000c001451100000c00300003100000000143100d0044d30000000f000400c00003300f0000000103010400030000000c0103000c00011000010c0000c000030100000100000000004040300000000003c0000043cc000000000030000011144001000000001403040000c000000303;
rom_uints[1007] = 8192'h10000000131000000000100010000007001c000003000000001030300030040000301c0514000000010000003003000c00001030100015000f00300300000010330000300000d03c00011001004001000304300c0000000000103d0000301074000030000000300000040000000301003030cd00000030001000cc003330000c3010000000300700003104000010000300003100000c00001030000c3c1500100310300000011100040005130c000030001400001c0010103300100030100030000000033000300110100000c000030000311030103307303010301c3000013030000000001000030000100c00003030003000047000003c00001000000030031010001300c000307000000030000300000000000000300300001c0c1001000000010000301000100034000000303000000c0c130000000000f000c70000300000c010040c1030300000100001000003300000301400370010010030003004000400013034003c0000101001000110400000000103100000001c100000340000103030041014003c1000300131301301000c300300003030000030001000301003001000040050003000100011140c1c000000103f00000000300000001000d03d303030300001c0f0010010301300f1170000300000343000101c0010001100001030c030001010300f300000001c040100c00300300030c430000000000c101030000000100003000000000010300c00140000011000f30071000003003040100d30000000300003130000001300000000100f3000300000101100001100000000000000000010001c0000030000003c0000303330103000300000000010100001303c30d33000000010040000cc1010300f303310000000001000010c03100c300330300100033031001030133033300310003000103000000001000c043031000103003330000030000000040c0c1f003010000000100000000000000000000003000000030300001100000000000030000c00303043013d0000c07030000000100000000000100300300c040001003330300c00300c1000000430030031000c10303030300000301000f0303030101013040000000000000000300031300f00001c0010103010000000003000000000013010301000010030000000000010c000f00303001010000031000000300000003000030303410030000030c01010030000300040053010000c00001000301003100c100c103000300c0011301010340000003300303010300004c0303001101f00000000c00010030001001f3c3030000000300700003000003000330000003000000001100000003033000000000000004010300030001000300000000c0000000000070c3000300040300450c000300d3010301000330000300300300000000001014c001010330d003000;
rom_uints[1008] = 8192'h410000000d0030100f0403c00000c010004001004040c000c300003c30004000003301000000c0404034003d0000040100c4000111034c000000040f0000000c000c000003010100001300300000000033400000070030000300030000107c031000040000100000001000000040c000004010404030401050030030c4003c0c00c4003000300f0000000040100000000c0000000000c0310000100cc311040c30c00000030c70030003000040000003034c010000000000000000300000003000030300000300000c00c3030001000000c0033c0100000000330000010000040000010311000000310045c00c0300400000f000010001000000017000000030c00c04c00103040000c00c00c140000000000f003c44000040004c000001410001010000c03041000000000004000000cc007000010300c0400000000d0000000c0000c0050d0000030004000d3c00030050000300440454c00700000c030300000c44c4400000000100011103070400030341000040040f0110000000300003030c10410000000300010030430300000000031000030300100041000c0114003c0c010c0000403000010c40413f010000010300144000000000c000005d0c0430000110030000100310000303007d40040300c0000000010000000001404500c30d030007041411031040000000c000000000101010003c4000004143001c010004d013000100c0010c07035100000000c100110300c00d04d30433010000310c30c0000400000000050143033050c0000701000c0003003001441000301730000404010000003000403130000000300f0c10000000000050343000410300f0070fd0130010330c03310000030050001040100100000c0103100040101000000030000000400100d100070100001000341f0100000300034010004000040000030c0000105001000307000000035000070001000c000710000001400030c001003000000001140003000031140003000001010f30010440304000000000010300000001000010004000003310300103c0004101000000000001100700000000000000c01400040000400d000400000310400003001340c000c3000000003c00100100000401000000010003100000040344000410c001c330150f00000414010100030c000c00000103004004d000030d000000000004000404100003d0003100001100000000070403000300010dc0000030000000004000000300c00f30000143000000000c34100000030300d4004d01040c10130003c40000030401cd03040303c0000000003300300000004d0001c0cc0000110400000000000310003040f1c100010d1d011011010104074000001701007c000300000000001110000000c0030000001400310000d3031100000000c0000330030343013100004100;
rom_uints[1009] = 8192'h303010004001011101000000100003103000007000c05001300000100f00731c440000300010300000031003c3000000040010000100000300000000010700403000700000001c00000c0c404c00000000010000003000c0003000000351001000000000304000000703300000401000004000d0071003470001c00c3000000003300300000000000300000130000000000300300010f0c400100000030000700400001103000040331c00100000103000c03010000003d400000000010000000004330c0000000000001000010100300010000404300100000000034000030004c1000301000310d000100000010c0c70000303000030000000000000d00040040c105100000340c0001000030000350000000c300100c30000005000cf0001c0700000000330000040300000100f011000000001040031000040000010003001131004c00000400300000c113000407040343000c30040000130c0030f1004000000000010000000d0013000100030311f00010d100f0000003000701c00131010001000000000300c0000300400001000c03000400040001000d010403000cf1300003010c310040310103030000c10000301c0d01000030c300300040000300000f40030000c0000004400001300c43cc103000010100040c300000010000000404030000f70c000001300033100c00000003000300050000330500003d40c0003000311300d000040c10041340c40000010000000c030110000130010c30011c040000c00000000000001031001011003000000d000000fc3010014c0301001030000100040000000100030040401000000000000003031f11c1010000000000400c010010343000400400cf0403100000c0000000153cc000040000000f3040030031004001030101400000043033000100010300030300003000c070030100030003000007c004310300100c0100000000000c330041c00300030100000001000100000300000000000030000000000f03013d0000300f030300030101c00301000000054300000003000334000000000cc0030030030001000000001003000300131001003300cf00001033000000000001000000000003c000000001004110043130100000000c0340070000c1030400403003010000c400000c00000010000130c00000000000001100400000004000000000400300000410000003070003030d01c34d004c001000030001033300010300000103000000050100100007c0030000410001f30003040001000500004c10310000330000530301003c003401003100c0031300c40000001c01000005000c04000003010003cc1300000000440003010000030000001440000050000100010000300703c3010100000013003030300000000cc0000003004400000c000031300300000c03;
rom_uints[1010] = 8192'h4103000300000030000000000000010000000f00000c0000030303030340000000010100000000000301000000000001430000000000400000000100000000000000000000000000414c43010c0000010300000003000313300000004300000c000000000001c304000100010000000100000000000000000cc000030001c000000300000000070400000000c00000040100000004c7130000014000000000030001040000000c01000000000003c1000f00c3000030000305000003030000000300030400000330000003000000000003000003000000000f00000003000000000101003001c0000101000000000000000000000100000001000c030000000101000000000000000301000000030000c03f00000100000303000300000000050007010503000404000040030003010000000403005000000c0c41000000000000400301000300c001000300005001005003010cc00101000003010100030100030100001400010400100000000000000100c0c0030003000300030000000003010000000300004041c003000000010000000000000000c000c30000010000000000030040004000c10000000000000103000001030c030000000000000300010000004301400000010000000003030d00000000000000000100013000040400434400c000000000030001310000000000000000003003003100030001004330000000000505030001000300000000c10000030003000000000004000000100300400000030f00000300000001004100030400000100000000500000c000000000000000000000000000000000030000000100000401000100034000030000c0000c000000000000c3000404000004030000000003030000000000030000000104000300110001010103104300000103000300c004030000010003000300000000000f031300030003000000000003010000000000000000000000000000000103000000010400000000000003000000000c4c010000000c00000000003040030003c100000300000000030c400000010300000001030100000103004000000000000000000000c0031000c0000300c001034000400003034300000000000003000300000001000001c1000500000000050400000403000000030004000c000000000001010000000300000001040000100000000001010300000301000300000400000000030000c000040000000f00000100000100030011000000030003034c00040000000000000000000340000000c10440030000010101c000c10000000400000d000000010000c0c001000300000000000505010100000000030000004000000300010000000004000000000300000034013c0c000300030300000301c0010300010301000100000c0300000000010000000000030;
rom_uints[1011] = 8192'h400000000c01044370000000101010430100f0c0c0c000000450c00401404000c003000070c000c00370001000004033300c040000c00000c34000c0004000070c00001301c000c0000040003001c0034100d3c000003041003100000003c05000745030c0000000c40c03c1c03003c03143007c0003004300000300c001504f7000000101f000c04010000c10c0510040d00000000c40c0c744014003407003cc0400000040410050c05400c0400440430000c0004c030000c00c00c0c010030110001000035003c74c0001400303440001c00330441000cc00010043c040004000004300c5700003400740000031040001d4c0c0000000c0000001034040070170c0400010404040c0000404030000300000d000c0104cc4000157403004300c100000410104000000c4c00000010003000300c100c0000401cf0001011c01c04d70300700c00000400140034000037000c00000000c0c414070c003434000c300400100000010310140001001031103c0ccc03130f40303f000000f471f00d330003100c0c0d7404300c4403fc0000000000000000040c0400030000000000c003000004010d00040c0003000c0400000001371000030500c000000000d404003f0000000010300c00000000000405070400001010ff00043700000400010c170370000000300c0d04000007003401000001003700000ccc0010300c00fc1000001030040c00003400104000c0153404000074400c100d0301300d000001000005400c0400100010003000100104001c170c0d01000000000004300017130130000c30000404003000040001300000001100310c0c00103c00410010cc0404141000300300001c0001040403000400000c0111000d01000000040700300c044430300000000037cc1c10000c3300c01c30000c0c030000100304c101143134030050103cd004003f013c0c0c44000c00330003010004d1040c3c001530000331000000000c30000c0000300400100004000030010001f04010043400100154000000710c00c0000340030c01000000000cc30100000c0400f000100c03040000000400040000c0003034040c0c010000d50301c0040004070004140c100c0101000004c000040007070c000f01000000000100003000370000000000050000100410000000000004003400003000000c00303403003433300d000c0c00000001030300c10010000000000400004c0500c0c000330c0400c30070000400103400c30001000030d01004f004000004010cc300040010001010c30c000c0030013c0401010000000400000403000033047100004300cc00000000000f0c030000010c0f00c004340c0004000c0c000004000000041300000001000c3030004000030c000c040c00030303d0000000130d0c00100404c033040f000c00034000;
rom_uints[1012] = 8192'h4000000044c0000c00cc0c0401030300c300000c0c000000000f4f00c4c3c00300000000040c0100000c04000d000100c00c001c000010d0c00c00c000401000c0c0c0000c00000c00000c0000000c0040c0c004c00003000000003000000c3000c4300100000000040cf1000c00cd050400000100000000000100cc0c030000c000004c43000003400001000000c0c4400c040c0000c3c001000c000000400c00c40440440001000405030c4303000000430500003000074c0000140f400000c00000c0c00000100c00000000000c000000c0000003c4000c3f00000010000000000000007000000ccd00040004000c00000000000000000c000000000000000044000000010000000500c0c0000000401700c03c0cc00040400004000004000000c000000000000003000000000404004000c00c00c0000000004c3c0c00000c03040000c000000044000ccc0c00010300000100040c4304004000000004c0000000000000410000c100000004c0f1040d0000c00303000c003044c00000000c0c000c03000000c0c000000000000c00000c00040040000000000000000c00040000040010040000010004c404040000004c0300000400000004000c404400400104430040000500c130000400000001000c130004c01c0000000001010400c0014441040004730c000fc1010000c70000040000000000300000000c00040003300070cc00000000c1004000000000c04340000d00000c000000c0030007c00007c405003d0400000300000000000004055700000000c404c0040c00000c0300030014000000000000000000040040000000c000400000000300004000c00c00000040c003c00000400d000c0400c100000c00000303004000400040c100030030300cc0000100000000c4044040000000c000000c54cc0000cc0c1400100004050001000000000000000300c0c00c00340c00000000000000005000000c000400c400c000000c000000c0c0000000000c01400c000c000001400400040300cc000d0044004c40030000010c03000cc000c000c0000040000000000c0001004c0404004c004c00050000c3000001000001000003000000000000000500400c044000000300000000000c7400000000000000000100000cc100000c0401004004000c0000000000000140044c0400000400000034000000040c0000004303000000400300000004000100000f000030400c00000000cc440c0000000000000c0443000cc00001000c0003043000c00003000000010303000000170047000003000c400c4000034000c0000101000001000507000c000d000000000004c0004000cc030d0c30c0cc0000000400000000004c030000030c00000c004c444000c0400004000c0000c00004000400000c00cc03030c00000004001400cc00000000;
rom_uints[1013] = 8192'h400007c000000c400c0000000000c0400000404d3000000000c0c10dfd400003000007c300000c004000c300004101001135000c40000000c0c003700000000107540003c00040000007000003c00001f0cc00c0c330000100103000000000000100c54100030300000000cc174c00000300030d000000000000000041000f7440300330d00300000004c000030141000000000000000000400041034f000000070000000300030000000100000040c044c0000003c0404000000100010cc400c00000000000000c00000cc0c0001000070041000030000100454340000000300000000000c000000004500c0c004010ccc000000000000400000cc0000000004c30f0704004444d0000000000000c00010c0c0dc7010303c1030041030f0000000000c00000000303000130330000000000410001000000300100000000c4000000000047000001c0001440000300030000400304000c000140400300000001c00001d00000c00043000000040040c0000100c00000000c00700c00c0c1014040c005000001004100000400c0c000000100000000c003c00000000000000000c0034400c407d000000300040100000003010300010040c0030000040c0003001001400c00c11040704000c0000140c1040044000440c00000000000000000c000c0000003c10001430104004000014c00c4004000000030000303000000440000030000000000040040041000000001c0c000000c44010000c040000040c300c440000f030300000040004030000140f00000000c1001011000404000000c0031c04003c00001c0000000c0040000010400400c0000400100000300000c0000c0030d43004c000030000000000c0c00001000400000000040000143f0000000014007000c0040d00400000000c0c00003430105000c4004004000c0010001030300000c0001000c0000c100010000003413000003001040c03000000000c01001c000000000c0c100c0c3030000c0004c0000000000000000014000000007d00c00000400000000000000000003030000c4c00000c0010000c030c00000040040300700001001010c000000010001c4010000c00c010000014000000000c000400000030c00030c4100c000400000c10030000400000001c000c000010000000304d00000300100000000000c000003c00041000000403d03c000c00c040c0000000000c001010040000110000c03c30140000301000000c00300400c00c01404c300000cf001d0c00c00c30004010130cc0000400000c003000000404043d04000c300040003004000c0c00000000700400c00000000000000000300c0000140700000cc04030c00000340000000000000400d00034000c040000000000c03000000400c00010000004011004010400000c3c0c0000000000041000050c;
rom_uints[1014] = 8192'hc0001000c370c003000300003000fcc0703000003000c0000000000030404100003000c131c000000030000000007cc4400110c0001004300000f00001030004040c0001000000000000c00c400044c00300c0011310ccc0133001040000c10000c000100000000400001c000300503000d01c100dc1001000111300100100001070040330000000003000c0cc013004c3000000000070000030f30040013c0003713000c0304030c0f030304c0100c01000300000010001c00000001050001000d0d0330000c350f0c3c000000043007000004040c030d0001c00c0dc700000d00001307400c000000000403d0000000001000400000000004010000300000000000700100000003140c001040000000000003000433000103c1010541cc1c010003c0010431004001c3400000050c01040000000300040000440f3501c000100000110c00010c04000000400d04004003301003040c03001d0cc1c000010c4100000300001c0000100105030400000000400100050c330c0144cdc1000000030300001004001000700000004301003040004f0c000dd43500040504000300011f00000310000000050000000c010010301c0001c1c000100444000004000140c01000000d030c0000033000c000004000300050000f000c00000101cc40d00d0170003c00000c000000107100c01d00c307444cc00005040703000c0000010cc4000104000d0c03034c000f4017c3033040000f00003404700100cc1000000040d040000c00c30001c1003031000000000010014700340c00040000300c01c40000000000000c0c000000000f030001000013000000000040001300d0000f0c0c04030114000004010303073004040000000007030c04010400100c00000100304000000100000000100c0c0c07000001033000000001c0000f4001c5000c474353000104c3030c0003040300000f003000300007000c401001003340000403130000400001010130c000003fd001400307000c3001040d000003500707000c4000000403011d0003030130c0000c000d0013700000c00040000000000300000000000c000c0c040c00131040000070400030000000000404c100300001000704000c0000003034000cc033000f1000100c00040c00003f00000cc00400010000000007040000000cc00f0c001000c40400004011000011070c0004000c0304400000c0d0c0030f00000c000000000033733d01300300040c1000034d010c0c000300000001c00c010c000414000f00c00010000fc10004010c1001030000c1040000000003c4000000040c000d1c00035044010000030f0f0c00030300c70403004104010007030000000400000100300040030c000c04c1040c0c1cc103000f0000400100100c00004001000c13030710000c0f03030c1010040c0004030;
rom_uints[1015] = 8192'h30000000043c00340000000c40000c003c3c0000010400340000000000500c00000000d4300d040400400000000004c0000c0000000000013000000030000000000c0000000c000c0c000c040c0c10040000300013cc000000000f0000170c0400cc50000400340000000c041c30000000c0001004000010000400340c000000030440000c0c10000000000004000001300000000004cc00040c300000c03410c04130040030100000004400000400400c040c000000000044040000001300000000000c0000004c14300000000000040400000044040c00003004040400040000000000400000000030000c0400d00c005c10000400000400040004000300003c4c0000404000303c00000000000000000c000c00040c000cc3003004300004001000000010000430f44c14000000000c04000004040000001c100004040000000004344014000c304000100c0000c4c0000404001004000c0c044000000c0c004410004c143c00c0000004000cf00000000c3cccc4000000f00004000c0c0044340c00110400170004000000000004100044300000000400000010040c0c00303c0c00370c0000000000140c00500000c0004000004c000000cc0c00400400c4000000c00c001000c00000300000044000401c0004000c00041004000000000030000000030c0c0c000c000030000c001c0c4c0000000400040000400000100cc0140c001c000430000c00000000c00040340007100010130c100000040000000c0c000030003c00100000300400100400300c001000000004300000000c000004000c000000000004c00000403000003000040000143000001004000000040c1000040c0030300000000010040c00040c10d0004c00000000000404c303c0000010000000040430c000d0000000100000350014040c30000003041010004c000c04c400333c4000140c0c001400100000000414011440000040311440000004003c00000004100000000004300c000440c0000c0400000000000000004000000003000000100000040034040000000000c0110c3c000cc70c000c00300400000000043c000c004c000000000f040c00000c04100000000000000000000c100c040000440c000c0c000404000c0c0000003c00100000040000003c1000000c0030000000400000000400000c30040000c004300c04000000000004000c0c0c40300400c00000044400003010000c04003c4c00000c0000100c00141400000c00040d000c00c00c0d00000000000410000400000430c10000140000040000c00004100400000000001010000000000000103000000010000004000000000030000440100030003000043400003400340004000000000000001000043000cc0c040000c0043000100030000c0000330000000000f0000c100c00000034000000;
rom_uints[1016] = 8192'hc30000000c040c134c0040c0003d30c0000cc000000000c1500000000010000040044100000000001c30000000cc510000c03d00c10c01000c00300040000c00000fc000003000034040404000004c00d400c1043440c4d10cc0040500340040010040c000c400c0c000c070cc000044cc0000c04c4000700010d0030003000000334030000000c000404000043440000000030c0001cc40c00ccc7014c0c000c0000f0400000400000000700000000010400c04047c00400440f000c00101c000c000070040100000c000cccc010000c0001c144010c00700c034700c4c0c00000f0104000000c0003003003000714110c040100030000cc00040000000004c0f034f030000700005c3000300100031cfdcc015000000700300c0103400000c0000000400c04301c00cc001030001000c00c00000000400410cc0c00000104040c0040cc001d00011c0c0c00404cc00c0010507c100000410c1000003000010050040400000c044f04013400c40004100000044040007cc000000000000c0cc010547000100c000430000c00004000000c0000440000cdcc1c00040c04441003040011000c0000105034000440300cf05c03431457f001400000000004004000c000000000000c01000400003013f100543000001dc00040000d00700040c050003044c01c10000f0003000000000000010000040c0c1d000014003450411c0cc0cc0c3100003430d000731cc03310001000000f01000c10044d1300000c5000000030440400007c000001000c04f04400300004044304c0310400c040c000000100000c00003000400304c00000101700001c0c10000000007003c00c1014000050130044c00000c4100000040c0c0104c0c0c00c0cc03000c000003c040c300c40404c0004100040741f041000010400010c34000040300c4c0c034f0444004c00040f0000110c0010101040c100104c001cc03000003f1f040000003005000cc00000140c00003c000ccf00001400301030000c5c001034000000004000000c501c00c500400040000c00000040401000000c1000000c00c00034001c3103c0f000003000000003c0c000fd100c00001c1cfc04001c0010f00c0050107000043c00c40ccc0334c0cc1400000030043104c0000000cd001c000ccfc00403300c11f0c00003300030cc105400000c00730c40503c50115c00000c00040000c010004c004cc00400000000003c0c30cc040cc00d04c1433001403c0001300410c3000004c05c00000000000100405001400000cc00c0c4740000100044040d01000040100f001d0004700000000070f00f530000000030400030001c00000c3501cc40001000000c0000400143c040c04400dc00000c1cc00000000c0000430400000000400c47c4c00000300c00000000f0cc00d0c004001000400030;
rom_uints[1017] = 8192'hc00c1000001004000500001c000030300d0400c13010c0030000000030c010044004000134340000000000010000c05cf1500000000000304400000c000000c0040004000003000f00000c1c04003000000010054410301000504c0c001103f400000500004000000410010000c701300000000104404041c301c000440c30c0033cfc04041000040000400034013440100c0001000c0040c000c00000f0000cc0007400300040103000300001c1003040000400000040c500d40004c100000000cf304000000401000000000000f0000000400fc0c000000f333041f0ccc001010d000001cc0000000100c1303400cc00d00300330000000000000340003000c0d0c0013110471c04300c004000000000170c100c001410c0441000c00030d7300100000000d000040000cc3000030000c004000000c0000044f5310f30444000003010300001004040004c44004000000001004000000c0030011000c00030001001001c3030040033030000004fc10004500040101300c0d40100010c030104101400ccc000000cd100007c0c030044004c4000000000000c300cd000100cc10300c00040000000000000c0401400c30000141f43007000010000c00503000054040000007000000031003100010003c00001000100000c00c000000004004000c7103000431d04401c000000000305000004000c04034ccc4000030030d1d4003c0100400000301000100034043dcf00040031d404c00010400040c00004003007000050000400341cc440100c00cfcc0040c00f043004003010c0000040f0004013000c0000c0c10010000400300040f00100000403000c10003000c04410010c00013c103030040000100040700400001000400040000c4000300000001030000c40433050000c444c3410c10000403c00100fc00400040c00400000340044014704315000c30f4c100030104000f0c00c00040000040000d00000c010001044003000c000000400403000dc0300c000301103c01cc004c0744c30047000000310c0000000010014144010003000c00c100040030c000000017c300c00030100c00040105001000104000000c01c30000000000c0c004010030030004440d00040c00400070001103000c103304031040000000000000001033000000004f000000000000000000030c000034000000c3c000001000010c00103000c100034cc053040005530410c000000cc00700c0000000c040100400000000000000000000c00000000003301c13300400140c000000000f00030100400000000004c00000c00043000000000030010400c0047000c0004040000400400cc001c010050cc470000c071c00130040000100030010004010040300000c00000000000000004000003030000100c41c0000140000000000000703c7000041300400004;
rom_uints[1018] = 8192'hd0001000000010000110303000103400300c003c3000f0c000000030c00c30030000031000000000003300c00010100000003c00003000000030100013000001000000000000c30030d0000030011c0000c0f00000000070f4300410001000010c1004013010040031041014005000100000000f3000300c0c00370000400430000000300001c070000c00000030000000040000000000cc0010000400300000000c003430000c40000c0034303000000410000000c333300000041030300010004000100001000c000000c0343000000005c00400144000104040300040300000000000101c3c04cc30c000c0c0000400000000000c000000500c50c40010405c10c000004130000000331300300400011070331000030000100000000000043000003c000030f40100c00000300c0c0c00000000000000001030c0007000000030300034103c3000000f043c0030701c001010c1010000100330303001550000300c0000003010043000333400300f34000000314010043400f0100500000040000010000030040030000000f000001000000004000010000010c100300c0000000000001030000310000000041000c0300010005000100000003010300000000000304c300000000000040030103030000040104050030110001010503004c030000030040000004000c000004044000001000000300404000d0c30400040400000013000013c40c0c04000f03030300000000f00f100c1000c010040340140f000005010000001000c0010c00004000000c100701400004004000000103000000000c0000c000000000000400000001000d7003000003010010000400c000030300000000000004000000300c00c0010000400300000104014001000301004000030040000110000400000fc003000000000fd00700011304030303040013c00300004f000f00433003000000000003000000040c00030000000001000000c00001c0000000c1004300c3000300033040000000c003400003400000c500000000000501c30c004333000300000000000001010401030000034000430000000c11000000000400000c000d000100000301000100000504000501000000f340000000c1c000400000000033100300c0000040000000c30f00010341000000030000000000000101000003c10001130401cd00001401c0030000000005c3000000000003000000000003c300030503300030c1000c00000000010c4103c00000030f4300c000000304000143000000c10000c0010300000000c05340400000000050c30000000040000000003045000001000000000303c000000c0000c00f000000470100000000040000000000000000c0c00300c00000030000000003000000040303c0000000000000000100001c0f01000000100300030;
rom_uints[1019] = 8192'h30110000c000c31000000f00000003340300000001c003007330000000350033404f4c00c3c000000000000000f1000504000110030000c30000400f000000c000054010000000100000400400000100400003104000f0c0004000000700050001400740010000c044400000010513c1d0c0004c100070000003d40000000001034000400c00000000004044c0100003c0000000001030c00400044000400000c000000303030010004000104000070303500000000010030d0000c00103000300030000000004c01700040000300000c034c001010073cf03cc4001c50000030000101d100003000400040cc034414100cccccc000000330000c0000400030040000f0000cc01000413000400000100c3031000c301004fc4000cc40000c4004130004c3101000110300130c0404cc0c00003000001000300000300000010700c00050131000013330000340003000003001000001404c1400711000003000000740030000000007000010000074100c0000000030000c0010c000000030133c04000001000003004000003c0c0030000004110004033000000000003010174430045c3030003300c031000000403040000401341400400004c00500303000c00000004030037d0030000c00000c00303000001704400000400011430000003c00003000400004001000040000013010030400cc3303003000011300400000100000000030000c04000030411010001400003000000013000410003004340000f0700000400400000100043030000004103000000004010010003000000033004030c0000f0000001000000000040c00300100003300c0010000010304044000c300013000103c000300003000000003030000000c34f00f30000451cc14c0c040300030000d03004cc00005033004140c00c3000000040004400730c00003300000000100d0000c053403340cc4000000000000001770c0333c00003300cc500000000000101031400000041000c0000030004003000c4003007c0c04c000d000000c000003110d0000003c000000010353500000c000300100040004000f34314034340004f040010000000043103004003030000040000000443000c0043100000000001010000010f000400030000300401010030000000100c0303001c030c0c0001000300010000330310110000000000c0000401c3030000000040c100001000c3004007040043400000100101000110c0411d000003c000034040400401004000000033000014c000301003004000300140003c00c0c31300c030730430000300100c000300030000030000001040300000000300000040000d00000100010040c0c40014000c003300040033000000c0031010040031cc01400300000000000000000304304300000c0041004f101000c0030000000000000000;
rom_uints[1020] = 8192'h4000000000010c010000004301000030100440c003d01001000110300030010404034071d0001000f00f50050033100103333000100c501010c01c3040000000c07700d10440100003000001001341100013c401c0300000130f00c3c000400043300030101c300041000000c004d03030fc033001c03001c1031001d0700100101030f000014000d000430000c0000300000000000003c00000070131030110314100400001d00003710003001300c500100000000ff3d3400000c00003330c00151000001c0c4010011003010170c00141c00441000013c30000034030000050000011f0310000d00300300001c030c033057c000030c03000000000013403c00013300100000343c310014330500c000000030430001000c1f03003705033110001317000000010d0304040c43101000000010000003000f0400000400d0140005350030001c00000100004c0300400004111c00010000000001000000100000041c7344c313110007500c300d04000000c103000000340f3407000004110301030300000000000000000000030100310300000c100c01000000100c0030010004f54103000003c0300001000f0c00003003040000000c003000330303304f3010001330300d100500003000013c000c000040000100000703f134c00c0000000030013010003ccc00030c001c03000101000100030001000010cc00000000000f00010104c400110000300000310100105000f10474000000c13000051130003c00413c03000045030100000000c00c000003030c1300043d00001c00000001010000000004331004001f100c00003f010010300c03cc014300000d3001500000c300000c00c040004c0101010001400400101040001000040433040c0400000f100c0005100033303430010303431f41000000c0100001003c0001400000040010003330010f0c1314c0140f100001000000030d3f00430d003010304001740000000003300c00410000000c00140000010513000c000c3400000f000000400003030003300010041c030c030000013400010100300000000010070001000000d05003013100000c0111000000003000030400700100011103000cc0103c00c00c00c304100004010c0000003030043403041c00330130001030034000300c370c300c0c033000000f00d03c00000010cc41000000010000041000c000c010040c00013c003001050001003115000100000431000000100003c0000105350300000000000003030013101c1050040030070030003000300003010010000d1010001f433c000c0004003000010040011c050000303030040001003010010040d000f00001003d300000410cc04105100000300000f00c3cc00001000c140017000c330000010000300100000104000f10030010013300070c00000000;
rom_uints[1021] = 8192'h33000000040c000000000000000003100c0000000340000005001000000443000000010cc1c00000000000000030cc003000000000c0300c141000000000000000c400300010100000000c04400000001c3000030000010c3f0010000c30043c301401003000001cc30400000030003000010000300005000000000000030004700710040c0000010030000000000c40003c000000003010004030040000001c03004000000000001000000c00400100010001000c00004000000c40000030000000000000030c0dd3000110000000000c704030040001010000000c310000010000000004104000071003400410c03031000c40045003003000000004000000004000010030000000000000700000c0000c0f0400000000c0440f374fc0c0400010100000300301003004040000031001000300040300000004000000000400000f00440003c00cc00c3c0f00c0030700107000050404d0c30c010434000003030000000100c030331000000c0314400005010000000004043100c00000030c330c3100d10000001c30030d300000050000030000040c01c00cc000311000003010140f100c0000000001003c0040000000044d141000040070000000300c0cf131010000000f0f0000c000c300300000000000334c0c0100000000000000c0000011000400c100d00c000100cc0000000000000cc0400cc000400100000000000000cc00100c30000301000110400400300000c000100300010c1c30000c01400c074034000440000010003070400007c01003000040c0000c00003000400001000c00100000003000000000005100430000000c30000c000c004013040400010030030003c00000300400300d0000000000f40000c0000c3c00100c000001004c030000000010001000000010c0c30010010c330000003c0000030000001001430c000003c004000c000c0030013010c000000c0000003c00003043000000014040000000010030000000040000000400c0000000000000000000000c031410000000500000000000004d00300000100400fc0c10010000030004000000010004500001300400000003c001c0000000000c000cc004400100001000000400000000033405c00000300003c4400000040000400c0000035000100003000000000300d00000000004000000100004000c00004300000004000d000000003f04000000d0000000003c01c0003000040404d0c501040131c004000100300130000054fc000000000f0000000000003000000010000c00c0003000100c000000450031c0300000000001310c001c00000003300330000101c0100000000000cc0c00340100000000000000d00c0001000000040000040004000100340d140000040000000000000040004140000034cc0c0000300010000000003000130000000;
rom_uints[1022] = 8192'h400000410d00c0000003000003010430000040c00001000003c0c000c00d000000000001010000001400f1000001c0000000000000c000400341000000000040001100030000000000c0030001c03000f0450040c00130000003c04017004140ccc30001c000334100000033000000010040d1010d000000c03000c30100000d00d0000131004100000045c00030300105000000000000040000000330400040c00000001000000000d0c0400000c340037000000000c01001000100c0c00003c300400000100040440003330000000010034101010144c30030000c400000c0000040050040000013030100c10003c1c041c304400000c3014000030000c003c04d00c00001c300000000033300704030c3440004010400310340004001000000000000000100004540cdc001404140030c01400100c03000000010004100041cc010c0100000000000d30000c30c0c0f3051400000000103c30100010f0700c3cf50c000030c000330010001000301c00001c01c0103007d00c1100000c0043040133101040030030000000000000000030001004100000303dfc044301000450000400000010000030140100140000000100001000000c030130000c000c30c00c30c0030c3000040000000001100c0030003004010010001000031710401400100410000c30034130000030c7cc10000c04000000040040300c10000c00004c00c00000011030440c35c3130c3c0d30000010040c300000340414c3144007100034c000100000040000000d000000d0100000000cd010100100001030300010400400f400001c1004c004003001040000003000000001300030100030304f4c30003c30100000000c11303000000000001c0030340c0410000110100000010004343030040301c00c0005301c1000003000003c04003000000c00c0300034100c0c004c40c100000431010000100d003000040c307000040400003000c010340000d000101f000000000c00000003000041033c0c3010400c01000004001000003030003410000010040430000030001dc40013000c04101d0c0300c000300400003000041d000150000f030033400c301400000110003030000c000c040000001c03000010300c000c0003000c0c1c00000c100c003c00400000000c0513000010340c0000300010000001001f000001341300041010110000000c35000304040c0400004c3030404c00043300100004000103700000c400031c3000071100303c3000010c0000010c04f100070410003c041c000f0000100c0000000c030ccc040001c010f000300c0000101000043304000004003004000f30001000100c000000001000004007d40040401030400c410000341c0f3c0c30000014c01000000030300c00cc1c000100000000300030003000000c3c1014000400000;
rom_uints[1023] = 8192'hf000030000c400030c00c001040003c0010004c40000000c0d000100040000004000d00d0004000cc10001c344300000030ccf00000500000003001000010007010000003003000001010c0000010c0400c43ccd0c000c00000000010c11040c1d0001c0411000000140000001030404300010000000130c030400000300014704100cc400004113c0000c040700001400c0c00000400131000000030404040500400000004040000000030c0000cf000000000c10010001c00000000003c00cc00000000100000f000c00050044000c4d07000c0000030300410c030c00001010cf00030103000400013031000c0103110031010004000400403001000d0c7300c0300000400d00c3010d0100003004400500040d000000430d010100410c0003000f0101003000c1010001001003104d000000030000003000010d0003000303c003cd0d0c030f000c010ccc0100000c000c01003017403301100003030c4101000401c00c0c110c000013300500003000000c400c0001f010101c030004000000000100000404000000030d3c01c00000030000100000030c0c0000000000f30d00034000000c0000000cfc000400000000000000c00003300004cc10040000034000100000000000070000d100d340c0000001040000003001000000303331000000000c1004cc4d0dc300030100040c00000000c40430000c00404d0dc000c3d0400d010000c0040001c00c403000100000000001000c53000101010004c10c00010000000300040300030000340330000104100004004003000c0003110000000c00000500000d000003400dc40c0000000030000f00000c00074c000c53000c03040000000c0d0000000c003040010103000000474010001041030001400100400c01c0011003cd000714010c000f040300c0000d000000000000074100c00040c00100044300410d00400c030d01c1040c0100300c401100c03001000000000001014c04000000000000400c0c500d000f04c1000c0000000000cc00000401401f00030030010040000000000105c301c3000004c30313040300004030000c03000000000110000041040100100400000410004c04000f400c0017d000000030400000430000040000030001100100130040010c0000c00100c30400c303000704734005c000010000000300000044c00000c31c0c000007400000000403c30c000004010010000000110340070cc00c10301000000044000c03030d070f43000000000000000f0c00400c0000000100070003000c03404040000c1103704d000c07100000000000010110010000000000000001010000450401000533c04004000030c00c0300000001000100103004c00503c11004040100040000c0000100300c000100000007074001000300030000001f00014300000d034;
end

reg [8191:0] outputReg;
assign out = outputReg;
always @(posedge clock)
begin
  outputReg <= rom_uints[readAddr];
end
endmodule
