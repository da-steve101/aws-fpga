
module DenseBlackBox3f4b5cb0a2(
  input clock,
  input [9:0] readAddr,
  output [1023:0] out
);

reg [1023:0] rom_uints [1023:0];
initial
begin
rom_uints[0] = 1024'h400000000000000000000000c00000000000000000004000000000003010000000010000000000000000400000c000c0003000400000000000400001c00000000000000000c0000030000000f00000000040000000000000000000000000000001c00000000000c00000000000000000000c00c0400000000000000000000000;
rom_uints[1] = 1024'h30004000000040000017c0100100000001000400000000130040c0c000000300400000003003000000000040003100000003000330301000000340003000000000300000c0010100c00000c00100400100c000000000000000c0400000000000000001000300000070000000000000000003000c00c04000000c0000c1400;
rom_uints[2] = 1024'h3300010000010000000000000010010c4c00000000000000003003000000000003c0004000310030c000c0010400003007000070004003c0000100c000c010000000cc70030000c00000000100c00000000000d040000000c0c00400040c00300033000c03000004004000c00000030000303000300040c00740000000010c0;
rom_uints[3] = 1024'hf000000000000300070004100d00014000004030000013c0c3400103000000400dc000000040434c040000c00000c04000000000000040c000130040000040400040c0000000c0010f00c00000c00340c00003400000030300c3004045000000000000000003c0010300000000000100000300000003c00101034cd3c100;
rom_uints[4] = 1024'h4f01000104101cc000000000c44c000000010410fccd0000c000c0c040401000040c00100000000c4000000000000004040000000000034c0000000043000c00000000000000000c0c10c0c003001000000040040000000000001000000c30000010003c0000c4000c00000000c0000000000311c004000c00000040000004;
rom_uints[5] = 1024'h30000000100100000000000010c001000040000000004000d004000001c300c3000100400010000000000000000c0001040000004000000000c000000000000040000000104c40c000000000000000c0030010000100f1000300000400000000000340000001000003000040c0c040c0c3000040000;
rom_uints[6] = 1024'hc1000000000043003001c0c4c003100000004000403000400000004000f040c000007000100030000041000041004000000400fc004330c0033050c3000c00000000c0303c00c0031000000070003010003030300030000040004040100040000001c0c0010010000050400400c0c00000f00070004000c030310000c1004000;
rom_uints[7] = 1024'hcf00010000000010000000000000000000000000000110000c40000000000000030410300000000000000000004001c00400000000000010001c0040001000000000000100000000000010000000000330000400100000300400000000100000000000000000000010400000000000000000100300001000000040003000000;
rom_uints[8] = 1024'h1300000000010000000000034000c000430003004c41000000000000000000c000c3000400c00000c341000000000000003000000300000300001100400000c0c000000000000c00000040100003000000000040c00000004000000000400010000000000c01000000000000000000000c00d000c04003000000d000000400;
rom_uints[9] = 1024'h400401c04003cc04cc000000004003400010cf3c00040c000c0000000000000c030000040000100c0004000000400400000031c0030000040007000000041000035300040701000400000700410c0400044003000404040000004000000400000003000100000d03040000c000000000000000c0004c0000004c0010001;
rom_uints[10] = 1024'hc00001010310c10000000300400401400030000301000c0000010003000000001000101401034000c00001010100000010000103030000300001000100000001010004c001000000010101000c00001300000000004000000040000010000010c10301010f000043130000000303030000000030004030000040d000000000;
rom_uints[11] = 1024'h3030300014000100011000400001000000000100000100000001010000000003003c4000010000000c3000034000000000004003003001000001003040000000003030c0000c0000001000400303003010030000000000010010130133c010000100000000000000000000010000000400103004000000c01000000000000;
rom_uints[12] = 1024'h4010030040000000000f0c00000040c400040c000000470003f00c00000000000c01c3030004400c00000050000000300004000007010c000044130001100d040000300300001400000300130001300000000d00300004040c4000dc0c040003c0001c044c3030000040000000dc0c00000000c00300f4100100000c0330003;
rom_uints[13] = 1024'h400000307000000001010000000400000f10000440c000000070000000cd000c0cc0000000000c0001000000000000030000000000c000000000004c0040000000010000c100c00001000000c00100040040000000c000000404000000c03040000c440010c0c0c0000000c0c0400004000c00c00000000c004300c001400000;
rom_uints[14] = 1024'h4f010c0030400701040044000c00cc0000303000000030000001040000450033c0000000c000c0c0ccdc0000100004000000300c000000003000000570700010000003000c003000700d000004000000000300000003000000043000cc010000c0c00330000c00c003000000c00010000000003000c400000f00000010341c00;
rom_uints[15] = 1024'h101030000004c10010c0000c0000d0100010c00000000000000000000110303000003000010000130000000331000000100000000030004000011000000000000000100000000050c0030030031000305000000050100040000000c5000000000000000000300c00000300300000000000000030003000300000000000400;
rom_uints[16] = 1024'h3000000c03000001000014004000000040000010005000001000003004000000000040100004031000004000c00000000000c000f00000400c00003040000004c000c0040004400000c000f030000000000c0000000001c001c03c400300004c000000000000040c100000000c300000c4100010001000300000000c04c1c0;
rom_uints[17] = 1024'hc0100004003000000000f000040000300000000403000310000003103000000040000000000001101000c00001d000000050000000c00010000001004000000000c0300000000000300000100000000000030000c000c30c0004001000510003000003c000050000000c00003000030000000000004000c0004000000010000;
rom_uints[18] = 1024'h130430000300000400003000000000000030001000000040100000030310c010003000000000c0000100004000003000000000000040000000c0000010000000000310000000004000100000030000000003000000000000000000c000001000001000000000010000000000000400000000400010010000101001040;
rom_uints[19] = 1024'h100100c003c0004041003c3000341040000000000ccc0470c04000000400000070000000000040c000c00400000040400c0400c000c050004004c0000cc0000000c40004000004c0c0000c010000100004000000000000000400000c003400000000000104000003000c00000000000c0300c0004040000400000040f0000d4;
rom_uints[20] = 1024'h1030000001000c0004000c00001000300004000400000000003000000000000001001030000000000000c0000000c0000000000c40000000001000000000000c000000000000000000000000010000000000300000000004000000003000000000000000000000000000000000000030000c000c000c3000000000000100;
rom_uints[21] = 1024'h3c01030d3c41000300004000000d03000103c13044c003110d00000700310003000c00100300c000300c30030d1074c1c0000040031110c330000c530010030003010f013004c1101f031000110004000301040331c00100003001001f0000000403000c0003030d00000033000003000001003007047d000035403000010101;
rom_uints[22] = 1024'h130040000d00000040d010001100000000000000c300000cc000003003004000c0040041004000030000000004300040004c0003000c00c30000100000000003000300400300530000000040c303c0000000000000000040000c00c10000c10000f100001001010001000100000300010000030044000000c0c10300c000014;
rom_uints[23] = 1024'hc0400000c00cc00003000400000000000000003003000000000000000000000000400000000030003000304000001000000000000000c01000000000000000040001c000cc000000c0400000000000000000000000000000010000c0000000004000000004000140101f0000000000000c000000000003001000000000000000;
rom_uints[24] = 1024'h30c000c04cc000cc440c00040004000c0000000000c000000100c0c0000d0003000000000c00cf000000400000dcc030000400000100c0000f3000404c0000000000000000c000000cc00c0410000000c000000000000040000500000c00040004c300000f00000000000004004000c4000000cc000004000000000c05000004;
rom_uints[25] = 1024'h3004030c00003c0c001c0400043c1c00003000004c00040031040404001c10000c0c00cf10100c0300100c003030000000040000f40003030000000000000000000000140000000c3c003004000c04011000033000001000000000300d00000d3300000c000003000300000c0103003000030c0c000f0c0000000100010c10;
rom_uints[26] = 1024'h400c140300f0040414100034c00000003000000000004000000300000000304c0c000000000000001000001000000000003000c00c0000010000c00030000000000000004070043000000cc000030004000c0000000010000000010c00000c004400c05030c0000000100004c000000000003000100000001000000400100;
rom_uints[27] = 1024'h4c000001410300000101340c000300000004c00001050000004c0000000000000000004400000d00030000400000000000000100000100000001000d0d000c10000c00c00c0000000c41c300000c0400410000010000004000000004000001000000010c000400c0404c00c00c000004010103040c000004010100000100c0;
rom_uints[28] = 1024'h40f00000004400c01051040000400000330d00c000c0c00100000000000040c0c000c3c00050000010c00000400010300000004043c01100404000000000400030031071000000000003000000000000f0000000001000000000000000c0c0001000c0440030c0000000004000c00040c000040000c0c000c010000;
rom_uints[29] = 1024'h1100400000000040030030000000030000100310c1005000000010c00310000000c010004000c00030000010000003000000300001004000007000000030d000000001000000000010010001000000001100000030c000000030003000000000000001001300000000040030000110c040040000503000000000040c00c04303;
rom_uints[30] = 1024'h4001400030c04040d010c00d10c00000000103c0c0404d0330c40000ccc000010003000031c00c000040c0004443501d00c0c3f000301000100103c000c04000300040c03040003c000000c04000d07000c000c0f07c00f0c0000c44000040c0f050030044413003c040440000c000000000c140f040c0f0430500403c0034c0;
rom_uints[31] = 1024'h30000d000000000000001410000300130010070103c10003300c0000030010001d41043100000c3000050000343000353004003000300000030003010000000140040c40000000001300000030c304300004000000000000000000003100040000cd30004100100043c001030010c001000000c000003035c300030001004000;
rom_uints[32] = 1024'h40000000c40040004100cc0310c14300010140c40000c00d0043003044010000000d00c0000003c1000d010003000d40100403000000c040000040404d0300c0c00000c000c00100000003030001000001040000000000000000000003c0000003030000c00000000403000000000000040003000003000000070003430000;
rom_uints[33] = 1024'h4000f140010c00001c3c000000d07f00141000130304401400140401cc030003301c0c3c00340000dc03000c00c01000104c3034050003c3133c000013000c0000c30c0000c00000000400001c0040000450300400001000441c00c04d0c3001000400000000000400700000300400010c300cc00000000540003c3014c0401;
rom_uints[34] = 1024'h4000100c010000400000000100003000001000c34c03000c0000000000110340c0104000334000c01000000030310000f0400300d10000c0400005000000040000000f00404401040000001000c000300c003300001110c03000303000000110c0707000100100001000000040000000000030333c0000000030000030010;
rom_uints[35] = 1024'h1c00000100030c1300040404000c000044000c0000c004000000340000300400004c000000300000cc00000c0f43030c000544040c0c044f040c1c0c0000000c040c04300404c00c0c00004c000c0c00030d40040c04100400000c0c1d1004000c10440000370330000c000c0100050000000d0100040f0043000f04041f10;
rom_uints[36] = 1024'h1000500040c0000001c0000000c00000c0000000100040000000000000000000003300c00000000000400000c000010000000010000400000000030000000003000000c000000000000000000000000000000000010000000000000100000000000040000000000000c100000000030000010000000000000003000;
rom_uints[37] = 1024'h3004c0f400000c0000004000c0100c003040c0f43040000000003c0030040c00c00000c400000100104400c50c4cc0010030000030c0004c0f00c0000c000010c00000700000000300c00405000c40000000cc00000014000074440c3004041000000c1074000000441d00c000000000040040c44100c040010040300c1000;
rom_uints[38] = 1024'hc000000030cf0100400000000040004000000000000000000440c300040c000010000000010010c0410c44040c004c0400f4000000c00400000000004000400000d000000000000044400000000000c000c00040c000c000000500000000cc000010300410000400000000040000000000100030040c00000000000000003003;
rom_uints[39] = 1024'h3400c00400000001000c01000d0000010040100000010000c003d0c130000000c004001401000c0d000000000001000003000000033010c0300000314004000000000000c100404130001000003400c30000c0000000000000003cc0303000000c7001000010000304030003000000c0000000000000300030000303000300;
rom_uints[40] = 1024'h400000000300000000000c0c000040400cc04100000100c3000000c1000000400000000100c0004400000000000040000c00c000c00000004000404000000000c00100c00000000000000000c000000000c30000004000000000400c00000c4000000040040c0000000000000000400000c00000400040000000404300c0c;
rom_uints[41] = 1024'h5030000000c0c0040400000034000004c00000000c00000cc00400040c0404000c0000000004000c000000400c00000c0000000000c0000300000000000000cc0000343400000c005c0004400050001000000000000404400000000c0000300000040c00000000c0000c0000000c300000000000000010004000;
rom_uints[42] = 1024'hc0000004000000000040000440040d00000400000410040700000400000000d0000000400000000004000000c00c004000000000c000000040000c0004000000000003000004000300c0000003000000000040000004000000000010010000100000400000010030000cc0000400010404000400004000004004c0010c404c;
rom_uints[43] = 1024'hc4000401010400cc140c1103100331100040300c100403000010c40045100cc40003300000000034c30000000430003000004d00c050000100304001c1040c0004000000043c50000c0000c74000300330000001000c0000001104300030000cc40030030440030000070cc00c0030c00c41004c04cc400700010400c0cf00c;
rom_uints[44] = 1024'hc0000c0c04000c1050c0c00000000c00000c0030c03001c4300000100007c00c3300000c400300000010000000000040cd00c004c4000c0404040013c0004c00000c00000c04c0000004004c00000040000c0000040c000004000000c000000044000004c0c04cc4040000000000cc0c0400000c0030000cc40000004c0;
rom_uints[45] = 1024'h300400000100010000700300c34031c3400400000300000001c3000100c0c00003010100010000c0034300000000000000400003000000004040000001400100000000030000004340c0100000000103004000010301000300500000000504000003400030000101300000000040400000c000000003c0034004c000400040c0;
rom_uints[46] = 1024'h10001470c0000000070030000404000000c4503c010c00000040c0000c004000c000c40040c0430000000000000000004000004001000d000000000000001000140010000000040000c00000c14000004010000cc003000000dcc000c00000c05040500000000000cc0000033070040c3010000000c040f030c00403003c;
rom_uints[47] = 1024'h10000000040000043c10000000000100003c0000001c000000040c303c030c0c003c0000140000000000300000000c0d0000000c30030000031004003c0c0000040c30000030310400000000003010003000003c000c00000000000c00300000001304001000003c3c00140004303000000c003f00030003001014000000003c;
rom_uints[48] = 1024'hc040c000c040004000c0000000c000000000c0000010400000004100c300000000000010004000c1c0001000000001000f0000000304003000000000004000c003000000000400000000004000c0c00000000000000000000000001000c0000000c0300000000040100000000c00001c000000000000001004000004000040;
rom_uints[49] = 1024'h4000000000004000004000000000000000000000000c00000000000000104000c1000040000000030040000100000000004400300000c000000040030000000010400000000000000000010001040001000000c000300004001100400040001000001000000000400000000000000040040c400000000c00001000000300;
rom_uints[50] = 1024'h1000100070041c3103011c030d000d00000000071300001400100130000170433003400000c0000010000100400003000003100030013031010c4003000000100000300c033330000011100030100000110000303000000301300340000000000000300000000010000000300000043010340000000007000133004c031;
rom_uints[51] = 1024'h3000040000001000040000000000030000c000000000000000040c0c00040030040000000001000000000000000c00000003030100030300010c0000000340000000300100010c000000000010000000010000000000400000010000000000000000000000000c00000000000030000000030700000010010c;
rom_uints[52] = 1024'h1d000c4070100c000000000000001c000c0030fc0400004404c10c00040030401cc304000000cc010034400300cc00c00c140034030c0000100c0100000000300c00000350000400000000030000c033000000000004000040014c00300050000030010400000000001c04000400070c000030fc00300030c014030c;
rom_uints[53] = 1024'h104010c00000000010303c041000044000000004f010140cc0001014c00c0000c4c0541334300000000000003c0000040000000c00cc000400000c404000043000cc1c00c00400c0000000000c0c40000000c000c000003c000000001015c000c00030000000000c000004c0004c0040000c004000000040c00404040000f00c;
rom_uints[54] = 1024'h300c00000000000003030000000000000000000300c400301411040000300400000000000030000033000c300400000000c0000003000000000001400003003c000000010000cc000000000000c00130100000000030000001000000001c03001000000000040004000000001000000000044f4000040f0414040000000010;
rom_uints[55] = 1024'h5014003c4030040003440c000f30107000c0000c0c1010f0000407c0f00c00c0ccc110000cc7010000000001f40003400d30000000c000c01000040c4f13000c003c1000c300c00000003d0001c10013000c0100010000c0000c340011000300c0004000100000c0cc1100c4047300000c3000010300f000100035100400003;
rom_uints[56] = 1024'hcc000004000c1034c07070400c401000100c004000c00c0003c00000000c30003400140000000010040400c0c00c00100010101000300000100030074040100000100000c0c0300030004000000011000000300000000000005000040c00000c00c400100030031c0000f00030c004001000000000305000000050c400000030;
rom_uints[57] = 1024'h4f50400040047c00100000030000001000000000c17073ccccf300c0c3000000030001007000d0c031c0100000c00d41003f001040d300c0c04cc070410140001dcc00000000000170040c0000007100000100000300f0c000c0c33041303df0000010000001030000000000100000430000000040c0f40030c0c0c00300c0c0;
rom_uints[58] = 1024'hc40000004034004000c001000000400100000000c3000400000000c0c0c10000c00c400040000000cc000000000300c0000000000c000000010000005101000000c04001c00001000140040c0000c0030000000c000003000c0003000400000400c000000100000040000440000000000000040040000303c0c00700c0004001;
rom_uints[59] = 1024'hc0f0017000003001013030000010000010000000000000000033300010000000000010100041030000053010035f000030400033000000500401003000004000300300000000c0304000c03000000000001040034300004070100030000030000000d00040c040010000033103030000701010003010c03001100003100c;
rom_uints[60] = 1024'h4000c010010100000400000403000000000d000000c0d030c007000007000000000030000103000000000000000100031000000300000004400000c3000000000000000000c00000000000000000040000000000000000c0014001c00000000000c00000000004c0000000f0000030000040000c4000c000000000;
rom_uints[61] = 1024'h10c000c0c01000004000c0c00030400000000000c0c040000040cd043cf00000300000000000001cf0100003c00030000330000000c04c00400000c030300004c0000030000000c0300000000000400000000c00030000000000013000c010000000c00000f1c000414c000000c0000000000000c040100000530c00c0c310c;
rom_uints[62] = 1024'h1350f0000c00044000003c001000440000c0103000101000000c0000300c0000003003003030000c000040000c000400003000100010000010c03035000000001c0010000030000000400000505c001c00000000c01000001000c00000003c304400fd3004040004c010303100c0000400000000300000c010003c0000000000;
rom_uints[63] = 1024'h1000004040c0c00400003000000000000540000000000000033010004c00000c00300030c07000000000c0000000000004300400c00000353000000000301c0300c0000000000000000000003000010c0000c001300030400000100001c4f00f30c000101000031000430000001f30c0000300005010000030000;
rom_uints[64] = 1024'hc0000000000040100000000030310000100014000404c000030000500c00c0004010100000003000c00000030c000130000000d53300300005c000040710000c00330c000045100004100003430500000c0000000000000000000001c00000071001000503014000000c0000000004000c00c000c4040300000c4c000c04330;
rom_uints[65] = 1024'h7003003000010003000001000030130340305030000d3000000031cc0c04c0040004030c3000000c13003000000c031300100c00000000010114000100400c0003003c1f00c0000c4c030030c304500030110000040c0000040000007000000001c1001000fc040003000c0000003c30000100f434c000c0000000d0000c0000;
rom_uints[66] = 1024'h43000c000040c0000300d04000c330c113f041c0c4134000c010000040c0c30100000340c001c100c001c00c3131003000c040400c030404c3411000d0000000c0c0cc00c0c004004000000d010cd10f0100400000c00001c1c040c3000140000143c403033100000000100303c00000040470c03100000030c000ccc000cc0;
rom_uints[67] = 1024'h3400310303fc0304000c03c10350414000104004000000000c0300030143000003100000c3000d0003cc4400c0c005310cd300c0014071000001c01301000000000000000300001050004c00040500c0c340c05003c300030340000000000000000c1f7141000040c000c00430030003c0000cc4c000000000c1ccc000430107;
rom_uints[68] = 1024'h301040004000d000043d74005404c04cc00000000c0c000c0c100004d0000c0000c0404c144003c0fc03140000000040003040c3c00cc0c04100030f00c0050050000000040000d014000000044040c04c04004030403000504004000000010304400400d140003000f5100030000000404cc10c000000004000c47000400;
rom_uints[69] = 1024'h310c00c4000010010000130004103500115011040c0c300f00d30013101f00040730110004100f0000c4003303035c3140d100300000010000701303511d0700703000000030001011303c00031c0100c301000000c000034040000040d300000300003030033f000004000030300003030c000c000c00030c00033403104101;
rom_uints[70] = 1024'hfc00003004cc0300f0c000c00c001000003f000034f0133003003c40f0303003100030f0140030300000000044400000c37400f00010c03c3f00530030f00000c000f07000413003500000004000f050003cf0000330000000c0104000440000c001c4c030c01003001370000030400000000c40100000304000007001500000;
rom_uints[71] = 1024'h4100000040c0500000000000cd0000c0f1030030c01001c00000c100003000000300300001000430c400440c010004c4c0005c0c4000c0041000003c000000000000314010c000004510000040c100101301000000300100c0c03d0040000000000000033010030c000000000003034000170000000031400000040000100;
rom_uints[72] = 1024'h3007c00003f300c400100300004c4003004c30000303000004000000004000011c01030d010f0300c31040c00c000030003c00000000000333f10c00000f00000000000000100000c0000000000403010000030000000003004140000030714000000000000001400c00c00100000000000c000003000000000040c000000000;
rom_uints[73] = 1024'h30f00000441000300541cc00001401003000300037c43c00c030333040fc00cc4c3300104c30704000303c00f0304400030074001c30743000000070f400017004f03400000034d0405040c030705000703404703040404040104c10c0000400301c4035045c0004143050c0000000f03044300040003010350034000c1003;
rom_uints[74] = 1024'h410000c001000c10000410071010000404dc1000330040d000f0000003300100000000c00000100040d00c00d13010403100040000d000c3513003f3000000014010310341010000000010111031000130003400070300c00010300044cc03000000000010c014040130005000300030033400cc033400dd14000101c010031;
rom_uints[75] = 1024'h4000003300000141703c30c00030400000c44c0c04345000303041000040f0703000001031100cc0300000003000350000301530300031001005c0070104303000304103c0c00100004050f00003000033300000100000000003000c01c041c330d00030303000000000d0000003700040004330100f71410000c3c000;
rom_uints[76] = 1024'h3c000c00000f50310003c030001c500000044c0040303400040400300c3000030c003733100010041c00001f07140030030004cc07000c3500000311050c1000340535000030c1104c030c1c0c01030000000104303003105c4303000f00041fc00310013f330c0d00013f000c1c000314c40c071341001f0d030003030005c;
rom_uints[77] = 1024'hd00c00c00000c40040030043000040104000404110c0004000000cc00000df00300013c0000040c0000c011000400341000700c40400000000130047000001c0c0c0000100440c000400000400000000430000004000c0000340cc000c000f0000000000c0c004000100004000030f00c4c000c00c000c4300c00010c0c0;
rom_uints[78] = 1024'h1300c370c3305040c40000c030040000040c0000030d00fc1040000700030130cc1300004100cc00c030000c404700003000c00c3000374000c04407143100d0f000033105c00700101c01100000c000000300c000300c0003300c0310303c00cc000100134033030d001c4c0007c0340003cf007001010000000d334c034;
rom_uints[79] = 1024'h4310003030f01000144000003030011000d031400014000000c003300040d01013304130000014c0003033030030d0c0001003043cc10000500030004040000400300011100000004d030130000070c00000040000c000300000c0c04010d0c4c00400f044c00cc000c0003000f300000004c1101313c0140004110030003050;
rom_uints[80] = 1024'h33000000000003010301000301503001040000003050c1103001cf0cc0043001000300140034000c333003c00c0100010f00033040000030000001013400004f033033030000031000000030f003100f000000000001000c111000500300c00000c030303010100310041d3000000c000010c0030104000000000000c100c1;
rom_uints[81] = 1024'hcf110300040300010f1713001000030040050001500000310007000104433503000107003037c010051f0040001d3dc440050004300c330d0100001531000c1c000f00004cc000104304c0350400c31df310000100010d00c0300000030110033c000030cf041d3003000c050010000143130007030000030004000003310c00;
rom_uints[82] = 1024'h30331c13014c10c0000000000001001000000004110044004cc000010100010400401c30001000040000000c0040003000040010003000000c0000c0000030500000000300003030c0000000010000000300000004cc000000001040000000000010d00040400000000000000c30070000c00000000000c040;
rom_uints[83] = 1024'h3100000f003cc000000c300f4ccc00043c0000010040d10330000140300404001730000cdc003070007cc4030f1c0440304f400cf04f00f0c54000c7ccc1cc00004c04000404000dd00003c000c04143c0010001cc4000000000c0c0cd034000c000f30001c043003c43000f00ccc0c00c300000034430070330c0040fc30c00;
rom_uints[84] = 1024'h40374000044000000001300030c0c0000c30000c0d00c0f0c0000000000001000300400000101000000400000000000710000040c01c030110c300030330030c0c0c0403c01300700000005303140303100000000000c00000c00000500000300400000001300401031100030000313000c0300000030000c003134000000;
rom_uints[85] = 1024'h70cc1cc0311000014c300100305f000003000034004c100c400003000013030003401000c50101301f300f0c40300100000304cc1510c3330003000100030040111070010403401000410c000131003311f433f100301300f035041f03c10000440010001300003343000000030c3f00c5017c003530300c000000dc104001;
rom_uints[86] = 1024'hcc00370cc311cf00c401011001000141c401d0003f40000000030f43000c34035c303c0303c04403004d00004d4304c500030014fd01f4403300414007fc303000c000070c303130c00410034f3030100cc000000400000001c41400dd4f4000011300c031c01000c40c3c0400000000100310c0034000010c30103103004303;
rom_uints[87] = 1024'h400c000000c03003c00001400300000040c0000003d300c0041103000003c13041d0c000c0300300000344c00300404000000000000050101000330001004001ccc0d0cc0c0000c040f1400005c03140cd4000000000c001300000c004c0d04303c30070c001001000034130400000000d0001c043400300c3100341007001;
rom_uints[88] = 1024'hc3df0cd00010c3c0001000000c70c700000000350c040c0000404c00c00c0000c0ccf000f000040000071004d10c0300c143040003030040c00400c030340000d000f40000000100c3c01c400c00c0c40414000c00c000040c0400c0c000000f0330134300c0c04040f0100300000011004044000c0c47c0c1c100c44c13004;
rom_uints[89] = 1024'hc00100001040d401c0001000000030d3043000300400c00c04c00050330400003010000030000000d010000000040c133c10307014000c00f0d00400000000304c7000000433000000c0030400101030100000000000000000300010c0103033000050100000033c00f0000000100040003030c0043330c010c0c40c1400000;
rom_uints[90] = 1024'h10000c304000430003454170d040c0c1000334000001f000c000030030c403f3f1c0c30033f001c100d00c04010000000043001030000000331000304340c4d0000000d343100040700000003c001000001000c00003000000000000c0030000c0c140301533fcc000f31100004c030c000000c3330011cc00d000c01140c003;
rom_uints[91] = 1024'h33700034003100000000710400000f000c000000000d0400c0710c1ccc000000070c40c000c0003c0303004000000000cc0c0030000c00c04cc73140000d003d40c00140c00f00000740410000000fd4000c00000000004001c3005c07400100000003c0033c130003300c0400000000043cc533000cc00c043d0100ccc00000;
rom_uints[92] = 1024'h1300033000000030010103000000010401000003000000003100c0c00004003350c303030440034510c000000c000000040003000010003000014000040c0010000030300001000003100000100403000000003004400101410040c00000000d0000000100c0000003001303000007003003003c0000410c000c0d13014301;
rom_uints[93] = 1024'h40000300c0130000000001c001c000cc50000000000f44000000400340410d0103040c130300f310f00004400051c0040000030101c30043000000300c03030000404453040041300400000073000cc0400143100000001010c0011000c00111040000311100000100040c00c00fc00300030003d001040003c000f000030;
rom_uints[94] = 1024'hcfc4c0000fc4000dc3cc44440f010c300000301c00044c030c040000c3c000474c000310000ccf00004c03034400f0dccc043fc00cc0000100003700c0c40fcc0004000104c00cc17000000400100f00c3000d0c1c0000310330c4310344030c0030000010134c0400440f00030000010003c40c0ccc1c010f000503103c4cc;
rom_uints[95] = 1024'hf1300000000c0030040000300c0000c0001001051100010000030400c0dc000c00403400000000f00d0000007000440000c00030031030c0040040f540400001303c000003000040110030030330300000311010fd0400004001d00030003300000030004040c000000000000000000300000000c300003100300000300000c0;
rom_uints[96] = 1024'hc00cc104000000303000440cc04001300030010000c0c0c0004040000c340003f000030000c0000ccc000000c000003d40500030004003c073ccc040404cf70000c0000001c00040000330400004000cc000040000000000010000000040000040004000f0300c0003c0c000c4000030000030c3400000cc0410c4c00c030040;
rom_uints[97] = 1024'h4d14047f050c0004003000c00f000000c003cdc01004430400d010340000dc301d00000c30071c0cc33c000c700000c00001010005c0c30cdf00041ccc00000104031000100000030000000000c00000c34000000c130000070000f070c00000c04400c303c130003040000c0000030000040000d010301043004c0040d07c1;
rom_uints[98] = 1024'h40340130c03000400000000100100000003010100000040000f41c070000040f001300000030013030000c04000014000c30040730005c040300100410100000400c0004f10000000003000300030c00031000403c0c00004100c003400404c0000c000000000000c3340c00c0c00303000101f33333c4000c0c0000000f0c00;
rom_uints[99] = 1024'hc0cc0cd300c004c000c00c00534cc4000040f005403c000c04c03100c10071000044f00c0001c0300c00300100f0303004c0000053000044310c00c44000c000cc30000c100000000000c001040433c000300040070030003c300cfc0010f4030400d041300f0c404300f3000010001004f3cc00c53040300030003c0001004;
rom_uints[100] = 1024'hc000c0000004c00400f4100000c000103000414000c0000000c010440030c04000c73004c0300f0000c0000400c00001c000100000440000400100d00cc0c0000c0334000004030000000000000400c0000000040300f0000005c400c0c100000300004000c10000000000000001c00700007100f04505c0000003041;
rom_uints[101] = 1024'h40037d0004ccc00c4dc004000c00c170c3c000004404cc00c10044c0034300300c0f1000000340040dd440001400044004030c0000000000c1000c000300000c4007000344004c0c00000c0000010400400c000c000001000004004cc3000000000c0000030101c3c4c110000c00c00c0040074c01040c0ccd00054000c1003;
rom_uints[102] = 1024'h343000cc3c00140c043430001100070004100013000010004000040100000c03101004000c0000041000000000c0100000710040300004101c34c001000000000c00000cc004000c140040000ccc0000f0000100400003040c4007101340300400000000000010000000c050c00000001c0040c0040000c0003307cc001c000;
rom_uints[103] = 1024'h4303000033c133041c00cd0001000301010c000003c00000001100000c45030300430d100000000000d30303000400010c3c003101c041c5100f01cc0000000300004304070000cd030101000300100305000051000c0f0001c030000033000000c0000310010110c00300003031000c0331043304f10300100007000000010;
rom_uints[104] = 1024'h100c00f000c00000040005014040114000000000000050040030c030f03c00003000d04040c0c5000500000430334040010000000c00100c1000003c0c004000000cc0000004030000033000ccc014c00010005001000030004000404d40c0000003000010003040c04003400000c00000000c00c0041000010504000370400;
rom_uints[105] = 1024'hc0003004003050300030c1c400100004c0c030000c0c0040103c305000000034f1145c043000010c00500000500cc000005c00c0000c10000c0cc0ccc4003000c10010000100100034f4014000405c0004c0cc100c100c01000c0f040150000000c0c004c0000000404c0c000000c0c000cc3000340400000100031044c00100;
rom_uints[106] = 1024'h40003040010700000d000034c4d04044c0c0c700004c030030c040000000300c040c000000403000c43030004cc00044c4c000000c100300144cc0c7c000c4003000300300000000000000004000030000004000444000cc00001c0400400000004004000d4400010010000c4040400000000f433004103c00110c4440c0004;
rom_uints[107] = 1024'h4c000040130010c00c1cd01c403c341000301000c04c1c300cc1003000100000400034000010f00000750c0400703400401004100000347f0700005f10544000310c1434130400fcd0c0003070400004044f043c50100c00011d00000043d000ccc400003400100c30f0700c04300040000c10001000007c3000d0704001f050;
rom_uints[108] = 1024'h3000310501c043004000000300cc0c00000ccc04c43100400001003c00000c3f10cc0c030007303034040004000c0400c44c0001cd400101000343000170001410000cc4000f040c0c00000011c0000014040cd500000000570041010073000c00004034005c001003041f00c434010003000140c3c0033c0033c0054c0401;
rom_uints[109] = 1024'h343400010c010000000000011300000300340c0000000003000405000043f0000014300100000004044f0104001000300043000500000000c004000400040c0000103030000000030c040000440000003000000031300f00000c10000005000100000000033040000100300000000000010001c10103000000c401004c003000;
rom_uints[110] = 1024'hc00430430d03c0c3303f000044500c01c100c53fc1100003000dcfccc00003000cd0344007c33d0004040000010c03013003c00004000dc3000003700103c3c30c00c00cc30034400f310c003014410f1301000c0100c0044c0d0051004c0433070000dc0140000040c430074000041f0c0dc00cc003000fd000c14044000;
rom_uints[111] = 1024'h10c000000700c3004cd443041c0341000c3c303d171c1c400044003c301f3c0f103ccfc0040c041430f03000304340cd30c3700c044300003fd40000fff40000c00cfc31700c0000d40400000030c000cc30003f0fc030700404007000001400400304001d00017c3d04000000343c300030003f004c000c5f04044cc74c003c;
rom_uints[112] = 1024'hdf0040c00003c00000f0f5010004d0340040000000030000c030407100c000c0310010000000340031c033d0044c004000030040c00000c000c00440000f00f0c0c0cf4c0001c53000000300400fdc001304000430000000d0c00035d030c000047004344000f00010000000507000305f3c40c0403400c400c00004c0310070;
rom_uints[113] = 1024'hc04000000304cc403000100007030000004000005000003cc043c0000003701000004d00000333045ccc0c0400cc017303011404003030000043c00003030c330404c000400000000c00040000100000030400000001c00041c40050010000000000cc30004045000040c104000300000007443c004000005130401d075c0003;
rom_uints[114] = 1024'h30300300110c0300000d1100010134300010d00004030000300001d03001003007300404130700300000f000301010f40010007c010c000010300000010100003f300cf004410011c70330c1000c0000030000000d03c10043010310040040000030000000013000110300310370303010700c5000100030037100033dc00000;
rom_uints[115] = 1024'h100c000000300340000141f0131400011003400000c040300300c33c000c1000f0100c0f003041011000c00000300310100c00000070000003504000141334010c40c000000043500000300400c000003010c0104003c0010000c0000003330000004010500fc00004c30d000004700007c00003330100d07040000030000103;
rom_uints[116] = 1024'hc00430f01100c104410c4011001d103c003010371c00303c004330000031300013004000000337c013330c01007000d0000d0037c040000030cd0314110401c0003430471030c05010000010c0000c0000c1003000f000300000014000c00000033000000f3001c0001030d00000000100c0040d00000030c0ccd073c0103f00;
rom_uints[117] = 1024'hc70000000c0000144c0000cc004003000c043000070c144c05440440004010cf001411000f00304300000341000400300000c0cc040440c00004001000000000100c1c000fd004000c0000000c0c0c000000cc000c0c00cc0005c3010000c0003c0437040000001000c000000040c0000001000d0c440000000070010f0c;
rom_uints[118] = 1024'h30d00010000103105340100007f30c000400000030c0303054c03040103001300001000000f0100300000341f400c000410000000000000100330003000c0cc13cc000030003300000c0400001c1000c00000030c0043430301100c011131073000003000000005100330000c04333300c070c4000001000d414310d343000;
rom_uints[119] = 1024'h100401c004050000004401730c0f003000c07c040c001df00fc0100c0000340f0d0d0c000004f41001fc0001c41003400d4307c00cf44000004fc41c0c4304040000c0cc030cc04c40c00c00c70140030050010001000c0f030c041c0c00131cc304030300cc0c00c0000d000300000c000fc0000000c0000050c10000400c3;
rom_uints[120] = 1024'h300c30000001300343400001000141000000003c0c34f000030000000003000c414133003010300f0c30c00d0013015003100100030100000030003400d00000010100000300000300043000c0010000010001000000000005000015000000000043300000010000000c0030000001010004000003000c000000000d0300510;
rom_uints[121] = 1024'hc00000000004103040f0300004c031300000f41000500c0c0c400c10004000047313d0043070f3c0cf00043010c00004031000000c400c4000d0c45400043300003001c1700403f0f030c00040401000030cd3100013000000300004d35300c434310010f0001000c0c00030c0000000003030f00043740000d00010000c013;
rom_uints[122] = 1024'hcc00303040000100c41c340000c0030007003000300040d01c040c100300c0330c070000c040c100c30003003100003000000030000300ff000010140000004010000c300c001400040300413f70c07000003c300000c000000004000040f0c00000c3040100000c0030c440000000404f330f003000043430000005c01;
rom_uints[123] = 1024'h100704c030cc0013040400004d310030300013010c0433030030033c0d0c0c0003011c30140300430000dc0c013c003304dc00000c030010000033000004040f050003001c000004cc400000070c00d0000403303004143000010000440c0000100d03050c010140001c0013033c00040100d30001010310000000cd00c;
rom_uints[124] = 1024'h3000000c0140c00040010000040400341000000000cc010000400cc040040300000300100000700000f000310000500304c001000000040f0070030004000000c0030003003000d000003300c100100000c00004c000000000c0000030000000003001000000f0003001100000000003000003c000000040000001f300d00000;
rom_uints[125] = 1024'hd00030cc0000c0003000c0c00100440001c00000c0cc400c0340000100c03400c00030cc0430101000043000c0410c4040c0000004c05c007004c0c0300000140c00443030401c0000000000c00340043c0000000330000400c000000c0010414050c0004000c000430001c700003030001044f00c0054ccc0500003c0f0103;
rom_uints[126] = 1024'h133cc30cc000c00c30dc00c010c44404c030000000001000c071003c00dc001005044300500000004000000040410000c430004030001400000000c1c003300040d0030f00001043000001013c00c3507000c000c000000040c0c000003c00c00010c0c0c00005c0c000c04000000000400040003c34100000000040c0000040;
rom_uints[127] = 1024'h3004104d000000100c00000110cf0010143000410c300010000300000310303410101d0003000f030300340000033000044000351300000c0000001300007300001003300300140043000400033000000000000400007033010000c000013100000c030030001c110030000000000f00000000300cf0000001000000040c;
rom_uints[128] = 1024'h10000c30000000000000c000130010100100c000014000300c00f0f000f000001400c000000003000c030000000400100030004000300040c0500330000d0003000300c00004100c00010300340001100001000000000030100040001005000040c01c0000000400c040004000004030300c00000004400000c0000000c00000;
rom_uints[129] = 1024'h74000031003c00343000000040301f07403c4000003134c000c00dd000300070c000330c0c00000000000c0300030010041000303000c401011300c0104c0c0003303100310c073c40003300ff0c1c04334400000400001c0004c00070c0000400c00003003c040400c00c010000000030000430f0010000044000000d000000;
rom_uints[130] = 1024'h40000f00000000033004c33000c330001300400cc0104c00c0000000c700c300c00043400000cd00c001000cc0000c0001c0010300003000c0400030d0c00004c4000000c000c0034000c000100c110cd500400000c3300400c07003400100000043c303400c00000c40c0cc030140d3010540c33101000030004100f0d00c0;
rom_uints[131] = 1024'h70033c03c333c3000030030c00004d3000015000003003030000100340030143cf1004c0c0004c0047007400c0c00301c0c303000000410000010013404100004001000003c0000000040f04000030c000400f00c3c300030000c0c040004030c0000c710d01d0000000d010340000c0000000f0c00c0100400000c00c030000;
rom_uints[132] = 1024'h4403c1003004430c04004fd00000414044cc010000c500cc00c0000c07510000c0003c0000014300000fc10001000305004c0000030040c00f044c403c000c000000000c00cc4c310101500000003004c0440000040041000040000000000000c00c47007131040000003010100700000c0004c3000000045100000f00000000;
rom_uints[133] = 1024'h300c300441000000001000c3d450304040101040001c0303000f00c0c0000c05f7001d0000000c105c00c03003300000301000c0000c3003100307c3011c040c310300100030001c1100000307000100000100000c010310010000040010cc0000c010000010f003000301000000001f0301c00000030300031100303010700c;
rom_uints[134] = 1024'hcc000c00c0000000c001300001000040f00f003004f0103000007000003303c3000073303040300070c04001054003f0000401c03014303c3c0000c0033c40000000f00c0000013000c01000000030130330f00000303031000310750003c0c0300000000d0c10030010301010c000030000c0030000c03150f100400054c000;
rom_uints[135] = 1024'h304000400050f14000f0001000cc040003f0000300c01001c3000000450000010400000000cf000140c3c044c000c000c5000340300500c00000f1003c00000040000003000000000000103731000043001044c00400c0c114f0c4400041d0c030000000000050f34c40c0003300000c400013000000c33003000304c070000;
rom_uints[136] = 1024'h3c000000300000310004c10017000000c3c10003330000040c000300000711d0133000d0f0740c01000000c010004d13f0000070000c43030f000c0030010040003000010c0307c00000011000f0000030301000300000001700001007040c5500000000101010030d000000040030c0030c000000001010370c01300c000;
rom_uints[137] = 1024'h400300400040040300001300000130130300c3c0d30143304c0000000004c04c0703030000c010070c00000001040470000103400d074303040100c003300004050307030c00004df004030c000701004303004300000004340503013d0000000c4100030371c4034d0300004c00030007040300040003010050030c01c0003;
rom_uints[138] = 1024'h400000c30400cc10000003301300000040101030400050d00c00d4c00300000031cc40000001000310c300c0c03000303000040000d070c340f00300330130c17010000300001c004000000000c0700030300000030010c00010303043fc0000c010700040000405000000501030303c10000c0c3304001c14300000f010031;
rom_uints[139] = 1024'hf003000c00003310005d04303d00c3100000000015000300045040300001d3000cf0030010000045d030c0300004000000000000d01030010430c01004c033010700c000300100000001000000003c0000000d0400000010c7f70140c34071010041c0c0f00033000050c1030010000073714140005000500351410cf1000000;
rom_uints[140] = 1024'hc00040f10000004303004cf30001c40040404410f1030400403000000330030334001f0301c041c330c003f13c710004103130000530000353c30130001101000f00030030000000031070c100c01370004000000c10003044403031103000004103311150033000d1371001003dc0c0000000c30100000130d03c03f1704000;
rom_uints[141] = 1024'h100c101c030000000470000010fcc0000004c004f00100001474000c004c001d3c1c1000000c00040c0000c010410000341000403c100c0007c0010004303c00100c000000040400c0000000100010003004000000d0000c1000040c000000003034c000c00c0c3c40001030043000003c404c10300000000440001004000c3;
rom_uints[142] = 1024'h10000434d3304030c31001c430000c3014400040030cf0f0103cc3043003cc00101000c00131c04d00001000300000073000c3003400005400044003100100d1c000030101c01700100040000000c301300000c7003000000330400310000001d00701c0d30c00334c0010300007c03400cc030140c10330300c1cc00cc00;
rom_uints[143] = 1024'h10003330f000001430003c30300d000000004004400000c4d044300c14100f1f304100300054005c30300333f3cc000003c0c00001c000400030104700401400f0001010c0403070000000f0304cf00014c0000400000000c0c0c3710cc100c0000030400000c000c100301030304000d4c0c01000f010c000c00033030010;
rom_uints[144] = 1024'h33000400c70000c000f4003001533000300000000440031010003c13350000000003001400040030000c0f000c000c013000030000300005000c00003000300313300c3000000000000301030003100014000000001030000010004010000000041c303330d0010c10331000c0000010000000000000041001000000000000;
rom_uints[145] = 1024'hdf013000000cc005000410000c40c00740040340101dc031004700cd045305cc003100003000f010010c0c01001d000040101300300300010134000440000c00000c03040f0000c00700f13004000f00030c030000000000c03c53113305000301c00040cc04004000030c050301000100000007c0004d03410004c00031f000;
rom_uints[146] = 1024'hc000c0c73000100000c00000c0013400001000000010000c004040130440040c400010000403400440d0003100404000c0cc3000000000034001304303100300c0000000400000d030000000400010300000100011c00130000c000cc00000003004003000003c000c00100400000000000c00003470c03000100040c000074;
rom_uints[147] = 1024'h31001c0f003000101000400f00cc10040dc51001000cd0373c070170c010040053000d404c0004cc070f040003101015300f003c0073443001334cf70cc5c0004c4c00c0c4040000100c00ccc0cc0113c0310400004c00000433c30001034c000300f00155c003003040700c00c00073c00000300054300013043c040fc340d0;
rom_uints[148] = 1024'h400c0000000000001030030000003c03003430100003c0f00d33303000040000304000050030010000010000000c310000004000fc30040000003004c00c333000403c0c0007000000c00c010000f00000000d00003030103010000003300040c00000100013143d10000030000000000c000100001000000100000000;
rom_uints[149] = 1024'h300f1c003100400c0c0c0044000330004300330430401c00300413000013000003701010c01031371f300c00440000000cd040000004c3300000000f0003c040011c74cd003000100041001000c001000130033100300344c1f10003000d0000030003000341003340003303300c0c1000003d0000c03000010000c003c0c1;
rom_uints[150] = 1024'h3c0c040cc4d40f00004005134f000001c00110000c74d00cc05c3344c00c05034f003c04c0c44000004c0000010f40f4403340c7fc30f40d7330013c340f0c0001f003340c034040c004103033c03010000000000700000100c01031cd034014010011c031c0c000c40c3c043000033010c014f0000000011044103d0f000103;
rom_uints[151] = 1024'hd40000010000170001033c40053000c0040c04003c000000003c033300000c03040c10000c033030c00c040c0c000004010047000000010001000004400000001c0c0c030004000c14030000000013000c440000000140001000000c004ccc34003c30000000000000300403c10010000f0c0000000000300d0000040000000;
rom_uints[152] = 1024'hc0d00000001dc1c144c4004300430700004000c40d00000c01303c0cc0000030c0cccc030034000300034004c10c0c400013011040000041c1c404dc0004c000c300c5000000c10f0cccd0400c00f0040004010d000040045c0000ccc0c00040033013433c0000000cc0c440c000c0cc0040000000cd44f00500c4c00110d04;
rom_uints[153] = 1024'h301c0c40000cc0040c1cc000f3003c10000000301030100c44000c50330431000300c440003400c40c100c00c00000000010307004004c00f00000c0001c0030407005300030c00400c10000100c104000cc30003000000c0f7c00000003c00300c01010000c0f010cc00300100ccc10003470c0043034f0d1c000cf101c001;
rom_uints[154] = 1024'h10000073c000430000510000004000f100300000514030000043330303c0c303c0c0f30300c0050040c00c00c10c00000053301300000000c700010c43430003100000c0400101400000000c00301000001000000f000100c1000340c0030000c0c04c00d50033c003f0d040c00c000f0000030000c000cc331000c00070d003;
rom_uints[155] = 1024'h30c030303150400001010400c04700004c0001030c0400c0400c1c000c40000410430c000c0c3d01c300740010c033c00c0430000000c04c0000000c4d003c40f00c00000c000044304103c00010140000c010001000010000000c14003000000040010c3c040000030c140040000007300103001cc100173d311000c10000;
rom_uints[156] = 1024'h30100c43000c00c0013101030005000000050000043101000000000003003013035000130000400fc500c31f00100003040000000051c005c003100004c50c00130c010030004000c00300000303330000030030300040010000300000000000400000c401000004000001100303030000300000cf3440010040000d03010000;
rom_uints[157] = 1024'h300c40303c40003c00000300df1c100010c000330704044030000400000510cc5400000100cf704500003144000000dc7400003c171330043c10041303c0c04000040545000c541c03010010043f40cc0c030030330000011000001d74000000d000c0ccd151000c00001f000c0c00053c000440c100000c033c000c11cc00;
rom_uints[158] = 1024'h100040c00400c0c00030400c310c300100001f04045c0301040c0303cc00444fc00000c00dc3010000cc50440000cc0c004f040c33001100100773c0c400ccd3040000f00c10f13c100c0737c00c0000c000cf00001130c00304014444000c007c0cd1c0104c0400451f1c03000405c00f07300dcc0030400c04070000000;
rom_uints[159] = 1024'h3070040010033030004000c0504d0000000000410000010000030544000000000430f7144010c03001400030000400c00010c03010d3001000314305004c00003030300000010040000030000000303030011000300010000031c000003003000030c0000100c00010004000001004000300300003000000f030100001000000;
rom_uints[160] = 1024'h300000f40000303d3405cc040000000040300004c0c0c0c0004c100c040004f0001000000004007000300014000c3c00140400000400c0400c007c0c7c030030c000000000004030000040400410c00400000c0004000400c003000c5001000000070030300300041010000434000000d000c300c1c0c00000100004400001;
rom_uints[161] = 1024'h4d000030053c0004c431c0cc4004700000c000001010430404c010f001d0dc0c0c0000000017104fcc4f0c0c40000000010c00cc0400030c0c00300c0000000030031014000040c0000000c0000f0400000400c00003000c040000f04000000001040cc04010c000f04001c030000000000400c000d1001040004c0040c0001;
rom_uints[162] = 1024'h4034c54000c00c4404010400001c4003104410100040440100041010d400040f044f400004300100004c0c000c01500110cc00c030000000470c0cc01010030000010040f00400001000000f0c000000c3000040c00c0c0000000000403401c400300000000000003c344c000000000c00c10030c43300003c0c00000c0304c0;
rom_uints[163] = 1024'hccc0c1713d030000c030031434cc4000443c005404c0d03000c0403f310000000003c03c00100c00000000100c000f001c000005cc43734f00003004040110ccc30300cd4fd0000300c000c0005300000040400043430000070143cc010c3074430c000330f004000d103400040004010c3cc1005344c00f0c4c5f10005404;
rom_uints[164] = 1024'hc000c0400030c0140034d330101103100000400001c1004d00c0140000f0c04030300330c330000003cc40001000c3c1c0001000c0440003011010130000000003033030334400000000004c401000c0000010041030c00c30311400d03003301300000001c1003000033000000001c4000041c00071040030c003140;
rom_uints[165] = 1024'hc4c044c013400c00c0c0100000cc00140c0c10c044401c1000c0c040004001c000c0f0000040c4040400440010400c040c0c00c003000000000001c00030730004c000c00000000c1c001cc0403c40400000c000cc00000c00c07000cc400430c0041c001000000cf1001410c0001000f0040044000040c4c0000c1404cc10c0;
rom_uints[166] = 1024'hc00740cc00c300000c0704000010f034005001000300cd003040c000013351007000310000304000400c0031300c00131004000000c0c1300000000100004c0304c40d01cc004000c1000400c000c0000c04005000c0c00043000001c0000c0044000000300100101ccc0c04400000c01d0310003043100001030030c3013010;
rom_uints[167] = 1024'h30c0c30000100000010010fcd00130413000000c0040000000100011c70530001001d0030370000c0d300730c300070013c0000000000100030c1014141000300000314073300014300300330040003003000017401000030f0003010040000c3000043000101101003c1330000000c000003030430171000114703fd04000;
rom_uints[168] = 1024'h100c003030c0700004010030044350405000041040c000304000c00030700c00004c1530000300030431040430c00040013000c300c0000c10000c000c004041c000c0000c0000004000f040330c0400c000c040c103400010400f701170c0030404c04050043040c5010440000431c000c0cc0cc7040003040034003f74500;
rom_uints[169] = 1024'hc03000300c34c033c03140030004100730d0400c004c50c0c05c440c0034f4105c04000004000054003010300400104f043000000010cc00000104c0000000000003000014043034004040005c0c00c00000005f100c00100c0400400c00000000c0c0000d10030000000400401c00ccf000300010c405c00f141400c000;
rom_uints[170] = 1024'h400030304d400f34c0300004001040040c003700c400000000c000001d0c000304d03000400030cc003030003c0c004414c000400000000c004f00c41c0c04033730300000000c00040c30c003f0c000f0400000400000cc0000cc00007c4000000c000040040411000000000054000000000f4300050010c10100074001407;
rom_uints[171] = 1024'h3f300440070c10c0000fd11c000370c00004d400137c1c000331017003100001400f37000014c0c004401c000c410030001370d40014403c0c4c004cc0c070300040c03010300000d0c004f0400c00c00350003c10034000010c1c0c00031000fc304f0034001000010070c3c03c000700d000040000007cc30c13404c013000;
rom_uints[172] = 1024'hc31000100000334034000000c4300004c03c0003cc3101001407001000f43130c00030c043004050000034040000015400071cc000000c3037000003cc010000403040403c03d000000010cc40400440000c0000000004000010c0000000c040000030040000100c40c000001010c1310c0410710134004030040400000;
rom_uints[173] = 1024'h30340001c0010003031cd0014010000100340c40000c300010330004010000003004000000000034f30300043030000100040c04010000000000000004c4010004500030000003030c000400303000003000000000005c00001c00c00c3400c0000300010c00000000c400103c000100c00000f1004300030104110040303000;
rom_uints[174] = 1024'hf00c0c530430d440003343300010050cc01c140c13cc1000000000103d0030030003c00040034cfc1f1f04300010001104130030100430cc1d001303040c00000030000c110c0343443004003000c00400310000303c00001047000041100000330c43d04c10441000001c74000310104030f0d03000003307310c0c13044000;
rom_uints[175] = 1024'hd0040c04000000000c143c001c334000ff3f00c014dc1c4110141c7c04cf3c00100ccfc0440c0114700df010040040cc3cc0043c047431003fd50404fcf00000f0dc3c4c3f0c054404000430303ccc00003c000f00c00041040414300c001400401f04c01d304d0c3d100d040034c03c430c007f047c001c1014104cc07c410c;
rom_uints[176] = 1024'hd00430300000c0000001313030f0100100400003330310000070707000cc30c331041f000030010000c433103070007000fc1050003334000310c47004030c0c040ccf003c00013c000000c040c0c000100070c40000cc00100000311370c00005043430100300c030000430103003001c4340003c0430c00c0000053c300400;
rom_uints[177] = 1024'h10110004100000cc0001000000400040001000100d0c0433000001c0400040044c01010000005f0000340001003300040104c0000000000cc01007030c03140000000000c0000c400400cc030d00000000000001000110c0c3130010c0004000000c0c000500cc0010040c3000000004040c4040001c0030000c07100103;
rom_uints[178] = 1024'hc0000001015c4700001d1c000001300300c0100000000000010c011c33000330033030001303040f141c30040f041034011d037cc001300014300c373101c33030f1010054103c00c0f3310d01010000000000010d030100403010100403430c00010c3000c003001d031330030d330001707050301000330031030301c00000;
rom_uints[179] = 1024'hc00c00000030003c000500c003041011d0030013013040000040c30003015303c4100c00040051005040c00000c000d010d3000030300cc003500000c01040000c400000000000030000000000300c00000cc0d0404000000000c03000030030c40030001000000373f301104040000044004003300c30004404000000000103;
rom_uints[180] = 1024'hc0000c0011005070400701c3011000c00701030cc307c30004070000130000033040000100030cf103f10c00c000000c0d10c001040000031c100000004c100c4044170143000101000050cc000300400010c00043000400004000000c0004030030401300030000c103010001100000c310001050300f000cc1c33c01440c0;
rom_uints[181] = 1024'h100030030d0040030f330000000c030000043004c40cd05c0005000c000000000104c0cc0f00007000000c01010400010033050f04c44d07000400000000400000000d4400d000c000300130000000c000000030010000c0c005c411000000000c0504040400301000f000003044c00f000c001c1047cd03c00040cd100c;
rom_uints[182] = 1024'h1f00030010c00103000303030034c3400000000040300301001710013c000001f0011100001cc0100071001c41c0c00cc0414013000013fc0001030003330300c10100100c0000300300c000430000c0010010000100440030301000f0101c0033030010c3000c005500010030000141f01f100f000033d03010140d0d003050;
rom_uints[183] = 1024'h4000000c30000000c00410c040c5f040000004c0400401cf40300503f040c040300010c000c00f40c43304000011407700d4014304c34040c574cc41c101f44000400d0f00000004c41c00c00c00100000040000401004ccc0400140c0007031cc0100040330c3c00c0000d000001050c000304000c04c00d0400c03300003c4;
rom_uints[184] = 1024'h340c000334100101001430000000000c00033000001000000000000100407300400000031c010001000071000c100140030131000400cc30041000010100c03003c00003003000013c01000001003000330000000c0310c5000000000000310400000000300300003030013100050000031000f144000c013300400;
rom_uints[185] = 1024'hf00040000040003140c0330000c001c300c3c0dd434000031c40c35000010004030300440040f004f004003013001413c31100040c40cc4030c00403000030c50cc301c5300103c030c0c000003004c00300030003130000003c0000c35fccc03041c400c0310000d00050c0c00000503040050000404000c0d0000003c0010;
rom_uints[186] = 1024'h10300c3c400c41000000c51130cc4340040c3c0000cc41d100c40c40000fc0000000000000341017c0040000010000c000000030300c10ff001f1c1000030c40500000000dc11403010010450f3c004000c040050003ff000000000f400cf0c040c0c304303103f004303c040c4440703c0003303007c40430004c00410;
rom_uints[187] = 1024'h100c0307c000d00000010030304cc033000003030100003003000430311c0000000330000013c00133c010c04031000000040c0030000001000c00030d0c04040f00000c301f100014004c0000040004030304003c304400030001003034000130000c030400041040000c0310040104040000100000c103000100003303c;
rom_uints[188] = 1024'h10070c00000c00c01d03410000403f00400000003c10101c040d00001000c0300c3fc010000000010c0000100c0000304c4000000000400000103010410c00033030000000cc000010000c0c0c0c0300000c000c004010003040011003103000030000001c00030d0000004000030c0000003304c00003034c00000c0110000;
rom_uints[189] = 1024'hc30030c00000f000fc10c0c001c100004040000000c10001c30c30000004f433c0030000040410d0000400001000000043f1000034300c007c1000f00030c0c400100400f000110000100030000030c03c0001c003311005000cc0010f001c010040c0400000c00c4c7000c40030c0300000033400401330c150f000c0f050f;
rom_uints[190] = 1024'h400303007040044000dc0c1100c0000304740000004010100041003000cc00000130330040c0000070000040004104c0c03013300040000040c040d1030f001040c00330003003430043000040030f00300000c00030c0004000c0300000000054000000000011c4c000004000030000440000004c3000d0000c0c00c0004000;
rom_uints[191] = 1024'hf0000405c003c03100c0c0000000f0000040000440003f3d00103001130003000004311000000430300300000300300000000000503c0000c00340010000033f00011c33001010100030000000030303010000000000070330130000000100000000f3000300011110400000000040000000000000004001011303030300c;
rom_uints[192] = 1024'hc00000c1404000000000000000c0c0000100c0c040c000000000014300010040c0c000c00000000000c04000c0c40010c0c0c04000c00000004000c0c00100c0c00000004000000cc0c0c040c000c000400100004000004000000000c004c00000c0c00001c040000000c0c00300c00000000000000040c1c34100c000004340;
rom_uints[193] = 1024'h70000000000000040000000030301334003010000c3000000000010c003400003300000c0c3010303000000430000010001000000000000000000001000c00000000000c000c000c000000000c3410040010000400000000000400000000000004000000500c3c00000000000000100c0000000400000c04040000000cc00000;
rom_uints[194] = 1024'h430001400000000000000441003000c000f03000004050000000000000c0c00010000000c0001004c00cc0001000037030010000004003c00000000030c01000c10c0040001000000004c0c103400000100040030000000500c040c0100000300000000000001003030011004400010050c000c0001040004c0000c14000000;
rom_uints[195] = 1024'h30000c00000041003444c0300000000000030000000100c00070000c3000c00c004030157007400c0100c7000004400000040000031c0c3000000000040000030cc00000000c00003c030000040c0000000104003000103300c0100000000040000c00040000004f0000000000400c0000c4000000d00c300c04007;
rom_uints[196] = 1024'h40c0000004004c00400010000000400500010000000c01000400c00040300c5300313c00000000c0000000040000000004040000050c0300000c10403001004c00000400c004000c0c0000c400000300040003040000040c00c41c0c00000001404c00300c00000400000c00004000000400001c0004400100000c00040004;
rom_uints[197] = 1024'hc0c00003000000000440010001c3340100f10000030000c00100007001c00000400c0000c00000040100000000000300c10000000000000000000000010000c010c0000000000000000040c04000100000c000000000c00000c000400400100000000000003000000000000304c00000000003004000c0c0010003000140000;
rom_uints[198] = 1024'h30000003000030000000c00050c000f000300031d1c000403040500300000000fc300300000033c000000000c0c0003000000040c000c3000001f0f040000003000003000030000000007000c0500030c0c00300000100000040c0404000c103003000000000c0107000c0c0003001030033004300c311001040c3000003;
rom_uints[199] = 1024'h500000000101500000030300c00400000000003300000003000000050003000100000003130c0144000c00000003040003000000000011001104010000300100013000300000010000100700000000000000000000000110c000000001000000003000010010030c000000030000000303000000000703030c000000000f0;
rom_uints[200] = 1024'hc000000000c0030101000040000000400101000330000000000000010044c000f0010000c40000004dc000c000c0000c4340000001c003c000000c4000c0c000c100c0c000400000c0030000c0000000030c40000000004000000300004003d00000c000c0000000010000000000000000c0000043c0000040c000000103;
rom_uints[201] = 1024'h40403003c40040000114c0040001040003000000c0cc0040cd000301c40030000003700f0404000300040040c0000004400003c00000030300c0c0404300000404c00300c004134d00c400004c030000040c000003040100040004034c00c000000000c0030f00030d0000040000034000c0070c00040401000000004000000;
rom_uints[202] = 1024'h300300c10000010300710001000c00000031000003000000000000000000000c000510000000000001000300000000100301000c000001000001000104000c00000000000c01000000000000000000000000040003000000000f00000000000031000300000400000000000001000000040040310100000000000000;
rom_uints[203] = 1024'h10030010030c00000c0000010000000510000001003000000000000000401040c000000000c3000000040000000000000000000000000000c000000000000c001040000003000000040000000000000c0004030010101004100000000000000100000000030003300000000401010334d010000000000;
rom_uints[204] = 1024'h14030030000000000031000301cc11100010000c0004140403000c00000000004c00503410000000000407000000000300000000000c040c000000003001100404000000040100001000000c0c3113000010000000000000040000000030070031103c1c05000000c00100000d00030003010000000f000000000c000003004f;
rom_uints[205] = 1024'h100000300c000c00000044000000000cd0000c0c700004000c000000040000000c101000000400070c0000000030003000000c0100000000000004000c001c000003000000cc100000000000000400000400300000000400000d0c000c041040040d0c00000000000400000c000330000c100330301030400c000400300;
rom_uints[206] = 1024'h100400001000400000103c0400000c000400000cc00000300010d70400003c00001000000030d040c00000000003000000000000000000003dc04440000000130000c00c0000c40010000010000000000000000400000000000f000414000100000000c0003000300104000c0700310010030c0000000000000c000000000;
rom_uints[207] = 1024'h7040000000000040000531000030000100300140004033000010000010401000000c70030000100010303000300000000031000000c00000000000104d00000000003030000000300030000003000000030000000000000000030000000030c00031000000300c00c0304000000000000000000c0000c0000100000000000100;
rom_uints[208] = 1024'h33004000034000c000cc00030100c0000000000004000000000000000000c0040000000000f00401000000c0000000000c00c00000000000000001000000000000000f01c0003000300000000000c0c01000000000010000001000000000000004c03000400c010300000000000c000004040c00c010000000000001c00400;
rom_uints[209] = 1024'hc004000c0c1330000100000040010100000005003c30001c00000030000400000500000000c00310000001001c000000140000000000000034000000000330010d00000301000c00300c000001000000000000000011000000000000310000000000000100000000000000300000501000000000f000310000130001000107;
rom_uints[210] = 1024'h103000000000040c00000c0030000000003c0f044000404c000000000c40c0000c0c000000400000040010000001cc00c00000000c000500400c00000034303004004000000004000f103c0000000c00000000150000c0040c0c0000000000000000000000cc04000000000000000000000004c004001400000044040;
rom_uints[211] = 1024'h1000000c40000000040300300005d0000010004003000040c0030c00000040003c001000400000c040c0000000c0c0100004000004c0000010040040400d00000000c0000004000100000000030410000440000000404000404000004c0400003000301100000000040000300000000007c00440000000000c0000000c00000;
rom_uints[212] = 1024'h40000000000100000000c003300000c0c000000040400000000004000010c400c000100013000000000000001000400000c00300000000cc0c00000000000000030004000400000d0011034000000000100004000c00c0001c000000000007000400000003100000000000000000c000000001004c03004004000;
rom_uints[213] = 1024'hc030001000010043000040400001104000000000000003110000000030300010400000d3400011013000310301000c300001000000101000303c000000000030010110303d000000130300001003000100010000010004000031300000030100000c0030000000300000000010000001010000300300f0000c31000000000131;
rom_uints[214] = 1024'h70000130c40040000000040010100000004000c000c0000c0c003000c004000c140c0000c40100400c3400000c4044000000c0c0c000000f0000004100c00000f0c1000c004000100000000f0000000000000000000c053000004000000000450c00c04000000000000c04040000c0c0c000cc000f00131000c40c00400104;
rom_uints[215] = 1024'h30700000100c0004300000010100c00000000000000000000430000401300000000000000000100003000000c0007400030000010000000004000000040000000001c40000000000c0000000000004000010000000000000101000000044400000030c0c00001400000000000010c0000000000000370c000000100410000303;
rom_uints[216] = 1024'hc00000000040034000000000000000000000004c0c00000000000c000000000000040c0400100000000c0000040400000000000000000004000c000c0400000004000c000000000000000004000000000c000c0000000c00000c0c00000c000000000c000050040004cc0044000000c00000000000000c0c000;
rom_uints[217] = 1024'h40040103001400c0c00300000dc000044cc000300040041c40400cc0c0c00c00c30040c4000000000000c34000000000000304400c300000c100000000f0000000004000c50000c003004f0cc04100c00000400005c0010c0000030c3000000040c000c04000000000000000cc0300000cc0c4003000100003c00040010;
rom_uints[218] = 1024'h30cc0000000040c000c040010100c040000c0000000000030c000cc000c000c4000c0c00004c04000000f0000400430000000c00000000050f0343000000c00300000505044300000c0c00000c0c0000000003110100000000c0000000c1004c0c04030cc000c00100000c030c00c000000c0010cd03001004004000c0;
rom_uints[219] = 1024'h400000000000400000014000010700000c00010300050100000001040c030300000000010000030c0000004000000300000000010000010000014040000000400000000000000004000100000310030c000000010300010100c000050040000001000103000001c00700000303030004000003000001030400010340010100;
rom_uints[220] = 1024'hc300000040000000000005304100c04000100000000104000000c0000000040040040001404400c000000100c00030300300000c00004003c300000300c000000000000000000000400000040c00000c0000030c0000001000c000000000c000c0000000000000000000000300000000c00003000000000000c000000000140;
rom_uints[221] = 1024'h50000010301300000000003001f001000000001131000000003010000001000001003400033403133c000400001c01c40000031130030000c00050c0f0000003011000001030310000440001c0000c00000000110000030000035010000104000010000c0000010100000003000000030000000310000100000000000c103;
rom_uints[222] = 1024'h4300cc04c0000000c300c0c0000040c0001c000cc04040c000c000400001000040004300ccc000000000c00003400c0c000300c000330000000003004c004c00cc0040c00c40c00003c0000c0340000300000000cc0000c00000004140004000c000000000400c0000404030c0000000000c0040c000c0c00004c050004010cd;
rom_uints[223] = 1024'h30300400000030000000000001000000000400301c10300030300003000000000030000003100f04000010003000c00000000300400c00000331003100000003003000000001000c00000000c1050030c130103030000000003010007030301000f00c0004030c000000f500d01000030010000000307031304340c5c10003c0;
rom_uints[224] = 1024'h3000000030000040031c00c0000c1040404c00cc0000000010040100c4440000000100000000000000000000340c0000003000000c00000400100004000000400000000c00001c13000000440005000000c000000000000000003000050c0c00000c000c10c00000001500000c0001040000007000000000000000300400000;
rom_uints[225] = 1024'h301030003000304400700000c000001000400000000400400010003000500000040000d0000c0f000400000000003005000404130000000000100030000010000040d07000000000000030000400040004000004000000010c000000000c030000f0c0007c000030cc00001c300f1004c4100040000c001403c00;
rom_uints[226] = 1024'h300000d000040040001440400000000030400000004000101c00003c0000000001f4010000300c000000c0003000000007000c30001000c4030000000004c00000000c0010300041400000301000000005d00000c0c0000400c0300000001c00000000300010000000000000004000000000003000003000000000000030000;
rom_uints[227] = 1024'hc00441000000f00c00c000f0cc40000c0000443401c700000344300d000000041c3000001000400c0400d30c000000000004040c0c03400000030403000000c00000c00010030d00c000000c0003000001000040040000000100cc414000300300001000000000011f00c00000100430300c0003470ff003001c04000000;
rom_uints[228] = 1024'h1000000040c4300000400000000400000001000010040000000400000100000000040000000000003000003010000500000c0f00c00000003003000111010000000010003003100100000000000000001000000000004013100000000000400330000000000000000000000300000100000000000010000000100000000000;
rom_uints[229] = 1024'h1c3003c403430c0c00d0004c00d0010cc000003000004cc00010014c0004040000c1004000c0000000004300c00c0cc0c000040040040c0c000000d00c40000c30c47000070000400000c00c0400c0004000c0c0000c0cc040000040cc00040030000c0c00400cc0000001c000c0c00300c4c030004000c0c4c00040000c0c00;
rom_uints[230] = 1024'hc00040c00003c040000000440000004000101000000c11000c03cc0c000000c0300000100030030041cc00000000030700c5000400100100000401010400000c04c0c1000c0043000404040000000000000000c0000c00000000034c00110000000c00004000000003c00004003001000000000001000000000c000c000c4000;
rom_uints[231] = 1024'h300000000c000001000001000000c000100000030000000d01c000000104100300001c000004c00700030070000000000c00003000c03000103000010000400000000304003333c140000000000100300000000030000000300000000000000030003040300000130000010303c001410001070000000000333103030000000;
rom_uints[232] = 1024'h1f400000c4c00f00c0400000010014404040005000000130000040000040000c4040000c0000c00140000000003c00114c400000c0c30c0150000040400440000000000000440100d3000000000d40c40410010001c0003000400040104000c03000c000000cc000c400000001000000c00000400000c040000400000000300;
rom_uints[233] = 1024'hc00c033000100000000c40000000000004000c000404104004000c000c0003044000400000004cc00c0cc304000c000004040004040100000c000000003400010c00004000000000000c0c0000000c030000400c0010cc0d003000c0c0030000c000400000000cc00044000c00000c000300000000;
rom_uints[234] = 1024'hc00300000400cc0000c00000030700000003000003c000000000c0000410000d0000000007000000000cc004c0000000000001030040c00004000f000f0400c000410001000403030000000000010000000000000000000c00000000000400000000000003000000040c00003400000000000004014000004004c104001d00;
rom_uints[235] = 1024'hcc30500c400433000000c500000003c100011000003300c004000073000000c14c0000000000c4004c010c00cc4040330000c0c4004000000000c00c001030053430c000000300000000000c40c003000000000000c000c000c0000000700000cc000000c0000f00000000000030c000c0040000004004000c0300300c4c0000;
rom_uints[236] = 1024'h3c000c400000001000004000040000c4000c00000000010030040010000000c00400000c40000000000000040000000001000d0000000c003400100000000040000c00000c070400000404c00000004000000c0000000040040001030c000400730300c00c000c000000000000010d4c0400000c0440000004000003003;
rom_uints[237] = 1024'h30100010103114010c0010300000103000f343013030300000000010010003000d3003001cf30040300000000000000000101001300030310c00307c3000010000001007000030000100000001000300300000010000010c000303f1703100340000043000100010330100100c00101000001000000030104000000013001;
rom_uints[238] = 1024'hc00000300000000000100000000d000c0000033f0000000000c0000000000000000c0000000000000001000000040000000000300c0c0c011000000000000000000003000c00000000300000000400010003000000001000300010000030000004115c0000000c000c003000001000000000000030001400000001040004;
rom_uints[239] = 1024'h10000c000c00000400d500000c3014000c3c00c00410dc000004000c003c0c0c103c0000300000344c0030003040000c0004000c000000000c0004000c30000030001000001c0004043000000000c040000c00000c0c0004000000100000040000000400000c4c0c3c1000300000003c0000000c000c0c00040004000c000d30;
rom_uints[240] = 1024'h1000400000c000000030003000001000000000000000134000004070100c000070001000000c40000004000000404010000000c0000c340003100030c00000000000300030300000100000004000000000003000c0300030000000301000c0000000300000000000000000000000000000000000303000001000000004000000;
rom_uints[241] = 1024'h10100000010040c000040000000000000040403c00000000000000000c1000000c000044000040fc400000100000400000040c0400000000000030000000000000504000c0000000c00000c0000000d004000000000000000010000000000400c000000000001400000400c0004000400000440000000000040c30000c30;
rom_uints[242] = 1024'h330000403040000430130f3310c1000000110001001041310001400133010303033000c300300003d01c30335350f03010000040010d0011d0f34303c011010c030011c100001000c40004010003000104000c000100000000000f03c134170c00001000c3000c0101004001004330400010000343000c00100c30430000c030;
rom_uints[243] = 1024'h4003300000400030001000000010000030c0000330003000401000f00013c0000010400000c00300000010101330000003103000000000000000000000001010003013040003300000000000004010000001000000007030000000000000000113c000500000000040000000000000000000c03341000000307010;
rom_uints[244] = 1024'hc00000031d00000001d00100010000c000010301000453004000400000c703000000000300c3000130c00000c07040000c0003000000004000c000000000000000000300040000010300400300100000000300004010001000010070401000030031000300004300c00300000001c000030300000003000100c103c11140000;
rom_uints[245] = 1024'h7000000c04110040cc0c000c000000000c000000401400000c4001340c000000c0000400c000000040c00000050404000d0000001c000440000c00000000000c0c0000000000c0000000004000000000040000000cc0401000004014450003c000000c44c0040c000400c000400c01000c00000c0cc0301004c0040000030c;
rom_uints[246] = 1024'h7000400000c0c0400003030371c010000010c00000003001000301f000000050300010003000000003400c40000044000001000030c03330000c000014100030000000004c4300c00400c0003003c04100c003500c000003f000131000c11c03033000000010c3300c000007000001000000c3430000000041c0004000030000;
rom_uints[247] = 1024'h50000000c000c0040100f0041c0c017c03100010cc101000c400400c050c0c003c0000000004300d400c0000040404003c3000300000d0000c0104101c00000030331000340000cc40000c040c1040000000000030000300040005000004100cc000005010000cf00f0000000400300c0030c0400c00c400041030405033000;
rom_uints[248] = 1024'h10c0300c0300000030303030105f00010000000000000303500000000001000030100400301130000000011000300410001000000003001000003000010010300001001030000003000000000000000100100010000000000000000300000c00030103100300001010000000000300001000000400001000013000f00c003000;
rom_uints[249] = 1024'h4c00000030000000000c000340700c004130001000004000c0c700c44010000040000000c0c0000031000000000000014cf00004000000c0c000007000f143001cc000300010cc4000000f000040010003000040040000400c00000040340c004000100c400c00000000000000040000300000000000c040300c000000c00000;
rom_uints[250] = 1024'h300000c04004000501301000110000c0400000003000000000001000000c404000000000001c0000703030c01000130000000000001040000010100000400000003000000011400000303010000000000000000c300c000000003000000300301100000400043000004030000000000000700300300000000000c000c0;
rom_uints[251] = 1024'h33400100000000004000041f00300000300300010003003000000003000000003100014000100000010400000031004000301000000c00000000c0000000000000004000c30000400013c000c30000000003001000100040100000000000000000000000100000000000000000000003000040001100400000000000;
rom_uints[252] = 1024'hc04000000000000000000003000040000003c1c10000f100d00000030100040c0003004000030000c000c000010000000000000000000000031450000000030c400000004000000004c040000000030040000003000307303000000100c4c000400000000010c0000400003000c000000000010000050004c000001070;
rom_uints[253] = 1024'hc100c301c00101000000000c01030000000400c0c0c00701000000c0030000030f00050000030101c00100c30000000000004000004c00c0070000000007c000000003030000010003000c0000000000c10000011040000100000c0000c04000004000c030000300030301000000400000000000c00000000c0403c10c000300;
rom_uints[254] = 1024'h1010000000100000000c033000303000000400300010140000100000301000003030030000301f00300000000030f000303130100013000c000030010000000c1300000000003000000000014c00001000000000100030300000003103000000001000300000000000100c000000303000000000000000010000310000100000;
rom_uints[255] = 1024'h300001100000011c0500c50500000000000c0440000c310000000104300000000030000300000c330000000407f000000000c044300000c01300000004000330300003c00c010000300030400000000000000000001000000300000001000000000000341030001f00101000000000000c0000000000c05110000004003;
rom_uints[256] = 1024'h10011000303c000017303030c13001033130400100004f70c00300310c700c0c00c0cd00f00000000cc100000d00005000c000c0000000044040300040700000000000000354010070000300010110040000001000c0040010003003c031c0030000000000000004f00030040000004000000300d010c0c000000300c03403c3;
rom_uints[257] = 1024'h33000000403010030c0001010000030040c04000403034c0000031000c0003000400131007030003c0070c030430c31000000c0c03300001000000040c4c0300100140000330000c400c0000c0001c0003100d101010000003000000430000000000310013d3340100040000c03c003004c0000400c00000003f00d000000300;
rom_uints[258] = 1024'h3040c000004013000f03cc03055303f01010030000c300000000031103010c30001000000031c000ccc0c0000500cc0000000030004030040003c00000c3100030c03c00000300dc1000c10010c01000c3030403004d000400c04003134300003030003c0000c0130040000000000000043003d0041000c0000003c30000010;
rom_uints[259] = 1024'hc007f0400300030001000f000003014f004001c04033070003c3c003c04f034004430001034c43000344500000c340fc0000c044004100c0000000c0030000034040404103004031310000c0d34770000c400d03434000c040d00000c007450050c400030140070030c5004000000c030044400000033303c50040035011c000;
rom_uints[260] = 1024'h47001300c00157000303c4403dc143710000000c00d00c11ff0cc0c003000010710000000330340f400000041c0073013d10030044c00000c04450753000304000f1c00d00430f1c000740f00070400c00c041034003304004f13011030000000300c0434051d1000c354000ff00101cc0c00400c03077dcf00c0344004040;
rom_uints[261] = 1024'hd3c0c03c110000c040403000004000400000000001d00040c14c00404c00030330001300300f0001c0000400300c0010450c00c00030100003100130400030000000d30040000000000004000400100000000050000000700130000004c00000304000001000c0000000040000000000c000000000040000000003003100000;
rom_uints[262] = 1024'hcc013000003003c313c3044cd17300030030c000d000030100c0c30000000001c331014003000c0410c0040000f300104c03c00543cfc0c0000100c3c4c0100000c303001000050100000700000004030703c00000000000c040400074400dc01c0000c4f10003014300c0030300c1000000304003d0030300400310000cc;
rom_uints[263] = 1024'h3c10000000000004d43c00000cc0000000f000000003310001041004000030000307000000001030000030040001000c1040030003000000c000f01710000003000030040000000c00000d14144000000000010001430000300000000004300c07300c000c00010030010000000000000100f0004410040000300c0000140014;
rom_uints[264] = 1024'h341700000003301000001000300130040070003040cf000000033000c0173000f000030001000340c3d3130000c10104000c3000030003c00303000000030000000133000014040c3004100100305000100003300300300000103100400340000d000004043011c00373030100000000410000d000f00003004040c013001003;
rom_uints[265] = 1024'hc00c00c04c00000c3cc031f000140070000000f110f4c40c400003000c00c00000403010104070004005700c014000000401f33c0013000030004c40003000c04c0330f010004000dc004043007030404000c00074005c000050147040f103c450c7000001035c0403d4014c0040c000003000300c0044703c700400000c0000;
rom_uints[266] = 1024'h403f301014cd1ccc1304c0003740301010cf00000404000050c1c53000c00000c0010040100c04100c301040100010731000050003cc73000040001f0005c03c300c3031d005000f00300001c0000c0100103045001c000c0c14000001f004004000000330301044f011005030000000440311011014000c05040d000c03100;
rom_uints[267] = 1024'h30003f0c00000c0040100000504413000000010000001000000430310300001000f0c010001400030000000004100c0000000033400300051003040fc33000001300000000c3000c000000f0343000000000c0000000004103010103003c011000100310030c040003300004010030004d3004c300041431000100000000cc;
rom_uints[268] = 1024'h40030035140300031040cc030001340f341007000c0c0000007c00cf400f010030301000f0104000c000101000c0000400c000c0c0031003300000700010f0000404100030003050140007000c00100401000011c030000000c430cc043c000c3d0c340000103000d04000c0000c0c00000000103000cc3c000cc000f4fc0000;
rom_uints[269] = 1024'h301f00c000003103300c340003300c003000000c4000c40001440004044030003003000d00007400000c00100500300000c003d00000000c0004000c00000000c00130000100034c0d03000700010c0001400000040003c000c440000014000c0300000000c0c4c00004000300400000001c00cc1004000000000400c1300000;
rom_uints[270] = 1024'hc0001cc740c0005040c50c03c43005000344400010f3cd00cc000000040c0dcdc00340ccc441000341c041c10140400004c00cc3f3010d030040005704000c00c0c0030c00440004100000cd00c0300000000303c3000cc0040c0c40c3cc000c0cc104000f0c4f0c0f00000cc04c000ccc0c004010700101c30c0c01c44dc71;
rom_uints[271] = 1024'h3000000000c310301000000f0c0400000000050001417000300d3400c311003000f003000001033031300c0c3c001013007100c00cc103c00007300000400000010000000400000141000401003c50050c040000000001c10000d0003f0c0000f4cc0404000c0000c3010301000003100001c00f100004d0000000c330403001;
rom_uints[272] = 1024'h3000c1710c7400041d0c00400d050c00003100010d01001000140000000300300003303d00034c0400400101401010700d000c303c3400c004404100000030000004000313404441303000c40c3434003000001000000040041c0301000c0c00c00000004000000000040000000000c10c000300001d03030c0c00410700000;
rom_uints[273] = 1024'h1001000cd1001d00003010033003003031c3000f3000000c001310c0f00cc1000000340040c000003cd000001d000037110010050000000000000f400c0000400f3000cc400030f00c10000300300004000300003000c000300c11344100000000030c3c05c0300100000003c0000100400010004c0005000000000000c00;
rom_uints[274] = 1024'hc1c404000f004404040017003400700000000c00010000000cc3000000c00c0000c00004010001c00c010000404000000300c00000000044c403ff00c410040003000314400000000c0d0cf0400000030004010000000400000100100003000400004f0000070c0000c00040d00cc443030000040341c4000310d3c1000;
rom_uints[275] = 1024'hc00140f000f0000050c0c0f0300000000300000030c0c043c033c0400000040170c0c401700403c403cf0404000d504004040000c1f013c00310c03000003014c3f310003044400c101000c043f340c3c0000053c00000c044003000c5030000000c300400003004c1c0000000fc00000000040c3000004003003300f040000;
rom_uints[276] = 1024'h7c0350c0030140000f0c300000100c000000400000330000fc013100c000c000000003400c300000d000001030011000d030000003000070000000000010004000000034001000104000400500000000c00000000000100000c001044100c000c00000103003000c00003000c0000004c003304000000c40c00001c0010000;
rom_uints[277] = 1024'h40f3000040d043000000cc001c03000043334400c00304d1007c0c00c0d103c000c000001403c3f0d00000000040c04000d000001030c00cc030c100c030d00003c30c4f100000c100c030c04000c0000f40000f40001c100c41c004704000000030d00000c034c00000c10c0000044043010303c100f0040000004004c;
rom_uints[278] = 1024'hc0c030004300c03000000110cc0c003000400030130000c3530310300301100570001010040030007c00304300000043010404c03000000001003070040034003000030101401f0104004300700004040070040004030004034c0043c0cc053000003d00030000004100003c0c3010000330000001040c00003000430003;
rom_uints[279] = 1024'h1400030c100000113c00000003300000070010330101f00050301030001001003401000000c00003003010033341410003000340130d00000000033400000034104c000303000000d0034430300500130010014000000000535c030100700c3030330004000050000034000003c0000c0000030000003001300c00030031000;
rom_uints[280] = 1024'h1000300400003000310dcc01140005000c0000003c00000040000d0000000404040030000cf0c0000c04c100003c001000000000101040003400140000000030d04000033c01140000004001000010340000000c0000003003003c0411000004103400440c00000c000000013000000000300cf0000010c400c00d010010343;
rom_uints[281] = 1024'hd0c0003c0030c0000000000000000100c000003c33000000004300000c00c0100030c0101c000033c001000000300140c300000d3000000300000001c0d000c4f000d0004000c000c0000040c1000001030430000c0000004703000010300304030c0000000000c0340000c00d000000330300010003000000000010400000;
rom_uints[282] = 1024'h4033c43c0330000114100c01c00c4000040015c70c300c03003c00cc30300c00000040000040007c1000000000030004003d4030c04010044004c03030f0104c0101034010751401000000c00000000000003c000000130f0c300c000000000c0400315030c0000000010004101000cc4c0403030d0010000cc040143d103;
rom_uints[283] = 1024'h40000070500104440f10d0400334300030c000c0100040300300300c0000300c40040030401c00001030c000001400003d50001003c100f40c000c01d00000c1c000c0c430c000f33040000c00c1f00000c0013000000000010010c44110031333300c03f0304030030000c030d0000040005000000000c00000100040003c1;
rom_uints[284] = 1024'hc000c0013c0c300001101cc0104c4310004000404cccf00030f001fc0cc340c700300000c300c000034001f0103005400c01010c4004400000411400504101c00040000304511c4050030000000103000000000d000000300400f04003c000c034c000001003c03140c00c00c010404130f0f303c00100404400c000400503c;
rom_uints[285] = 1024'h44000000003015300401100100000c400000034070f00c001300000c331000000010000c40000000300030004000440310000000010070d000401c0050000c0000000001000000000040070000304f040004001000300010000410070430000000c0043070c00000c03004010000c0300005c435400004040d03400000100000;
rom_uints[286] = 1024'h30000000cdc001401c0040000000d0034000000000005010f00030413c01c300433000000040c3000004c30004305000000540cf1000c0c00c0031000d5d4100c0001c40105010004000cc3030300000d0c00010c130003000cc41007041c400c0330110001000000f00000000c0000c04c30c0c004000330400c0003041c400;
rom_uints[287] = 1024'h341000000c10040004700003c0310030001033100c000303030001ddc00000f4030010000000001007c00004c03c10400130000000fd0000100034400c004010c10d050000003301050000005011000c0031000001030000030000300013c00703133c003110000103000030300c00000c3100400c00074003000044cc07c0d;
rom_uints[288] = 1024'hc03c00c001030030000000300310010000c00000433cf730103000c0010000003000000000000033001340c0504030f000104000d05100c0000003030530000001c00030f0000000010000400300c004c000004000000010000003403403000000030300003003000000000000100000000c300303c0030f1003030010401000;
rom_uints[289] = 1024'h500c00000f0300100100c000000d3030134d30100101450000cc404010000100cc101103c0c03400313314c00303010000000c43004004014003f001cc00d00044030101c400000000100010100054303304430040400000404000301001c3cc0030400c00047f00330003000701010004c044f0c00100010000040303010711;
rom_uints[290] = 1024'h130040001300c3004050014001f00000f00113030c1c000003300030000010104100c0000103003340c3000000000d003030034003000003011440010101c1001030330300000301000000300000d000041311003010c000013033700040c00003c14100100000000300c1000341000033000c0043303313310003003030111;
rom_uints[291] = 1024'hc40f01000010000334010504350000004c0c0c000c0104000c001000003c0005c00f0004001403303fc0c0107013000010040000f100030313043c3030d00000303000300704c00dc00033103010000033000004100001003010470d101000041334000c00c400300c0330000000001010030f0000440000441433304400dc;
rom_uints[292] = 1024'h300000310c00c4043c3c000c3c0000000000030c001510011300141130100c000054000c00100c0000000000530000000d000c00000100140c0003310d3000c0000d000404003dd1001130040000000c0c0c040c000003000100030100404c3f40c10c00000400010000f00030010004405033c0040c0c004c4003c0040000;
rom_uints[293] = 1024'h300010000000300003000c10030410000030000c0014c0000000003f0500000000c4000030110000103000d00100070001100c00704710000013003000041040004004400cc040030c0100c501000030004300010010101040000014010000000000030304c0000100004000003033100001c130c00000043100c001300033;
rom_uints[294] = 1024'hc000100304003000300c001300400000444044dc00000300100c00401300c0001010010040030000004dd4000c003000400400003f00040030c04040004173000010c00c00cc0c7044001000cc053100000030403403000000043070040fcc0010cc00040c0300000c030c0300003034c4c400c0c00c00000003000d10000000;
rom_uints[295] = 1024'h150004330411c15140010030040401000003030c1300c303100300000000040001010000c100c0300000310430000300000033000030300000410000000000010070004101000000030004103000000c300000010400103c0c4004000c00c030304010004000030c0000000003030007000000001c00000000c00004;
rom_uints[296] = 1024'h13000030003000000004300c00301c00004004000300d03000010000c0010003300310c0000133014000c00430304c14300000030030100011113030040000000004573c34000430130000300cc01000c0000010000040300d70300040000000304c0d0110000040000000000030000003000c0000040070001000030000010;
rom_uints[297] = 1024'hc0cc004040fc540c050401c40c440301000034c040c0c00110000003f0000000040f00000440010c00401c0000030400040f00cc000c0010340c0004c303000000000cc000c010003400c113000044000000c0500c50030104000303340f30001030cc00301f04040043c00c00c0c0c000c0c00c000400000000430000010540;
rom_uints[298] = 1024'h1c000cf00301000101300100004100004c0000300034000000001040040000100040000000000001c000c000100040000000000c000003010100300000c400000040030105400c3100000000310010000004c03000000000003050001c000400000001000000000004c000007000000c000010041000003000c0100040000;
rom_uints[299] = 1024'h3030001c00010000301c100000371000350f03c14c0c3000000c010410f00030030c004010c043fc70030000303c03000007d000c000000c03000c1300007030010000d1003040030031030000030031fc04701000000333c0130003100310f000c010303000700433410300d0030103110000003000000000133000d03000;
rom_uints[300] = 1024'h1040c40c10400400c303000000c00000101010000f0030004c000000c00c0004f130000400304000134040340530d0100000c0400000c0004c04040d4c1000004070000040001000d00001c0004340404000010c40c00040414c04440034000530c000031005c00f40c00104f00000c0000c3c04fc004100000401000000700;
rom_uints[301] = 1024'h4c301cc001d050040c000010c400f01000c0400c0300040c7030000c003c000c0010100c0c3040341040701030c4040d1c0140100004300400c00014001030000c0444041c140313451000100000300430403100c0c00001c0000000540030000000030c140000004010000004100c0d4070000030003300701004cc043c0;
rom_uints[302] = 1024'h1000c0030433c0000c0ccf0c0004c40d000301c0033c300014c00f0f1c0c0c0c403cf04404c000c000000000003330cc000310000047000000010404300003000f00000f0c005040050000043ccf0d000c007000000c0004004030000000c00404c05300500004000005000000070c0004f000cc000c000c0cc1000000c0010c;
rom_uints[303] = 1024'h400000000000000047013100004c00000003040010400c13c0003c0f0f0400000304140000003c053100000340000003003c00030000001030030300c000003030004c7071000000000000f0000f0000000c0300000400000043030c001004030000010d0c000004000dc03000000000004f0300110c000000000030100c;
rom_uints[304] = 1024'h40c0030000113401c0000030000000c04000c0000c300f400c3000c3001070000c00000c440000c500c00440457005c30303000030cc00000030c0c30cc010000340700404000010000070c00000000000430c00000000cc003011f3cf000000000405030000400004000000000000000c0000300c04000000400470d140;
rom_uints[305] = 1024'h40000000040d0f00c0c040000410cc003003c0c3300000000300000030004c4040c000400cc440c00cc043010003c040010044c00010c000d00c404000000040c0001400c00000004004440101cd000000000004010c0000470700000cc00047cc11cccc31504004000040070000000004070c400004000dc0000000000c30;
rom_uints[306] = 1024'h10470010d0001351f010c0000003100d71000000010300c040103003003300430010000c47040000331000cc01400000c0700030c34c70000110c30000000410c0000040000100003013c400041000001c00000000001010c0000100040003c0013f0100000030300003000d0000050400044000003001030000003005030;
rom_uints[307] = 1024'hf0000130000001004150007140cd00003030410007310000f4f0c001000014004003f0400011003010f0004301cc010300f0c10000cc150001c0cc013000100333f1000501f00001030000000d100300100d000000c0d0c000c0c000000004100c0001d330c000030014030000000000c0010070c10117003030c04003100;
rom_uints[308] = 1024'h7400001011000040410070010000430c000c55040000403300000001003103c433c0400f1000f3000f33dc000c00400fcc0c00c00140f0c400c30000c151c13000000c000030000c5100000c30c10c000013c03f00c0000300040140030d0401c3305c004f0c00f001433f00cf1000000000037000f0c0c30000003300450f01;
rom_uints[309] = 1024'h700000c40000000010c40c000000050000000030101c00c000104400010c34c0004c4030040030040c0000003000300400c00300100010004fc0007500c40c00d0003000400003004010701040430030c00000040003c000d0001000444000033c00000c0c01000300000000004000300000dc003017ccd000340c30150c05;
rom_uints[310] = 1024'hcc03cc40d00c0c001043040004cc4f00010c00030303000004040400003100f07c0c0c01530400301c3c300c0400000003000400c0000000400c307c0001000c0c00d000040c030f003000000c0c000c001000140c0004003c14440c1000c400040c00000c300117c1000c30030c0030c4c470000414000014140500010000;
rom_uints[311] = 1024'h10000d0c070d000c030730c0000304700d530cc0015050fc0c30c0100430c0c301c01000005030103130000034c34450010c000dc00000000003003c004c1000c30c10000710000350000cc1010000c1c3003000000000c01cf0300010100343c00000030d000c00304101c00000c30000405030100304301c1000040007000;
rom_uints[312] = 1024'h300004c3300001c0f00000c0dc00100000c00000000c03100000340000300000c0005400100cd00004f35000c0441044040cc00000c000c00000c0f400100cc0c0dc1000c0000c000000c040c4000030304030003100000001100045d0001c0000cc01100000041000703c000030100010000c3030001700304c0c343c010000;
rom_uints[313] = 1024'h107000c000100100c0c0c030001004c40cc000104030000d700000000000c03400000004010000d3001004d000c0c0041c0c4000000c7cc0001034c000c0c10000c0100c0000d000000000c0001000c000000040000000c1000c000010c00000003000c0c004000304000000040000cc00400040c0300000c00004000034c;
rom_uints[314] = 1024'hc000c0030fc00c0400c1cdc1100c0400400104000ccd03cc00c0000003000c000d0c40000000c0040101c0c30c0c00040001c000000003c000000c014045000040c000003040004104004000330010030000001000000003000c0000100000c0400c00030100035000000000000c440000c3030c330f000c00c0000cc1000d01;
rom_uints[315] = 1024'h300000400c50700031303030c1c0030000000000300003000300033030003400040000d0400000c3d00000001c031401003040001000c001d0070034300001700070730000c300000410000040301000c000434010000000d00c0000041000040c4000c500100041d0000300300013d0400000430000010031400000001101;
rom_uints[316] = 1024'h30c0100037000c111030300000000000000c00003000c03c0c30f0300030f0041c30c1003001301504001533000c10103040ccc0000c000000031400000010c00040004070010040c000000400c0001000040000040000040000c03c0100340001005000f4c0500004c500100c00000000d0003c00100c400000c4001000;
rom_uints[317] = 1024'h10500c0c0d3310400001000000440c00100c0001300440000003d3000000000c030c0000000130c3047c0c3000300030000c00c00004000434c0000c003c000040040030001f0030001000cc0c00000c0003001000c0010d0000c01ccf04040c000c0004030c04144300cc000c0c0c003100001c04050c040000001c100430;
rom_uints[318] = 1024'hc04340c0c0c005014003c0c00c00403001400303cdf5010000000045000105c3c04c40001000000300000400000000000300040301c030010003030041330004010131010f5030000400c30000000003c0c10040c00c0300000003c1c03000030103c3003100000005c00340c3c1004050010044000000c00100c0c30310004;
rom_uints[319] = 1024'hc0400030040004344c7000c00c0440000014014c000000000000030000c00300c04004c000c0c7703034f00034f0c0004c0000100040f0003100f0004100c0003030c00000300c01c04440030030300000000440100cc000003000c040c040000041c0c10004cccc005c4000c0000040400010c4000000400c0700000c10700;
rom_uints[320] = 1024'h5c010d3030fc0550470f37300f3c4047117c43010d5c1c70f033143040704c0c373111403010430c0cfd133d3d375450c10df0c003701003431c30300071f01c11c040d13353500d40113330f41151350030cc01f00d0300003333c31df10103300300005f433400ccf01c3040f00100f0c3df1000401c33001c0c04f1340c03;
rom_uints[321] = 1024'h3303c0344000c4303d3c7d74f340531c1c0c50f0cc0c33c000c13cc33000d33f34c013033700c400cc034f30c500c0100c0c000100f0001ccc1033f10f5d100c13017d5cc0c0007c73330700f0111f00335c4d0f4400d000070000fc73c10001f4c071dc5fd734000c00c040c3cd0030040104c100c00dc1000cc0d0f0c03330;
rom_uints[322] = 1024'h700c3c43444401d30f100cc143100cd11cff1c30c0d34c30c03c00007010fdc03134df4ff154f104cccdc07070331010001c7543c04001c0c00100ccd0d000c5c001cc13f4c53c1f1c05cdfc7dd01031c400413000003005f5c374fc0f00070d307fc0cc0000f030537c11c040fc530004c404cdc4314c0c30c0003cc00c5fd;
rom_uints[323] = 1024'h303430770c37d304013f1c03001c70c300454cc31317340000ccd0c000133030c047077103d00f0403c30737c3030d010c03c0040074c000d13d43110010c400700005310c01030043073400c0c703c103000f11004700004000131030074400411100350d45c0c0337003403013c003c001300404100c1000d000c10cdc0013;
rom_uints[324] = 1024'h7d03305370040c07330437d00071007431000030400150034c33f3d300370040103133000000c0070c41030710dc044001c1100343400100303c045035f0c0300300f1c000c030cd00030340c3c0031100f1003104703330007101005dc70000001441377000500dc10f30400c000c001df0000503c30d340cf000f010c000f0;
rom_uints[325] = 1024'h314c000f0df3c10dd4ccd3cf10c47050c0171d341155c00300031410031f040d037401310f0103001007010f03001771041dc330100f45000471130301010f007d0000040f3030001d3c3143031c01000c050005c00110333013c300300f000073c7cc0035010f0434034003300c0333cf3504714c501417cc04cc770f1c44d0;
rom_uints[326] = 1024'hcc0f014071d47c030013d0441000430333f173030301f040c0030c000303300d10003c0140030410c7100cc450030307c0031fc03140c303f000040033c4c300c003c0000010130d7c1000004030310407c3030cc07013f000d133003d7010c110114f03d3cd7030017711000700f33f33d0c7c14d031713370037005c40037;
rom_uints[327] = 1024'hc004c3054cf51c04103013010c0f0c00030f00c043ffc5000d071703074c040001431000010c134f404c074c0c0c100c0043c0040005000f103c0c1340034f0341d303c7000c0c0705004143034003413000301f01430c004d5d0f0cd1007cc31330100c000c0d0c330003040443100c31c4f1000450c313013300000c00c014;
rom_uints[328] = 1024'h370400130003701400d31341c00d00070c3c33000fd37f010007f010310030031c0c73c00104034033100000003034340c3051030041330033f40c0000330fc3c0c0033030140403350003c1030377401330c33c0040010307cc4dd3400f710c1d4cccf3c7304d001000030100c00130000340303300dc00004071d01fc30003;
rom_uints[329] = 1024'hc0c0ff030f43030dfdc50d130454107104331cf10034030c370d0c0cd3003441d0013317030001c43004701c011f300405040c7c0f1c75303c005f00303c0ccd3003333c1c0d103010014c000f300110404c373073340c04534047000000c4c710051c0c0107130030173154303d03003f3704337c0144310c450430010c04f0;
rom_uints[330] = 1024'h3750f33c014d1100013f0d0c433733fc040f340300070411000d130c3c0f013c3d00d4003d40110c3503310c3d0d10030434fc500cfcc7c31400c00cf70c0c04c40c34105d070007f04301031c3007011c0143074040070c05c10130344c01000033000007000d00530d00f50f0030000c044001cd01571ccc500c13fccc3011;
rom_uints[331] = 1024'h7d0010000c00331c5410513431f010000000cc00c1041314f3140c30c04313c513f330ccc0c1c43410c3044000040333c0300071f00130c0003c1013c0010004f03c3101447540c0df0100001401f37077fc00030030c040c3f00045cf40114503450000c0c0430c3c0f0003100500f003754143040030500f000100000300c3;
rom_uints[332] = 1024'h433303f0d000300703007c30d11d304341115700301f3430034c4cf0040040c570051700f100000450cc1007f03034f351f03013c330404f033300704000f1400714501034c0c01040d0373033d050f0c300c011c0c4003007353c3015f3c00c3d0c340013cc7411d001033000311000fd00105c333c1d7c3400f013f4304040;
rom_uints[333] = 1024'hc1407dc4003301345cd30c1cc03004c00c14c40004d1004cf047400c040300ccf0ff01d1f4434030dcc001000c03340000000d0c0f3000c40400c00c0400000dcc0003404f0437040d0c70005110cc0013000000430700fcc3c0473dc135003137030014cf1c003c0dc401f00410003170c00f01037004700040030cc001c74;
rom_uints[334] = 1024'h1000c40c343df341050c73cc4c03c741334044c3440f35d3cfc014d43c7300dd13c3c1cccc40dc0034df05ccccd4747407400cfd330004d3740000c44c750fdc010f40313310410c71110001c1310000004300077c3c47f004533307c03cd003c0c0c040113004f307f31070c3c43000c300c0f400c7cf000c300cc41f44dc40;
rom_uints[335] = 1024'h45c3433040f1400cd73003003030051cf44d517043407140f5f04433d053044cd0f07d010d5f070c4070033370f411d0c750c3f0c03500311c1030c30040c040c0000340130300405d03300010304c4143c30044c30000010cc4c5c3713cd0c5f1c40000404040f033c1fc31c00340c341d4c110d0f4c4d031cc01ccf04f3053;
rom_uints[336] = 1024'h3730017c1034c3071c4c51c03c100fd01330c07c0030c0010f403fc10c000c345010f43170044c0f0d3300300c10100011f000303000c00403fc005410c03c4031310037030c00f103043000403dc4003010010130ccd040111c1fd5340c0c040f5103f300f5110cfc4041103c11000030100cc5331104543f0c30004f00074;
rom_uints[337] = 1024'hc000405003350f01c0c5c701304303f003f31fc10cf110004d30c445100730f3107c400f4000c005357cc55000111004037c1035c14cc0010100c0000c0004c00c13c3040fc130c31f04f1754443001cc00f014c00400000cc4f44c01f05440440040003f3cc11037070300d00c001010004010004cc030750040400400003c0;
rom_uints[338] = 1024'h3ccc001f7c0cd130007c535c4c4cc350300130334d31cc03cc00f400f04d300cc300cd1cc340000d40dff4d310c77745731d4c3ccc0000f430305f007c30cc00010d3c3000735cfc3c3c40f4c51d01003c30003011114300007004370dc11040f3034440403d103401cc00f00047000c0370000000500004c07cc0105c3fc334;
rom_uints[339] = 1024'hf741d40f3f7c0000000fc0df33ccc0043130c13033700c073c170073c07c4507d30c700c0341f440343c05530313d404f04fc34d3c0f30300504c303cdf0c3303dfc304117010c30c0110f034041310c7c3040047c0003c3ccff4307cc4f0000d4c13f00f540d3004cc030cf00330000103d0145400031f403300f030f47c014;
rom_uints[340] = 1024'h40cf530c53f543345f1c0300dc030c0434133031f4c000000005c107f1f70cd7703100001c0140001c33500cc0c403c00003434000f0c035cc1f04f0050ff17f00340304315334134f530035713d0030f000f10c0dc00000c00004c341001050d330f3cf00d0c51c173c7f03713033d000003043041c14f10c0f313d000c05;
rom_uints[341] = 1024'h30345c104d154010fcf0300cf3310030043137f4100c400c5f4400c4cd0d3c70f3303c4c050110cf3f0c1f00040034f0c01c4d0f0134c31030fc5000c01cf0fd14c13441c030f0400c70cf7710f51000c407f001c000000df050d4310313040f00010cf13c50d0345fc00f0cc0c010501550105010f0404fd41f00cc300044;
rom_uints[342] = 1024'hc30c3ccd3144fccc0f115140114c1010031130c7370000003001f73130403031f3033cf03001403307d0c0c7d53c0f3010311c400c3300c003c0110434c4c033c013c041f3101031f000400473c3d1341400440c43005010dd3570fcd03030411c4cf30310c1f0035033d0001301f0303330430007035c10f05d4310343030f;
rom_uints[343] = 1024'h1100007ff1f10141140030341c3f1c0003c0054330c30303c0cfdd03003c00403340d000304c043300d3c03133d414510c3f03f04c7cd303c0100034401030030500d003301000304c03354303c7500130013c13003300000534fcc050f303f303d33700100475d30c3f1c7010337030fcc4f000051703c073c33cd040301400;
rom_uints[344] = 1024'hd1037003035c30c1741014043c3403d00000040000140d0f71313c3f000f37f4f0003fc130c077c33017c0301c3d30100cc0034c0010007134d45003000007005c00333c35301073d0c0403c03031004004030003ccc0310007031f710333000343c0c141cc0000040000030001ccc00107370050030051004c001143df3303;
rom_uints[345] = 1024'h3001c0c1c1c3cd01c01010000310f011303000000030300003504301035c03c30000f0f0d303400740c00cd00043303040cf03c00d0030303330c1131100d103c1f340c310400003c000100170c1f100c100033000c000d00d43c340f0d0f0074043010137000073c0c73011004101d0034303710040034013001371c1513300;
rom_uints[346] = 1024'h1c4433104000035437504530d11c00c10cc040005013f3700040300003c7c3d1f4010f03f7c0011157d14054013c313fd1500014430000c003130000544303d045dd00c333d101504c50001033034c33000000c310000000f1003f50c137c100c5c140301103f0c0c0f3010400414300000fc3f347f0100000400cc0d143d033;
rom_uints[347] = 1024'h740130c03531004500010d04cc307cc10f5c344f017c400000cdcc1c300f4f0d770040f30000cfcd011f0045d0c0040c7fcd050100710f0070c33070000c103cccc30c0c401fc30f7500cd30cc0c03d000cf010000300f400003311173c10d3dc003c1c03f031407c031cf0543cd343044cd050c015ff0f0f0cc05df1c00031d;
rom_uints[348] = 1024'hd013fc30001cc3403051010c4103c1010310303c0404cc3c033d0cc00f0130f77157d3330dc04c0074450430410c300700c30113330107330004017403001303400501c03c0101c1f10014333dc713300010103313d7400051700c44c0d31f0c4c5c33c745107033100c4033004003c3c013df003300107103d0df4147314300;
rom_uints[349] = 1024'h30401450f3c543000cf0c003cdccd0313350c30004031400c305c003013043c7013040c0c0c400075403035440fdccf1f03413300cd0c03040f0c0c1f0ccf5c430003f104334f01013440c0444400010f1300101c030c0c501cd0c401040c103c0c0d33fc0304000cc100003007c0cc01d0c4043c47000001030c040404c0c0;
rom_uints[350] = 1024'h30003001f0043d5c7d31f40c01d331311c4103f43447d3c0004c007c7d130047c05f000473dff410c31c05c4004c3c1c7500fc003110001c7c04033d1d003cfc03110c001c304d41310031033070f0fc0d011ff03411c01fcd30314731000cd3c30d3c5010f01070c070c1003d0cc054fcc000301034135000c003f05d000d;
rom_uints[351] = 1024'h7001043fdc3cc371044f40414fc01003000c03010001c30313f001040000c0730401cd0cc00cc3410d7f044173c0c40400d0cc4cd0cf1400c140c304ddc100434c1f0000c0443c4cc35d0001c70d00c00c03001100c000c30013c3f55f350cc301744010430004c00df3400130000000c4030005f001007400300f344cc44000;
rom_uints[352] = 1024'h43030c04ccc113c44c030c0c04034f000303c405001f430003c70300cc000f03341df0030c0030c70d0000c007c7001401d003cd10c04003410c373414d00d0ccc0003033c0004c30c0c34100111003f00000445c30050310700c7c0410c30430f30000f4340004d0c34c00305c1031030c30000c40007410001000d070c700;
rom_uints[353] = 1024'h410110300c310111dfc00033733730304cc3c000cf57500300c401f00033d17c11014733010c0003d370d0313300d00001003000030070040030f45000100f0140700c101c3003c3100105c10101403c300c010c0144f0f0043000f74c003300ccc00c337100c403f351000170d0330000d330d111c33010013d0d007ccf31d;
rom_uints[354] = 1024'h3c340070c0301c34000000100010300c00d01c0530d030300d741c00005fc00077111c500400333c303c0030304c000c103c303400041c0014cc003010141000041c10c43f3000001c04340530c01c00070c301c130ccd3030103c340044003035003400ccdc001c00310c00343000000c0c00cc7404003003dc0f303007010c;
rom_uints[355] = 1024'h30000c03400103300f404c500c4cd4700000000110f00c0c74c330c00070c0001045fc0c1401cc300df03001330003f0401003034314003003304413434d103000c0043c31334c001040037101f10c00000000400000400c0040043c11d004004030540c31cc0c0430003f40f011d00004040530c1044430103c153d144d3d0;
rom_uints[356] = 1024'hc0c0f0043d1cc4c4047d4d101f7dc7510cccf5c33dd0c7134c4c04041370104fc7c004000c00507c074f000010040400004d001c00100003371000c0f1fd4c40c00cf00403471cfcc100103d04c430000c0000031c40301cc7cc4c00c04d4c4cc340c0c100041703dc4fc1c1c031cd0c034043c3d0141c0f037f4cd0d0054d01;
rom_uints[357] = 1024'h40cc00013004000cf571104044300010003003705034c4f040fc0000c040c0145d00c0001c30110573110c0011cc01f00441313004305000c000500c30744404100070f0300004400300d03ccd340000141000300c014c501040c040040d04000c04403340f4dc000430013c0000d000cc040000f0c10400cc34000c41005cf0;
rom_uints[358] = 1024'hc00c700cd003d1400003170070d03043c400c00c0f0cfc00114f74000c3470704c100d300c330043000c13400000300cd01533441cf001113430f01014c4003c5500043c54710314fc7c15400054000503d430dc041cf10305d5c3d53c033303003c11303c030dcc003f0110301000303d3000107030cc00c1300311c1117004;
rom_uints[359] = 1024'h33c1c1c71003004c1155d000d40d0007441510cc37004cd00030301334403140f00305303030000cfc040000c340c403c4000004d00100533d01000450003100010430047d0300d50000c3303307d00010000004c003c07000d05c0010c0000fc013047174104fc0c074d03003d00000030c00004303400c000070304100f4;
rom_uints[360] = 1024'h1303403d033c03031434330400771030000c10313140d330100f00330f300407743c100431073430043014003f034c140100300d0030103111d4703101013014c003035f3713310c1310300fc131d00130c0405301034f30047c00331d310007034031c0100f00500c40334001300330f000000cf01414f0f010330170000c0;
rom_uints[361] = 1024'h1c0f040433053f0f5fcf1c70000037000d034f003c040400cf43000f30c0430f41f5f303f43c50c005101304003c403000f31ff4333431c470100f0003753050d701d30f0c4d0c134300c0c0f4050410100d05703131301000103c375030000cdc03103f54c41001343314c34d0003330cc004000040c300dc0530144f00540;
rom_uints[362] = 1024'hf001c50f331333c0c4d3170c1c03001700043040305400003010040d0003043c344c310c030cc4000013c04c13310531407010007ccf044535051c0470007f300cc30400c7111f3cfc110c3d030c01c0030000400003400c100003000f001c005d00c0001504030050010c0c00030cc00f31010400714114c03000140f34f3f7;
rom_uints[363] = 1024'h7f040017130313c50041d100310c07d140330c0010730cf14c4500010c1d3130c7004f4f50d0c143c537040014cffc7c4d53030403140030304f05c000100070c13c0000d00000031f000000c3307303c00c040053430c00cddd1fc4031743433170cd103140033c0473330f34cc0f000040400010313c01307353f0c0d53110;
rom_uints[364] = 1024'h31443c030005c1040c370700c70c0d0003317dccd5f530c414330c301c0300c043530d4c033003000004144717033c4111d00f44000c3cdc3c313f030cf100001310f73d00000cf13d005c1fc71401c40004050c450000001713d0d4710300005340170d31335f00000304100cd50130003340d10313043303c40004c73f0401;
rom_uints[365] = 1024'h44c0310d5430700300100003df0010100cf0000333300dcc44004000003030310000f03007f05330000475153c0044d003c040001c000c0c0cd400000100f100c000071300d0cff7010734047c01c10dc150105010d10df1c04040000c00100f00c103000434c01c0010c030003000000c0040300f50070f504404f00410c;
rom_uints[366] = 1024'hc10c3d5714f413000cccffccc007543c1ccc1400c3cd0500340001dc00cc400c0300c04104f04c3cc30c00000cc400d0000f003c1057010cc00030037030130d00000cdc03c0c303440500041fdc0c47cc03ccd103cc0c4f004703c34400f100070044100dd0c710fc040c474c070c0c44fdc1cc07cccc4c53cd01cc03147d10;
rom_uints[367] = 1024'hf0c04c00c304f3031cc30314f10071c3003000fcd7c0134100170c0c00cf7fd750f3f3c0041001000f05c00040130fcc01c35333037033313cc0054cccfc0405303000f04f0d0505c3d503007333c013f47c103f07c0f140300c003c0703d144410303c3fd3c000cc143f1c00104c1c05400503f0f0c0500443c073cc30c043f;
rom_uints[368] = 1024'h1c00430f3300301000ccf00c1033d501104303030000cc401f7043301ccc300001001c00f00c753034d530300070004c003f14c00c7330d00001043013d300f0d000c30c5fc5c5c01010034040001000d000305033c000f3d03333371d30cf331035333005030000c0c3111c10330c00003f030403f5000403f07c1531330043;
rom_uints[369] = 1024'h3f400f0d04c411733ffcf0031133330c470033000411313dc473001350c140004f4100030034005500dd7c01d1cc731307511017304003c0c00fcc4d73303c0dd4c0004443c000003f4700101d11dd05cc040304c4150730c1374403740d0d33434fc003cf0c05000453dd44000400300007370c004407404c030fd1c00cc073;
rom_uints[370] = 1024'h7f00301c1c0d4310341c351d0ccd103000171003110307f000c534300f7000f0f0305437c40071c1d14f00cd7cf10037000c303d430c07f0043f3dc03c5c4c00700131d4f4403010d3c071c3f0005f11407dc1737ccff0c17030c01113c1c1c1f4c11334471700c00dc51c0c03111fccd730c154c00df0f0c4c1c1404c004134;
rom_uints[371] = 1024'hccdcc070c331030cc0c511341414001130334304f0cc4f33037043cc035c037044110f40440101c014c10f00014303df14cf00cf130cdcc103d04007031f00c5ccc00cff3040130f430c0c433cccc100301003d3c3c3100000553307410cfd004141c41fc1cf4444cc73c54030c533c3773f3f037f010501703330000543010f;
rom_uints[372] = 1024'hc0004c0cdd00c00440707dc0ffd153f10c7f100000fc3333c0400000d4f1033f03f44cd010fd37c0003fd0c0004300c000010cf0c054c3f003c003d0c101c0f0c403307f3530005c5cccc5fd43c00c00c00400f3003c0030c3c44c403fccc340077315c0433014f0401f30010c0000f103f04770c4003f300303014300443305;
rom_uints[373] = 1024'h334000c1c5c4cc4000d414f300c040053f4f0030f10300001005004000f1c034043f0c10c1004374004f00440050c1300f10310300f54f13033354c03040c4334013403fd00c7410013014300000335000c3c30cf033c3c000c3c0d1330174c010f043334340c10c031103f00003000431000001010007c030430400000013c0;
rom_uints[374] = 1024'h3c03ffd50101dfc070300431310f05300d40c00400cc0010c05041000103140f00cc003fc573000700c30000004c0400053031d110c3c00340303f003034110fc3c001001c30f030c07c070101143cc01f00004011c0710cd3f11030c0040033c540f0f33110c0014cd070c40500c3331c4171100011305005455010c040000;
rom_uints[375] = 1024'h401035dc344c1400c13c700c3c30fc070cc033d44014d0d0c0c000100040004cfd50d403cc04700d0413041cd041017031d4f00cf3f344040044f00c00c03c4453ccc03cc07530043300c0ccd000544c5c0004144015000000030d0000c000710c357c0037101cc0c0fd101c000010103c3100451cc17000c0c0c1004c0c4cc4;
rom_uints[376] = 1024'h400333300500040c013100000c033000d030c0c00003c301001130007000f010001000033dc34000c30500c30100400334c0140330501f114030c040000030040000101000c0003040740c000400040440000001001c0335000101c304000d1fd03c1100d34003c00cc00303cd000003010104000113d0330d40c0c3310001;
rom_uints[377] = 1024'h334017000dcc010314300f0c0c403f034c4c0f404035c3d034d41d0503011c4c0040cd43c07cd3010d34030c010cc34c40713f0000c740040c00030c700cc04d00000ccd1007000d0f03c075c1054d0001101d01000170c00f43c0cc0fc5c0cc470000010f0000440cc40073300000430c01c70d005c300c0f01cd00000c0f03;
rom_uints[378] = 1024'h170400c00f73c0f505cd0d405f0c57114c0104011d5c001f007c0100001d0c4c00c04c03f001f3401150c0740cf3c0474f013f70c00014000013cc31c105c040c50c054c3003c3cd01003c00400043c4cd0004c0005c000fdccc4cf00700730fc3000753103cc313440300c05c03400043404300f00c5301304c430000fd4c0d;
rom_uints[379] = 1024'h3410f13300143003cf1351000f4d0010030c3f0f0f0d03c03f00d3430340f11c0044f0014400dc10cd1c070c11c0014c0333040c003000c4cd13433073000c07013700070000030c70440c300000c030001f033703cc0000073000017c000f0c40c400101c0131300d30c1310300733d3404c03400171010331c00d10040105;
rom_uints[380] = 1024'h30154330000c30c44cddd5c310c0310100044040d3c07000300c70303c03303cfc043c403d401010c3d5c000d13c007f34d0f00c5c31000c704cc00007000014c500301c331001d5001000004c0100fc300400343f3f000cc0c43000f00c0c0cf1d0c1005140fccc4c7010c40cd0c000004c3f3f000c0000004c0ccf10015c00;
rom_uints[381] = 1024'h7c33113f0317c4dd4c0000440d001000c001c0030003f303030fc00c0d4d00571f0000cd00c3447000000c000305cf0d00030c0400c700003c0fd33cf1004404000f0001dc4004d03c3c37040030c014001003f0000d0cf0004103010500c00007140f0c000407000c00cc03ff00040403033005f0000000000d030103;
rom_uints[382] = 1024'h3307030c003cd1701033fc0d40d4c07cc0d40010f003010cdc3010000c00007c3110c703417c00330cc000000d101104c4030070104f171114030c1c14cf40030003c03000010fc30d300c500043f3017cc033c00073d10c51dc0100c03730c00104dc00c30451d00333071100c004f045cf3c077c15c33041c30130c05d0005;
rom_uints[383] = 1024'h3403003104000330137331300d50c04000c133333071c3430c7013d000001033034000f1c0f713700330f30334c010f01cf007c001010f4010f440510301cc47373411ccc0030001f037300f50f03300f3100314cc300347170140f40c0040035c70310030c33f140d030003314003000744000000d0c0510c310c030013705;
rom_uints[384] = 1024'h5f41103130fc05100c3f333f4c3c100f110c0001fd1cd0f000f3140030704c0c3731110300cc030d0f3d1331f137c4500c0d33cc03341000005c3f3440700000400700cdf70310f15041333035035130cc130030cc0133f0037330c7117140333013f050530c4414cc300d3d10fc01c1f114c3d001070cf0700c7c04f7341300;
rom_uints[385] = 1024'h7001c134c3300031307c04370340430c5f4c43001d0c31f000c50cd33410d030c00003c3c300c030cd03410004c000100c1c3001c0f5101ccc5003c1035c50000c3c0d1dc500007c73730000cc3d5f70405c0c33100f03304330010c77c14c40f4f0305f531334000c0ccc74303c10dc340d05cdf1d03cc1040cc0d104d33301;
rom_uints[386] = 1024'h401d0c333740000c0f10ccc00fc03c1010cf1dc0c01f4c34cc30c30f34103d007130d3700054f001dc00cc3070300c10031c71430f4000c4cc15033cc0d00104cc00cd0cf000c01f1c04fd3d0c0c1000c71344304000043534fc04cc0c41000c307fc0d00d40c0fc1f7000f130c014d004c000f0f4f14c3000c0000cccc14c1;
rom_uints[387] = 1024'h3430770034c3443333df03010c731fd405404013d734030cc0d000401341000c000741011c0c0710034303030cc0000003033500700000110000101010c00040300105f1f00000430430000303c3fc00000000c007dc00704c03c030174400400100000d4500c0f04403403003030000c030c4000c00d043c004d00f0c3003;
rom_uints[388] = 1024'h4031c3400000703033710007d5177310053310cf00d000cf034c4403700001031303d1007fcc3f00003031003c34300f011c003404003300c400431f10030340030c30130713c40000300043030d000f50000070001000041c1c0510000000c1700047033101c000c3040000000c411c0d00403030c0440f0000400d50cf7;
rom_uints[389] = 1024'h307d30cfd100c04d43cc10100fd47000c4070104111400cf00d7140703dc041d03740c3f0010c40010050d7fc707077104d1037c0c0301100541001340050c007d0700003c3100151d7c004303dd01000d3501c400d1c1037033d34031cf3c0003045c0175073c0404330003fc1003100c3134014c0714173f35d3070f0074c0;
rom_uints[390] = 1024'hcc0f004c70d07c730010cd04d4014317c3cc730343c1c04000033c0d70033f0153c07c00400040c374103d000000cc33c03110cd004007c3c003130fffc1f3cf0403cf013013170d7c0000004cf071c007c3c0000004101004c503000c40c4d014103f03d0cd440315c0113c0341333733c0cf0c4017d71337d003140d40fc3;
rom_uints[391] = 1024'hf0c4c04100350d45c430df01000f4c0f030000004f03f4301d030303044c0400000f01c0033fc34f470c754c4c0c00001c43c0450c051d0fc40ccf1303044c0311c31c0403030307f543014f3c5003013410040000030f0c01cc4f430d03300303c0030cc000010f43330f410407400f74d4c1737003cf03010f300f50c00f04;
rom_uints[392] = 1024'h3704004d43437c040013031ddf1d40370c3037405cf37004c00c304c710030031d017cc0003c034030dd0c40000dc004d03c00400001070030c03c3cc0f310030700333c001010f0740003f10d004400430003007030c000031c7c00454c703c01300307c7030131c07cd34000103103013c3c03000dcc01413f7cd41c000400;
rom_uints[393] = 1024'h4003cd70c5330ccfd04303701141701343c1c31c134100d030dcd00033c31401c013f100300410431347ccc301f01040433107c0fd334300d355030c03d000043477cf00c001100dcc00c00c303001c70403700733704035000030100c3f40700051c00013313347007311300010f3c3c3000330c0d447d1c05533000cdd4f1;
rom_uints[394] = 1024'h441f33c3440c1ccf0430d3c4f47f0f0c41cc057000404ddf00d134f0c0c1d3f3d00d30c4c70110c3503c1cc0c0d3003c40f30400cfcc70f1407c311f3030c07c400070341033700f00331f30f003430000543004134011fc101017cf40cf10c0cdcf507d7033d00534c13f103003c0c0c104501cd1d53d0fd404d1c3ccc03d1;
rom_uints[395] = 1024'h10053cc00403f00d40057ff00010fd30000cf00c104431003101400c000330103c3f3cc0001043400ff04000344047000301070f30df4c04000dc140304f34104cc040000310cf1ff01440140f3f070443300c40130c000fff00045cf00515113450003c0c03f0c3010c003d0d4000573050140044000540f010d03f1c330d4;
rom_uints[396] = 1024'h430330f1013f000303434c350101340311104400331f0430437340c0300330007101d33371d0443047d31cc030f000f751f030d00330704300c300700010f040d305411030d0001007d037fcf010340cc0d30051ccd001f00430313015f0c00c3d0f74d0401c3001c141003d0030f0f03150131c303c0d70350ff100343000f3;
rom_uints[397] = 1024'hc4107dd40c00103051000c001030c30003c0f043041dc00cc547004c340f000c30c011c1f77341143cd4c1c0d07c743000103d0c100f3cc44400cc31f4f1030cdcc00000430404c4c13c01005010d000500000004000300cccc0400dcc3100713370c737fc1c0c30014311fc0300d01100404f11034030300440034cd375004;
rom_uints[398] = 1024'h100d113c703dc301014c4ccc1c73044137717013140c31c3cfc000c0707f00ddd000010ccc4d101175dfc50c30d4307447331cfc333000d3310c1004303430c0010f10000fd0110070100c3104037010010303434f30035cc343f707033cccc3c41040705031d00707f01c040700007403c0c3f501cccf40040003d04f05cc7c;
rom_uints[399] = 1024'hc3103000fc000044000c003c45311c0541414000403140f5c01130dd10003c1ff04d0c3c5017005330d30370c400d0c410c0fff004c071100003104050c040c331030c1373f0305d03003010f0c0f103c70007d340c4000c00c1c071cc00c0f1c0c0004c407031f3c13331c0c3000370d4c0c300f0c4d041cc10c330530453;
rom_uints[400] = 1024'hc04030030dc3107000c4c40dc3c10fc41d433c13ccc400401034703703c010c370005f4c00cc44c300d0003f143cc03c110d100f00c001c4400fc405001f00000c17130c0004c40c0c0000c130131040f3d1001c1c1cd1c01011c1cd5c00c5c040c40030000f51000f0017010301100f30c1001c47050c4540c0c004d4340f44;
rom_uints[401] = 1024'hc004071000440c0000c40300c0031c3300c0d30c03c5d1c05130040143400030004c44030043cc04c13cc1440041010003434005c00cc3013133c30c4c0000c30c001030030000cfdf44c14100407010cc0c0c300c440c33c00f40cd1f05400371c0cf07f3c050000405704c0003400003140070040144005f3444304ccf0000;
rom_uints[402] = 1024'h3cc034dc000ccd03033c4f000c70c347717c3003013110d00c0400010071340cc4000ddcc30d000177dc34d010c0043173cd1f3c0c4c00c073005307707ccc400c1c30317474133cc000400415cc11c00d33c030dd114050174301041cdd0c0c03004c0c733cc3300dc01033000301000071000400040cc4143c0dd00c0333f0;
rom_uints[403] = 1024'h3150030f003c000c000c100f00ccfc100105010013711c073c175443d3004403134041101f00040cc4fc041c0f134c15017cd30d307f0130c534ffc701310f344ccc330117003c00dc00c0030fc1f4c30c3000004c4c00c300f33f04dc033c40d3043f3dc1050f003c10300c10034343d35130450c0431c3d3310f300f070cd0;
rom_uints[404] = 1024'h40c35c0c53f144705f1c1f3cd31f003030c03c003403000300350113f1050dc300314300d00500340c3f534c33f700000d1c704000f03c35fc1f143c400ffd7c33300017310c30dc03400034303d0c3cf000f000f1c01330fc1400c0000c0307c300ff0f00cfc41c070d4000300171007410304401c004300003353c1113d5;
rom_uints[405] = 1024'h300d745c100d504c40ccc17130f337ccf0303133c0c74c4c331c340700f1510c4f307cc00c01111cd7fc014c0044003530c0000d0f0000c310000c5030c01330f1f0003040003cf0000c401f3300c0101cc5300001c03000310400d4703f1300d3040100f5004c03001cf13f0cc010105c1140004c1330045cd3dcf0cd34304d;
rom_uints[406] = 1024'hc030030f00d44f3c000145004317cd310431030d00450000001753430354f30f0c003f0f0c04140000710c100157c030050314f400d30000003c01c340400c043d0030001c300300df00c30740f0301041010001043070010d00543ccc0fc00405011cfc313c0f4034c0310331301333103400fccc4405014f04143d0f100103;
rom_uints[407] = 1024'h1100007000300005400c30300033100c03dc0d4333c31c00000310c331010000f444d00100001400030fc130c0c4c01000303304007cc000d111f0304710f00345c1103f300010004c033147330050310011f0000000c00001f53fc450c300c3471730d11c1035043f034344003001f333c4c1d4040703c470130300f330d040;
rom_uints[408] = 1024'h4100703031c5c30c1331110343c4317100030040f10140c0c71313c0c30ccf7f0f3003c3000c30c003307c0c3117100104f00034003135101341341300030c7301340f0fd30444c73d0c040333f07100400403100ff00401040403d07d33f0c40053003441c330003000013000c1ccc0005707100cd304501c4c001d70c33103;
rom_uints[409] = 1024'h33000cc10013000000d111c0c305f041f434000330f3c33103174301cf1043c3103530c0d00370c44cc04cd10043c00137d0030301c330304330c04301001133c0c00000c3743003cc000c10310001400c400c330cc143100c000040f0d0f0037440c00134000c30c0c73000c001c111134303700c40004000441040c1003130;
rom_uints[410] = 1024'hd543003c000330430510400d150c0c110f340045c40f33303473c3003c033c1c5f10303c0d0010050d1401001fc003f0040c10403030cc1035041ccc44700c004d1c0dc33c011504f150103300300303300000010000140f1f10f40c0f0c100c4c15040d1c3f1c304f3d140c0410303000fc0f3473014c0330003c0d144d3f3;
rom_uints[411] = 1024'h70010004000000110cc1dd04ccf073cd435f30700c03400304f10c1f340c4f0137104303000dccc03113dc54d00030304fd14401403c030f4ff37170000f000fcdcf0f3c301f0c3c7401c130000c03d00ccc000050000f00004301d144c53030301311c00f43d403c101dc01100d001c47f0004cf013fcc0003131dc10c100d0;
rom_uints[412] = 1024'h1004fc00d01cc0340011fd000030c500030000300303c13100700330cc0df0333004d704003340c43040c0300d0ff01300d370d70310174003c4003033c01300150000cc0c030004f1341733fd00d000c01010301000430011f40c4c1107001c004c040435000043100040033000001010131000f30040313013030144f05030;
rom_uints[413] = 1024'h37cc45703051f44ccf0f003cdccd3fcf04fdc7403731040c3c0307010304303c53440cc13f100007400031450fc43ccc543c334c0f0c30c44f0cc0dfc0c000400c033101031f00fdc040d043744001075c001c4c041f404d1010030d000000dccf3d0ffc44450c0c01041034034007010300047c540c00010f000440041d00;
rom_uints[414] = 1024'h3000c400f0010d0c31c4f400300f40304c00cc313457c0f0404cc44001100057cc4740d070df341dc3d045c00300300c7504f00c0300105d4cc407315dc00c0c000d4cc000344d553d013133c070f1c01d047cf07401001fcdf1011735030cd007017c4010f41030d000f1103c000550f0c003011cc41c1400000ff041017c;
rom_uints[415] = 1024'h304d07cc103cc371007c444043d0c040001003015000ccc3df34c405c700003f0431cd00c04c0341017f070140c4c40304cc4c7ccc0c0313c54c0c041dc030404d0f00033400400ccf411301c4f00c00fc071000000d0703471703045c310c030174000373c001d40ccc40c130400cc0030303c531f50037c074000443c54004;
rom_uints[416] = 1024'hfd7fc3f0cf103c003030c3f04030304130300051d1c714cc30400030f100343040df3c30c0330c7cd0704c007f3c10405d34c00000041c300c30740170301040c000000cc0004f303000115054dc03003000001c00f4043040d0403700c03030330000f000401010dc1000c040111004cc3c4c000000300300100c10700000;
rom_uints[417] = 1024'h5000df3000304d00030cc00c430770c040d3000d034740d033c44df0d0c0113c113040303010d043d370dc303030c14001330cf3c00103c40370f01c03cc0cc10f400c17d0c074030c0c041dcdc040313040010cf147f4cd04f300f74cd37340c3c0dc333c031400331100010cc04d1c000001111dc3301f17000c0c3cf3f01;
rom_uints[418] = 1024'hc3400331030007411c000d00c10300cc00011113cc0300001341c00401cc03044100c000000f43013cc0000fc4c000c003f30340c041c0000cc007310d0000c07cc100400110cc4500037100003c000c3dc3000130ccc04040400744003c0007400341c00d00000c07dcc0034f00003400c30003434053070dc033034030410;
rom_uints[419] = 1024'h503cc0304003000cc444d0d0f4cc1400013000100300d3c07c030c3dc7c00c0dc47fc0c04c00d010d303d01333003303f00070000c44001f03040d35700013f0cc0040c0030010010401371c1c03c01c0373c33300c00514c54073c150c37c344fc504c7103d00400c13f440c5101003703c503c4c444301030153d001d400;
rom_uints[420] = 1024'h104100f5cc0c0033c41000f3dc341000005003d1117470c130714d071c04f03f30703030d144c344f000f10040000313d0f1c3011013c00004dc0f1f14c40c500300104073ffdf50d103c0300c00300000c3c0d04700cd3cd4c0003404c4c0f40cf33000407031c5300f1030000000f5f5f070f541f1f037f4d13c0350d01;
rom_uints[421] = 1024'h4700c0d300070000c134101c540c0c1000000444510403cc40c0c101000031171c5034000c04d0040110c00011f1010000401c03040410400104503c40040400170344c000004401c300d401f040000004c0c00100014100140c30010f11f7004c11401004041c0c0733007c000000053c34303534c104c10c05001150cc10c0;
rom_uints[422] = 1024'h1f714cc033d14f004307004cd03003c030d00cc3c0f101313f004101f400704c133d0000044003141d1370000c001010d500770f030c0034c00c104405007044010030514c0004c040511300c3c00573d50c100411fc3000c5c3153c4c40030f7311c03c0001c130cf401430101114cd0300007000f0300100043141100c00;
rom_uints[423] = 1024'hf00f0c1c01400004f1145d03cd0cd5504341500d033003cc01c3003100444304c0030300c34334010fdc000014344f040d400c300c1c00c770000401400000030310031437c00c0d5f000c0ffc5c00000100000170403437fc7d34ccc000cd04f00030771001d00ccdc34d771ccc4370cc3cf40c04700401040d3703c104304;
rom_uints[424] = 1024'h140f003d00c030003570300430335530400c10173130c000130c0ccc50331003740c10403c073430343000c03c130d141d37431c0c71004d101533701100f00100330c50c414f13c10030000030c1000c000400c7d040433043000301f303047334031051c30c3100031c003113d3cff0d1f100cf300173c3c1c3000333c0c0;
rom_uints[425] = 1024'h4c0f14043fc503401f001c074005030130030c343cc000010f4330030c0f54135d0133cc043c103c45030c01303000414cc31fc503350dc043000f503c044113c431c00000401cd3530000c537f540030000c044c5303c0005d43074047cc00c1c03140044041130343140d000f5353c1c3004730001f34700000044003c100;
rom_uints[426] = 1024'h3101c4ff031040c007d3170f3c7301d77300f0443045030341d43711f4c3340c047c003c0c43030d315fc04c134504314370031d30c304410431d3043401030c0dc304c0c7043100f3101d3ccc0c11f0cf0400440000031300330c050c0100000111c03015300c4010f0503cc30070003f3000003c045014fcc40f1133001000;
rom_uints[427] = 1024'h3f400c4d3005fc40001c100300f77d17003033c137f03c13f000c31431c0130c0304f030010cd43017003c304d34070000f00c4c01401700c73c1c00000307101301034d030003013040000d0004fc3c00c000c134300c100dd10d0070753003170d04031031300c447310031131310044c430030013c0034704330d0d13110;
rom_uints[428] = 1024'h31000c030c05d04000347300f70c3c30103131dcc4f130d310370dc00f74000043130c000031401701c0040f1303c00111d03044000c010ffd010f0fc0f100f01045033c041000f53d004c13d31301401011050c450503434c4014147cc3c0005f730334310c4f0c0013071c00c410043c00300c000304330fc0100037037001;
rom_uints[429] = 1024'hcc040fc000c5030000c10104004cc30d000fcf301333cf4f0c04404001010f07004cdfc000000f0470433044414300000c4740c4d00dcc0cc0c00c0c0500c00300cc00cc0043000cff04d4700173c040c411000300004d11cf1cc0540f04300141f11000cfc3400c05c4014c0340131400c0c0130444014000f4014010410c4c;
rom_uints[430] = 1024'hc1003c0304f00310003c3ff0cc1404ff01cf143cc3fd301040004dd005f3000c1740c00514fc0c00130c400000c433c10003003c130700cc000d07c70c00103c0c3030cf17000337040c001303dcc007cf003c03030c40030457030704c0cdcc57c144d17d0c0710ccccfc470013000f40f1f1cc00d0c00c033dc40c4f104011;
rom_uints[431] = 1024'hd0034c70c04433cf00c000c4c30140c3c03cf0fcc4c113403010cf0c40ff7c0450c0ffcc74c301103f05f010441000ccc1f45043307d04c03fd10440ccfc040df000ccf00f0c0400c0c4070040030313f03c00fc4303004033fc070c00000454011c04f0c03c0000f057c101013400304403133c330c0513440c04000400310c;
rom_uints[432] = 1024'hc0c43003001001100cc3330c13f15010c0c0f030f00cc30d3f04f33030f300005001dcc003c4501371530f03433005c1033051000333000041005303303000314c13f5c4fc4c5c3cc1c000c00105100c0153010000c0c04154730331dfc003011040c30011f0000f4ff10035033000300331304300503040fc00c050c330703;
rom_uints[433] = 1024'h34140500404103330ff31001c3330004430331004010c0dd07300c040c040144c551c003434305543dd0341d103711f44110004f34003c0f00cc1404730330cd50403004000c0d13f700040cc071c040c17004710110430040443c0334c1073703fc403ff3c01000440d174000411110007071c4000044f0c000cd1d001c174;
rom_uints[434] = 1024'h30413111430d0010301c311d4ccc103c305317031c1000f300c50430c43d03f0f0305004003074c1d55ff0c10dc133070070c131000d3c3c04303cc03f134f3c7c0030c0f45c7110d3c005cc30f04fc0007cc00c00c04001707cc01c0c04f1c1f0c11c334317c4330dc15c0cf01c000cd435f100c034f0c0f0c1cd7050103c34;
rom_uints[435] = 1024'hf1ccf4000f0130c00044044000400d1070040c0f4cf7f0013403ccc734c0f0d70050f03040c0d0c14c10000104330cf04d305cc130cc1100fcc157013cc44010dc0cc0373c3d1c0000d0c030fccdc0030c10004c0c3150001150734401f3d03404104dc010f4447c07fc15400c40fc3743f3f033f0c00047cff44010540c103;
rom_uints[436] = 1024'hd00040011114fc140031311c3cd113c53c3015000ccf0f30c040040051f0303c3ff00c0013cc34f034ffc1f04c470310f0cd1cf0d050c0f3000ccfd3f101d0c0c430007c3533f00c5d00c4cc03cd1d04cdc44cf0000d0070c3c450400ff00f40f37315c14c3f14f340130cd00c1dd0c400c4073001033f331300010000454305;
rom_uints[437] = 1024'hf4000350104000103d017c303c44c040f4f000cf3530000d314dd4000c4f343054c7f00c1040f40304c0031004100300000043040004fd30c4307c0705f011370005033c000434f0030140071404c007010001c0070dc0000c4c4cd004547c4000c00315c730100031113c300000001fc00000130050300f004044c00051cc4;
rom_uints[438] = 1024'h3301c3c1401000c3030334cc0343cf0300c001007401c1c10c050411f0540000f53c0c00c053f414470c00c041c03053035300110133330034530ffc00074100f0fc041c00c303470010c14051017cc001300070415144c0fc371040cc011304f3077053030100001cd310000040015100d3101c10041000cc105000f000f314;
rom_uints[439] = 1024'h44d0c5dc004c0000c03c071f7000f040440030c44014c5d0030cc5d5fd0700501d50d403cc404c017417401d0001110000c0cd4f03f010043540004d00040c0040c0000ccf0140000050c300cd70470c403400304054040c44003c0100c340710c01400435041cc4c0c1d40c001010d4000400550cd14c00dc0131005f001cc4;
rom_uints[440] = 1024'h400003f3030504c70304f004100d03001100003cc14003cc55704d0311441007cc001003003103000cc70530c01d4f400c3503571030131f0040c30c0040133004c00303d03000c03000f45c10c100040440400000000c03040c01c100101c0cdf0cc0403f03000cc00c00d0c3f004131301401400415010004d4003c331c301;
rom_uints[441] = 1024'h3f000440c1c001430cf0c70c404f330c304cf340043500d0f0d01c050300100cc0410d00333cdf0c0f05004001c0000c40710fc000070dc0cf11c3007cc000410040010c00001c300f4300700d074c001d010d4c007104d01007c00033030ffc37d3040d000d05350000417303400d014fc0c34d0300f40c0fcdcc14111c00c0;
rom_uints[442] = 1024'h4c401fcc033c3f50100cd00710f17c11c0404001c51f0dfc000001504cdcd400303030f070d3c40015cc470ccf00c57034c0c300c031040c010ccc1fdd40040c0300141f00300001100c000000314c4cc04c00f00404c0fc0f13c0c1300440f0f40c000103c37035c0743c0530f400047300000f4104f313040430000c15701;
rom_uints[443] = 1024'h340c10044013703d30311000c710c4003c03c0f030003003f1fd350034034100004d340370713130dcf01500c303140000c070c000f0cc7c1100c00030000070407c0030300030c4000000c00c0dd3700100304010f0000447033c13c0700007317000c0c0101341d0010000fd0737d070700c41003000d331110d1100c135;
rom_uints[444] = 1024'h51400d0000300100ddf70010c771d0f4300000d4003030f04d30713f40330330043c00303010d014d40000d03cc04cc41400010c3d070c3740d400040000c70504c34c3f0010d100114d053c050030fd070cf0c3000cf0c0c73010f30dfc000410c003503030f3013f10c43dd03003c0033c3c0d0003d0301c0000d301d000;
rom_uints[445] = 1024'h3037cc311700010d0c00d00c1450103040000c1d300000030c3000fff40417d30770030303c00cc4403300c0c100004c3c114030f040107c0310c0c000c00007044430f0005dc30050c0c3c00040070c01410100c00000100c01c40cf01d100d00c00040c0c000413003c47cc0f3301c010070300050c3c1310000c03f433;
rom_uints[446] = 1024'h3f77407c00301c40503ffc0d00d3c17cc4c700c03c03711cd030c0100030057c7104c70301301d3331c00c410c010005c00f0073d04f001010cfcc0004c3000340dc00f0300000c34074504010000f01300c00c00303dc0c0dd000cc0143f10700c00c33c30441d40f00c30030c0100005000004701107c041f3cccccc0130c4;
rom_uints[447] = 1024'hf400d031f4300431007300f00c00313300c103000331005ccc40101000001730430df000103313331c0037033000000310c007f001400c3010044353c7cd0307f700c003030000013003f3035030f334f3d10f000cf05047d70c50013c0c4c401c403130000300010d4c40003040000003300014001c13503c0140033353400;
rom_uints[448] = 1024'h5c40c00003f00000c07c000c0c0c100000c01001000c000000000405c0300000c0c0d04c40000c0000300000f0040c1000003040c0044000001cf0f14000000000004300c0407c3c1040c30001001000000040c000000030c0300004c000000000c0001c000300000040000040000004000c0cc500000cc0c03c000000440000;
rom_uints[449] = 1024'h700f0037300100c010300c3733000000000c100030003400000000000401103c37001010cc011000cd030040300703100301f73001f11c0003500004004c0000c00c4110c50300cc4033003030311c040f5100030000000003000030430100000430311c5f1330000000003000cc00cd44010000f40000014700000001001f00;
rom_uints[450] = 1024'h1000c0000544000003000c000d0f03c043300000000350c0c34000110000f0401000c0314c001000d000c000001c0f300001053000400004c0100000c0c04044c00cc03c001cc00c4c04dc00030004c00703330070000014043000d00043000030000000000031000340000000044140000103c0c01070c1101130df3000403;
rom_uints[451] = 1024'h300330000000c00000000300004f400300000100104030000000c00300130000c403c031001040001340030000c003400400000000000300003100d0030000400040000103000041d1000000c300000c134400c0400300000700000300d34100710410c30100c000300d100300000310040000c0c0004000403040c010004003;
rom_uints[452] = 1024'h41011000000140c00001040300004400000000c301c0c000330005400040014300003cf0000370303030004cc030c0000003000040c3043cf001005300030440000000d00003050070000f701300c000000000c0001030040cc0c50000000000701300334d0000000340000000c3c1c0000040000300410c00c0440000f00;
rom_uints[453] = 1024'hd7c000c0000003c0cc4c70007040fc401000033000404cc01070300070407000300c0300404100000011c03303700010410004c0c001c1003000013340000000d000d0c00040001300c0c0c0f00cc0000c030f00f0c1503c0130300310c00000014130000300d000c0700003c0c0003030404000c4703030f040000100c0000;
rom_uints[454] = 1024'hccf0c010000cc00000307313030c413330ff00303303dc04004030001437000340000000300034003300031001000cc00001100c0141c13030c0010030f00000004033c30303313cc4c001004000000000710f01c0017041013c0333d000000051000000303c00003d0c3c00003010330003000000013c001040004004000100;
rom_uints[455] = 1024'h14000000350d5400000001000fc000c34000000033c0000c347c0000000300101030c003030300034000440000000c000000350c04104c30000000100030004500100400004303c040015330000011040c050030003fc0010c30000000ccc01703000c000c500000000f100400010c010001303000f300010000000c000000;
rom_uints[456] = 1024'h4c00040000004000000001c01400400303000403300001c00000000400001c00000000001034000d100400c00c0f4000c00010000c5d003c000c040000000000000000000104070000001c00000000000000300300c000310010000014000110040000400c0000040000000400000413100c000c000000c4040c011003430;
rom_uints[457] = 1024'hc0003300f40c030c1333001541001047003c01cc0040030d5010003003003010033c0f0707000410030cfc0000c3000c0003000103030710c0144003000300c703330c3cd1104d0000004c03c30044c30c440700300104040000000c0c0c004f1000c0dff304030d3c00000010330000000f3130070305041430000000000;
rom_uints[458] = 1024'h1c00cd0000000303404c0330400100000700000000300000001013301c000031040000034c01003100010000c0000300003c00000c0000100000010040030c0400400f0000300000030000000010c00001030d00000000c0040030040f0c00000000000000c4004f03100403000c000400000c0d004000c14300110cc04000;
rom_uints[459] = 1024'h104003f0051f3304450000f301004c00101c00000300010c01d0400c01cc00003f3fcc300011000c00f030000040030c000004003000300043314c4000400003700000d0f005401cf0104000030f003000000c000030113c3070c05c0000141400404f400ff0300005c00030000f300334041400045401003414d30000007d0;
rom_uints[460] = 1024'h54c30030000000030030034cc141050c0510004c30000101000c0c0f4c0f10003101144000001300c3000004303c0004300040c00030043301000030031033000005141004c000050000030c0c310700010430010000003004353c0c04305400310f30d30000400d000130300c300330100400100001300004003000343f00c0;
rom_uints[461] = 1024'h3000c1000000000301000c0400003c00400001303000d3010c04000400003100c50c0110d00700000000031000040100000000100100000000000100130000030cc00300310000000013c00000003cc0003100010700404000c000000c131000003000014d010003c4104013000000010004070010c404000000070000700300;
rom_uints[462] = 1024'h1000c00c0c00300010000400030000c00003000004030040c0031005cf000000c04d005000004cc4044401001000040c310041000444500000040000030c0100050000001004300030003001070010000334000f00cc3c303f0000000000c3c0000f0c000010440000f01c0c401000000c40000c043000030;
rom_uints[463] = 1024'h4014503c03c07304300000003004310000701503104043333010100011501c00c0300c34c04403001030c00c3000f340040000c00000000f1000f01040000cc00430044c0c0304c0510000000c3cd30100c00000c40004000300000030000c00f00c3450000c0000f3f0300000c4100003c0c0030000c0c0010000037010c011;
rom_uints[464] = 1024'h303000300c3433c03c00001c3010000100c000001000c0000344070c000011031000f0c00c005c001173000c0000f11000000c30c010010400c10010001030303040000450100000c000f0000001c00c0010000040001000c5000001003c4c1003140000c0c00000004140000000000040400100334000000c0c01404301004;
rom_uints[465] = 1024'h400100040030cc0000c300000c13003000000400dc0000000040000330c0000000300100c00000c0000000300000000430c000004c000c00030004040000004c00000000131001001c0000000000000000c00000000000030000004000000003c0003c1cc40000000000000000000c0000000011130000004000000d30000;
rom_uints[466] = 1024'hc000041c404c100040cc4030c040d340000f00c040ccc1140cf530054001c4000700c10c304c4401371c00c000340330301cc00c0c0c00ccc0c0000403030140004c00c04444100f10c04000050300000c40c1c34d00c010c0404d43cc110000c0f04000030cc4010cd00c00004004001100010700043c001440410040044cc4;
rom_uints[467] = 1024'h3104000f000c00004c00000f41300110000100000031100330070004400704000300010000cf00001430001000130c0100f0430100030400111103c3c001c300003c310003000100100103c0030c41000c00000c0041c0030400030440100000c3c03305410100000c51300000c00003c0000041000400000f0100703fcc0013;
rom_uints[468] = 1024'h40000000030c44071f0c0000c00c0cc0330000ccc01004000405311301303c100c010c7015040c300d30000c00000000f11000000300c034010c04dc300000300c300000043030004000000000314000f0000000000400003cd03103010c030400303c00000300c000010300300d31100013304000140010d0000000004314;
rom_uints[469] = 1024'h3030030030000100c0003310c30000000000003000100000000004300305007330111310001001c00c00000000000003cc0c01000300001101001333d000003100003073030c100000000003010000010003003100300001010000105000030000300000000000c003003000000000000300304c0000100310000003300031;
rom_uints[470] = 1024'hcc7030c0000000003031010c0f54004104100300003c0300003330301000c00cc0040c000100f400000030010100100c0000103000001140003cc5030040000101c4015cff0f03005c00c41403003c30c0000c4004000c040304004cc0400c0c440d040c5c4000000cc30104000000301030000c000001000300004000031130;
rom_uints[471] = 1024'h40000003000000c000000010000000000004000c01c00000c0004100500000f43110010000c0434400000000000d0003400040000c70000d3003044d00c000000140000000000cc05030040001430001400000000c00000000001004404c04000000000000000300040000000010400000005000000000004010400001300;
rom_uints[472] = 1024'h1000030c000000010313030004100010000400001000010040c13c00001034000400030004c000c0030000000030000003000000030c5101040001001000001f004000c03000030310c04000300000000040000000010010444000000c00000101070004000041030c00c01c03000c0030700c000100000000c001031100140;
rom_uints[473] = 1024'h50400110330000000100c300100001004304c00040434003000000000000001010000400c000000cc101000043000000100033003400c0730100011c30000000300000f00300400000001000000030310000000000100003100f000400c3000040000000000300c000010000f0000000030340005000401000004001000130;
rom_uints[474] = 1024'hc100331f00040040045c400c04c0d0500c743005c00fcc00010000003c3c300cc0004c0c000c00070c10310003000430040cd03030f00c007144130c740c00c00c3030403011540401400ccfc4040003000004000000101cc00004000040000c0c0404004030cc010c0c04004400f3300c0c03470c0c00c401c00300c440304;
rom_uints[475] = 1024'h3010400400000001003103c000304401000300000003440000c0001c3410030034030000010010030d00000003000000001c0400003001400f014000030d0000510000001300000031001130000000140000300310000c310110000d44000430000f100c013cc000cd04300c00cc101f34c3003000c300300400000000c00d00;
rom_uints[476] = 1024'h300400000000c0c00001001050040000000001043000030f0010030c000c30004004f30000000000044030000c0f04100000104300003043000400c0140000000000000c0c404000c10030130c000000040000000c001004000700004033000c4300000005000313000000000301000310030300000353000010000114001100;
rom_uints[477] = 1024'h30000450033510034c000cc0c1cc0001000c0c00003300453f000400040c03001534300c0300000c0403001400000300054003041000000d03f0301dcc040000000003001c0030031c04011400003007010000c70401c00405c0c0011000c001c030130f00000103030001000314044010000043410c340010c000040040c00;
rom_uints[478] = 1024'hf0000c44100c100cc015034c00dc01000d0410003004404f000004540411c0040c044000c0010005c04c00400400c3c00c504c000000c035cc000004c000000030300500000c000450000cc00000000c3000000c00400000031000000044000cc130c00005000c0c01000c0c0c300040503000c000000c00500100ccc404000;
rom_uints[479] = 1024'hc4100000000c0410c4000004d040c430015003114000c333c000000040cc01300410103c01050340170030430c01c130004400c0cc0df000c0000000cc00000400c0c00300c4001034000000417170c0c001030001001044000040c000504007034401040000c00100004000f00d400000000000ccd00000031003040000300;
rom_uints[480] = 1024'hd73c0c4300330003d00300c0030044404f00000c0c314000d0010700000000c44130c00000000000000000043030000143c0000c00000000040430500000000000403c00000003c00000400341000040000c00000000000300c000c00c0000000000030000300c00c10450c00111400c00c07030100030c0c100000404000;
rom_uints[481] = 1024'h1400030000000040030030c400f00003000c01010030470040c0404000030000f0c3141400000d000d03100000330000c010c04f4007f03041c0c00003010000100303000000c00c0000001003000003100000004000410c114100c00400c0f0400000000000430033040c000000c00004c3000003010001000004c0004c0c43;
rom_uints[482] = 1024'h34340007f000000001000010100010000005003003000100303043140f000030000100000c0100040030340000000000030003100000000c0000031700000c04000005340000000500000000010d00300d0000000310000010030040170c0030000013010000000c00000000010000130000c333030f300000033000033d05;
rom_uints[483] = 1024'h300000c07040000000c04401030000010003000000c3c1d0c00c03003000030001c00c000140140400d3000000730c0300c00007000c000003c3054c0430001004c00043c000100c01000070c030000000c0000c04400005c40000430044017c344005001000040f030d10000000000004703000f000430f00004503154504c0;
rom_uints[484] = 1024'h3003000c0300003d010c00f10331407001040010000330c340100031030ccc0000c0003d13000530000000d4300400410f4c00000003000001c001000c0000003000c003000cc500100000300300000000000100003313004000030000000f00c005000000033003003003030001104c1307c0100300c00c0cc3f0000001;
rom_uints[485] = 1024'h400000000000140f4300000054c00000101000011040400000104040c00001004c00c40000c0c00001104c3cc0c0030000100000c0000000013001c10c041413000040c003400000000c04c00000010044044c0000c0c000003c000004cc04c0fc010c300000c300040310c000c00004f44030c03000c0000000c0001c0cc333;
rom_uints[486] = 1024'h70c30000004503c030000000c10000000007400c000f00c0030000040f1003070100d0000300000000c03301c010017041400140c00010c00c000100040000c3300f000103c0010347000400000c000c01001001400140003d4044430c0c1003c3c14003c0c0011010c00003010040400c0000c733001007000040d0c001c00;
rom_uints[487] = 1024'h33000c001100100100135013c010c04003015030000f30cd00c0300054440303d31003000c03f0351cd0100010fc00d00d100000010c01d403010000100003300c100300033fd0105305000031030d000c0330004c000430300034c0f0000000f4000077001000cf0cf74103c0c0414d003030330430c011033004c00514301;
rom_uints[488] = 1024'h3d7000c3100f1030330304000c17010300040100c3011d10c003000001c700003303040c00004f30041300000400007100c00300c0037310c1000777040400003300303400005010c1300000c000013403000c030310500300070000010f00000734c3010000c00400000000300303c300040004cf000047c40000300303c404;
rom_uints[489] = 1024'h3000000000fcc03000f003c404030000000001c00c0003001000405f000c0000071000010030010101100000030000010000000300000100300000050000000001100003003001003500000300c000007000c0340c0300000000034304040100040301003000c4000f430000300040400003000040000003010043c4100c0001;
rom_uints[490] = 1024'h340040cc000000000dc1c0c000300d000000000c00030000010000d00000010004c040300001401070c030d1c04700003301c0c00c0040004041c030000001000040300c7000000f0100040000015000c040007c00003000033000000000101401000030033000010410c0f00c0000000c000003040500030040c0000001d00;
rom_uints[491] = 1024'hc00000000100d00f10101c0401c070070000330c0707c000101000000100000400070c040dc044000050300000033004000c0c0c010c0004df4f00003c000003431c300d001c0000343310c01410000000000000000c0c000c01100437040000441c0c03430000001000403303c0003001100000c000000c0004030c1cf04c4;
rom_uints[492] = 1024'h40400000c34004000303c0007000c300030310000c1fc00130350c00cc40c000010000c0000441000304400001000c1c01030040c400d00003000400100003040440000040034c03d004c10033000000004000034001000004000040030000013300400300c401cc000001000041010000400c300000400100010004000000c;
rom_uints[493] = 1024'hc04503300005031403010130003c30000000c04013c3c04000c7003300000c0000400300410000300070d004001010104c030004c1000000d310304000c3c00100cc0c04c0300700cc1405100413000030110010c0000c30000c3300000030004000001c100343400000701cc04000000030301310040113003000003c000100;
rom_uints[494] = 1024'hd1000100000c043df0030303c34c40d00cc040c034d00c0f0010010043c00000c00000c00030040400c0010c03403c10004000c07044c0c431c00030000000c0000000c10000010040003000004d404100c3000000030100403003300401100040034011c0330000c000c0000031003000000000c100c0c0400040c00f01c00;
rom_uints[495] = 1024'h400403000c03000c003cc00004c0000c30000400c0000c003f0040cc0c015530cc0000000d003c0100000000000c0000040c00440c003000054cfcf000000c300c0000000004040000010000c01c000c0cc0000c0004000000000000040401004000010c4c000054c1300404000f0000003c4000010c440c0000000c4103;
rom_uints[496] = 1024'h100c40c0000000110000003000c31100000000000040130100004f0f003f40c000c01100300c4433300400c003033010d00301000300340303000000df0f0004c0c00300000101000010001040000000000400c0300c300104000030103cc00310c3003001000010300000d0110000330000000000f000c00030000530701433;
rom_uints[497] = 1024'h4100000c03c000000003c00000400013030000003101040300010434300001470cc300c1cc0001000000040000044cc030ccc300c0c000000300c0000000000000005010100001000010000000040001044000700701100000000070cd10030000040000010003011030000000000043044001c0000101cc00cc0;
rom_uints[498] = 1024'hc000400300d000000cc31001c03103d00000000c00044300c00453700010300003c4003c00070c0144c01000000c300000cc031000c30001500000030134c007d0d0c140010001c131c01f000f04c100c41000001cc0000417000c04c300000300117000000000000000000c1100000100001000004f00d1000c00010c40000;
rom_uints[499] = 1024'h300c0f4000c0000c000143000111000000000000300070000010000000000340100100c0f00cc0000f1100010100100c0004010c00000c1003000043000000110004000c07000100f04000400000000030c0000400000440c0140030004c00001041000001000000000001000000000000033307704000000cc0000005330000;
rom_uints[500] = 1024'hc0403c0110000440040300070dc130000301000000c403004400400103030c003c000c0040c3000040f10004c04000000c000000014003000000303c11100300c30f04003300011110000c004000040cc0430000000003000c0100400040c00c3331000000c340030507c1000100d0140000070003030f05000003010000000;
rom_uints[501] = 1024'h3400400040000000f10000c0c1000400000001300035000100400040003c007c100434300330073004c00300d010c000341000001c10010000000304740c000300c00430000501000440004000000003dd0140000041c04001300c110444cc000cdc000003001000003400000c0004000c0003030f400c0c133040000c40004;
rom_uints[502] = 1024'h30c430001001034000c000303c1310300010000413303000003000c030300003011c00040404f00003c030010000100003400000c00c00c003004f001000c1001c01d0007033031011001043300300400103c31f0001000000100014c0c1000013330000c3000400f310305000033140013000004000d0004000d40030141000;
rom_uints[503] = 1024'h41010000004000010300330c0000d507000100c11c01c103c30305c0030301000c00c0000000430003070c0003010c4000c0100000c000040001030001003000000300313300400d110d010c000041034000000c700000000000c0000d0001000c004044010103c033c000cc00001004010001441dc040031d01010003000330;
rom_uints[504] = 1024'h400030c3000100c030003000c340c30000000000001000001070010010010000c30cd4030000000100f301c03000004030310000100313034010000300003300c0100010f0f300000000c00030000004f40430004011500300000000030c1d400f00001003070010400d0300003001301041513030405330c041110000300c01;
rom_uints[505] = 1024'hf00003001c3003000000003004000000000c040c0040cc030d003040000000c03400c000400c000c0300401300c0c0c4001000400c000000c10000070c030003030c000030300000c000000000300000fc01000044000c00004000000000cc00010c41c000c03000301404000000c000c04000c00000000c01c000004000100;
rom_uints[506] = 1024'h340003007000f0000d0d000c0d14010c1010001330333cc03000003000c0400130030000400000011d00300c00000400500070003014001000100c0111004030001100f0000000d0000000033000043001000300304c4cf000000000040000000c00100100031040400c00000000c00000300034034000c040000000c01000;
rom_uints[507] = 1024'h40011c3400d003000c000000011c3403000000030100000c33c0050c03000000001003300300030c100100000401001010070c0c0c10c300000c001303003000030703030003010040040000000100000f00100000000003000301000030030c0400000000000c0d300c0403c000010303030113100001000000000030000;
rom_uints[508] = 1024'hc0d000000400310001c31c403000010001003001000300000300000040c3030030430300000000140000544010f0000001100010c00000c000c0400141000c10003c041c01017100300000430100000c3000010c001040000c70103c04c0c01043100004c0037001c00010400103000013100001330410004000100d303c100;
rom_uints[509] = 1024'hc000c30000110300c300400c00030001030700c000d0c000000000c04f0d00003c00400000400100430040000000000c0000405000030000000040000044c3004100040403c0010130000c03c00140003005d300110000010100000100c0001000500c000000c00300c000000010400303101100cf0110000c1010c1c0000300;
rom_uints[510] = 1024'h1c040301300d0000103d003c10340050303400313c101000000103030000c41030041033100c0011301010700030030000000000040c7710d000330104133000131c03000031000030340074031000100003000000003010103300300300010034013c0000070034001c000030304000100c10004004700000103d000cf30000;
rom_uints[511] = 1024'h30000040140c1030004000003015000010010c0030000c400100c3000000c003030cc003400300400c30300300c000f01f00300c0570c000c0330000d00000030403000003c0000100033300004c003300c00000000000030300000000404000003000300313100001400304000000d10400030030000000304000004f13010;
rom_uints[512] = 1024'h404000cc0030c00100004030c00304410000400031d04c300303c0000040000030c0c0000440030030c0000100000310400030c0c03013c0004f300c4000cd00000000014043003050010000310dc3140c30001103c3003000030000c101f003f000000c001100030c00000100310013000003110100c0cd00303300c170300c;
rom_uints[513] = 1024'h300000c040740000000c304d0c0c0300000f7010003000cc000103c001000000040000003400c000000001433037c350033c0000100000c0031333000c3c1400004000100003003c404c3000c3c01000c00401c0001000003400403400010010103031100fc304c00014300000c000004000000000040c000c07010330003000;
rom_uints[514] = 1024'h400000c00000000000d000000040c004100000103300050100031140c000c000030c10000503300010c0000103030000000030004000000000c00030c000030004c00100c0c0000030004c00030000c4c07003000000c3c11000f00c43c0007c010000000000400f43000000c000c0003003d03000400000000000d000010;
rom_uints[515] = 1024'h3130c00040400403010000000c0c040c000000444000030000ccc0c751500f0100000000030000000000400000cf01c0000340050041000000c100d1000303003444400454404c03000004c0c0030300404431004440000003000000c4c3140031d344c0303010003f040000404c0000c00000cc0370f0c000031c00001cc4c0;
rom_uints[516] = 1024'h14d00d030d0403fc37004031c0434040c001403c1c0001f30000d044d3501071d010440333004c4c040004d00540000054f34d34c031c0fc4404050010c004c035c01030737c10030300034040410040cc0003c003404301000040ccc03100c000c4004c14010000407000300000d4cfc00c130c3100d003000041040030;
rom_uints[517] = 1024'hc30004c001c34000000c30404003c400c10000010cc0000c000000400c0004c0040303c0000c304d000000000f400000000030c043c000400003000000440c44000c004300330c40c00c040000000300c000000000000c4040000040c00000400100c0000003000304000440000400000110000000000000c000004441000c0;
rom_uints[518] = 1024'hc000007100d00000c01413c44000403003c00000130c300000c0000000c004004030357100130000c010c0000000000000000cc00543c003003430c0c3c40000c000c000030000017000c00044300000001000000c40051010c0400030300000c040030400010c00c14000c000c0c0000000000000c00000044000001000100;
rom_uints[519] = 1024'h4030000000c400140030103c00c03010000c003034300400003043000100f1c0100000317c300100c00040000c0003003500400000300303003100403000005100034010c00c300c4100000400030100c000100004000003110000004030300530000000100100300107103000100030000c300110003000300000000cd000;
rom_uints[520] = 1024'h131043400013001400c01030000d40140043004140734000cc03000031033433340000305004004000d0c440d0c10544000c0003000d0c0030c411313030000300c000333015d53c71001300103000d003cc03c14f030010000d3c00400000000100c10004300000cf70f031040000004033000300c00c0333404cc01c00c030;
rom_uints[521] = 1024'h1c0c3000000cd0d000500040440cc0070c00104c0c40c4403c0001f00c01010000f10100000c000054c00000300c40401007c0410307000044000053100000d03303c0c0c0c00c0010000cc70000c0c04003700004c040053000044000304504400001030530434c0c44c0c31c0000037003c0c404440000000f0000dc4c1;
rom_uints[522] = 1024'h3000000050cc50010304c00400530000000c00000400c1001100000003c0000c0310334c0401c0000c0f1000030110001000050003d0045000030000000004000c0c750c1007000c0000041dc00400310c0001540000400003141000003004000000c3003c4c300400100340000c0001300100000004400c0000cc0c00000c0;
rom_uints[523] = 1024'hc043d00040000011c00c40010011f000000004c0104c000140400310c0000c00030300010000c000000000c000000004000010000000400100304c0c300000c300000001000100c103c0130000c00300001000000000000034400040000000033400010000100000303000043300000003100000044130503030403000000;
rom_uints[524] = 1024'h400700340003050703410300000dc10c30100310000d0040004cccfc000f147c7c01c41400cf03301000130400ccc030010000c301d0140000000000011c30004707100f300c000000c000cd3c0733c034010010c000030c04f5c00c0400c40c010c031403503fc1134100010c0300000000004c300110330000c00034ff4003;
rom_uints[525] = 1024'h4ccc304031100c3041f3c00000400040300c30100304c000000400000d00c000c00c00404000c3fc00000005040f003310cc00000000c00100000300000cccc003300c04300c0003000405003003c030c40000003340c1c03004dc140100c30034000c0cc00031000010003000000000000000c40300c0044c00cc04000d;
rom_uints[526] = 1024'hd0cc700c000004001c00034000510030400c4000001000c00c000000f0dcc000c10010411300701c7010001004710001000c0c0000c030040c003c710f10000c3000f404000070000000000c00d00d00000030003010000000340c030000c0c000400100d00400f0000c104000000c300000010330000000c0101c04d040;
rom_uints[527] = 1024'h40000c0000c5d00103001303c4570300041100c0000400000c01010c0c0000000c01c010110030c057000f00003d41004410cc000d00000c0173010505040c0cc00000410c0f34041000cc0034013000c00c000d01000c010003010004c0f00c4c3040003007000c1010c01000040000cc0c00310c7000030000c0040503000;
rom_uints[528] = 1024'h43d00050030143301000c0003300000040c010d340103040001c104c03010c4c50c0c040c030043c0030c00040ccf000c000d340001300c000c3300c1010000000403000000033103c0c00104cc000004110000040005dc0c1030000c03000000030004000f4cf00c030c00c0c000010304300c0303030c00404300401;
rom_uints[529] = 1024'h40011300014304c030c0c0400f0073100010703030000004310105100030001033031000c030010143c403001010010c70103140000043010000000cf040c00400c300d10000301c00017040400000c501317c0033004300000cc013400cf0400d00030000100003007040014000000cc0c0010000000003f0304050c00300;
rom_uints[530] = 1024'hc1301c0040000c3000400000400f0c000000000dc0c310000030d00001001c00033100100000c00c10300000300434001410301001430030030c0c00301000014000f04c3500000c30c000c10000001000000400110050c0030000c0100430c0c040400003100000c0000f0040300010003030100003143300050110311000;
rom_uints[531] = 1024'h1141300cc000004c0c4cf0300000400000000c00000040c00c30400c0440003503c3cd3c0470043700c0000cc04000400000c00130d000040c003040043400000310404040000c0000000140cc0c00c0000013100000300300c000c0301010000c3403000100000013411000300c400010000100d0104003000030f074c14;
rom_uints[532] = 1024'hc0040c01fc140410c000000c004000000000100c00300c30c00410300044c50000110031c0000301040001030010000c00000000000c5000010050000c100400000c040010000044c403c0100c40004c00035000004005400c000045000c010303c0000004004cc0000001000000000030300400cd30400c0000000310001;
rom_uints[533] = 1024'h440031c001031033f000030c34cc47040100000700010c3d0004000010001f3004004040c1000ccccc00c0001f400c000301000401f00300c30f4010000030c0c47305c4f0440d40040f440c3400000000000004f000030100df000404031f03011c0c47100c0004000c10d0f0000130040000cc031cdc0400c00c04f14c;
rom_uints[534] = 1024'hc00035400031000cc000005010300000000001030c0000430004c1000030d0000000c100030000000040000000040000000c004c0000040000400000000000403340004010100004030404000003474000040040014000004c040c30000c0040c0400fd00530400c300140c000030000c00700000c400330c100000400310;
rom_uints[535] = 1024'hf101000110c0000030cf00400000013003cc0000000f000ccc31004f30701000300c140000034d400001003400000430000004000010000033cc00c0050001000003000c0000000303440100710100000030c0030500c0340000d0cf0f0c0000000041003f03000003f0000c01050130440003000000000400301000;
rom_uints[536] = 1024'h10000c001000030000000100040104040100c0000303f04300000c40074103000001000000c004000000030300c130cc01c0000d00000001004000000000c00003431700c100010000005004c0c300c3c300c3000303c00703c000000c0040000000004000040c00c00000000d000003031000c3000003300300c0d00343;
rom_uints[537] = 1024'h3000c0c1c11000d000c100000c0cc034000030300704000000c00c0300d00010330400000014003333100000000000401004030000001100010000000000304000301c10001040c040c001400000000010303000004c0000400000030c100301c0000c003010000000000030300c00c000001000003010004304;
rom_uints[538] = 1024'h3f0031000001000010103c1000005000000005c003f30030400030000071d340103000010f0000401001d00300030000003000000c01000040330100f0c0100000000f301005d001000003c3400330d0c000c1000100d3c000300000003000000000001003c0300330000005100000003cf300000dc010000030401000134;
rom_uints[539] = 1024'h4000000110000000100103000c1000433c00000c74000030000c04000440040040030401cc1000c3100100040001031104011000c00f0000cfc00040010010c04c00110cc00074450000000000101000c000c0c00000000f00c0401000000c03c000434304030130030001cc040004040100040300c00c00c1cc000003c0;
rom_uints[540] = 1024'hc000c13000c0c0003c40dc0c100cc000c000000c0f00c001340000010300001000c00051c300d0c700440010d00000c30cc0003041000000041103030001000000400103f750101c100030300031c03003c00000000004c0c4c0034100000005440c00441c0031040101f100000c400100c0f3c003000340030c03001004343;
rom_uints[541] = 1024'h4403050010000400000c0001000043003c400414c1003c0013cc030c01104030c0005d01c010000041004c00c0004403300fc1000000700c04700c3403003430c000540400000cd0010d001c01300c001c033010c0003c00044300004540401010000000443100000000001000c0c03040000401000000340000500010f34700;
rom_uints[542] = 1024'h40010430001c0051004300c0104003c0c045004400f010f14000111004407030000000d10010000c0040305000300000cc000c0030301130100c00300000031033005c410001003030c0040100c0c100c0c0003cf4030003013740040033c3c1011100f0300007400c000100007403000000000003000040003001c50f;
rom_uints[543] = 1024'h4004000fdc00010100030030c0d0000000100010c00000000000001000000c0071001000dff30000300c0000000403000c003cc00000c431100070303104000d03000410003000100100000504c000030000000c030100300000000101000071300300000050000000000050000000000000040000c03400c0100700300040;
rom_uints[544] = 1024'hd30010003104c00c005031305710030300000400c030703c04300001fc1c000300cc0030000c000104100004304010040000c11010000c0000340044010c100030430c07003000040034000010cc3500400010f0000100004f34000100000040300000100130301000000334100000400030040c003004300030011041105;
rom_uints[545] = 1024'h430000003070011010000fc00c013c00011400110104400040440430003c113c10c14030400000000001000000c0d3f00700c000003c300c043c0001c01130000c004ddc100c7405000f0104304000303000f0040000130300004c10000f33000f4040000100000c003000300c1000c010000c000c0303c40004003c0c03040;
rom_uints[546] = 1024'hdc000000100000000040013530001300c00010007000c30003000030040103037003c003013300300000000000013100013001000000100001100030c110c40000c00000100003000c000030c300030010d340000000c00100403070d03001303003411010100100000000004300000140100000407033c1000100000000111;
rom_uints[547] = 1024'h340c0c1c0700300c350034c43010300c700c10000000040000001001000103403c0cfc00101404300fcc00037300100000040000c000370c000400333f1100cc3000304047173cd030033c140013040300011f100000000c311043c0001000000c3400000c11010c0003f100403033050000403005004c040010430000c0cd;
rom_uints[548] = 1024'h70001000403000000000c300000001000000c0013030c004c40007c100c04331300c07010000000c00000030140000c300cc000100300000c0030010000c0000007044000000540100010c00c00000000040003000010c0400000004f4c3340c10c0014030030000c00003000000040000000000c0c01434000cc040c30;
rom_uints[549] = 1024'h340404004000303000000c1c030000001000000ccc040000000100000000000c3cc0000030100004c040300000c003000c100c00000350040700c073001000000041000500c0000330000c0400000005000c000100031000030000040100003cc070430000c0000000033c00000007000000d031000c00040031c04d000033;
rom_uints[550] = 1024'h300000f0400000000000300c0000000400014000400d00c000f00000030001f0c00010004000003040004003f000000000410c10000c4c00300040030000000001004f0c40300410440c140cc41000100000004000f4000c004013003000c03000f04344300050030cc030040054100c0000000000c00011000030c14000003;
rom_uints[551] = 1024'h4000c300d51c030000c0110c00c1030c00340001010f474c0000c330000040404001030005000000c0301300000300000104000f0000033c00000c01044000000003430000700014110c00300300100000030040c0000000003010300010000070f3c1000000004033000000400100c10cc30003000300000030000000014000;
rom_uints[552] = 1024'hd10030000000010c00c00040000c000010400300000400000440040300003d3003504000000c040001c000c400000000c040cc0c04d0304013313300030503000400000403000010cc0000fcc700000403001000004030100c0430001d00003c000001001040000c030cc0003000400000010000000070c00030003000000;
rom_uints[553] = 1024'hc4c00100403c00c0c500050000400c01000004000300c00d5c00001400030700000c34404000c10034110c000c000400703c00cc5000301004001000003010c00ccc0000000400040400040f0c0c000c00003014300cc00101000c0000000c001d030100051300000043c4100c0000c00c0000c7001000010c00001014001100;
rom_uints[554] = 1024'h4c00033003c413000130010c300100030c0000300c3000000000100cc00100150000010001000000040000000000000300140000300400001100f0004034000040500f0101003c00000000c4000010c000003000000000043000430400c00400c000010000c30030000000003000030c000000001430c300000c000054c00;
rom_uints[555] = 1024'hc00333041c0c000030311d01000cc40000440003d03c4300000000000300c10005030c00400cc10000000070110330c3000000045004c0400030010c0040000000010043010130000c301c0040400f10000000000000000043014f000400700034001100f03010000004000330100040c010000000004030040040001000340f;
rom_uints[556] = 1024'hc004000c01001003030140c0010c004000c001000330000c00c300000c00d034400c04010130040013010500404001c10cc00004104cc0000001444000c0000c0400c000100044c40d00400040000000440100000000000404140f440003000047030001010d4000300c0000400400000000000003000003000000000000f0c0;
rom_uints[557] = 1024'h4333c3c110141c300000c000010d40000040000000c0fd0003c4400770d041003000007c00c4170040005003d103004043c40004010c400f40400c00300010431000003703400d003d30103001d440c01400047310000c01100c00000031400070000000300c0041c330000174c10100c01410c00407000001400010cc000300;
rom_uints[558] = 1024'hc0103000000000000c0000000100cc0cc4003300f34300030000c003011c10c030150400100c4f013000003004300030003103040000000100003030040cc040010c000c000301000c03030f3000c000700000000004c10400000000110503111301000004000d0500000c0c00000100004c0040000f0c00000010c00100;
rom_uints[559] = 1024'h3004003f00000000000000000000f000030000c000000500300000050f000045000030010c0040000013f000003400000000000303000003001000030300000004330c440407130000c000d000000000000c1000000001000000003030c00101003070000001000c0400001003004c000030000030001000070000000001430;
rom_uints[560] = 1024'hc000c000c000c0c10c150000c000010004c0c0004c000c0c7000f001100500c401000004c0c0c10000004f0001000003000300c00000000000000030c101c40040330500030010001070d00043040000040f00000400c000000030000003000000d51043040000000000000001030f000000c4000070c30040c570c003;
rom_uints[561] = 1024'h440001c0000004000c0f0401100030c330003c00004f00004000040000000d00c40030000f0c0000001004000000303340c10440cc0100000c34300400001104000000000c000c0cf400044015100000100000000004010004300cc004c00c0470c0000cc004000c00c0070400c000000c404010000040000c0c01011000000;
rom_uints[562] = 1024'h400001d00040003005f0000303000c000c0c0c0cc300c0400000300c40043c001004043704000404100000c000400001c0100000030c0410100c30000003400000404003311031701c300000100010dc00001000000013c4c0000000100001010c000004000030000c300c0030010010004040c0000d0034d0070007003;
rom_uints[563] = 1024'hc00c00000433c0000050c001400140003000004cc304000707c50330c0c0d3030000000d0700c00010300003400000030073047000c0003c0100003c03000000300dc704000000303000000cf100004300c030f0c000030000c07000c00003010001c103330000000130300043c0030000040000c0000700400000070010c;
rom_uints[564] = 1024'h4000000010100040041300c031c0330000f540000f043330000000400c0c4303c0030505001c330000f050c0cf00c0000000000010103f3000c0000005100000003004000300c0054000001300c000030d0c0cfc000000000c0004100300040f34c5c01430010033040c0c0070100000000003c00c0f0000c3000f00000c305;
rom_uints[565] = 1024'h1040000c04c0004c0000040cc0c4004000f0000000c0d103c0140044c04c3400d10000700145030000004440000dc003f073c000010000c00053c010700004304c1c0000d0d00000007010301030330001100030040000c0dcd3c004cc000c0400300f0043700d00030400000300534030000101000004001004001c00110030;
rom_uints[566] = 1024'h10c0003007047ccc010404300307104f00003c00400304000c154000000001130c0c0c3c0c140400450c4c0000040004000304100c07000001130c010c0301140c0c0c0400041f03030f3000040c000c0c40140004000004000c0444c00004140c00000c0f0c3c001331010c1c00000c000004410d0014000000300101000130;
rom_uints[567] = 1024'hd0040d00005c00000cf33f100300003000030000304d100fc03000031341100000c0001000440c000000d3000700000000301010c0101000000000000031100000c00010c400300000000cc01d3010010000301003000740000c0000111c1340cf373007010000000c130c000030000010401101010350300c0c1000c000003;
rom_uints[568] = 1024'h3000000030300010d00000c4000c10c0300000d0003c443004f00033c03004c00073003034f01730c0001004000004430000040000d000000c00000000d31000c1001c0c0030004401fc00003000000040000010001040440400414010c00000c00c00100000c0000000103000000c00c03040c000000000c04030c0;
rom_uints[569] = 1024'h4c0c0400cc003f0100000034440000c000cc000403000d004040010c0c0004cdc40010000c0cc010d40000c0c000f00000030c440010074c00000007000000000c4c0c1c3c0300c0f0c00400c01010000031040c00000000000040c04010400000003000c0003400001437000004300c004c00000100c400304c00007000000;
rom_uints[570] = 1024'hc0c4c0000cc40c0400010f00c11c440c004d04004d0c43004cc3000403030041ccc0001000040c0001014400000300c4c001c1c740400c5c40d44000000501c000c000000300004105033040030cc440400c000000c0000fc030000d000400007cc00010c110034cc0000040000d45004003030f03000f0d4c03100001010c00;
rom_uints[571] = 1024'h3000310300f000c043530c3d100000000000000300c3300000c4300040c00c3000d101304310030100000030c0150c00003400414000c001130000431073000033c0140000031c004c0100c0c04000000400030100f0cc043110000c4000100014c00c1001f4c00d0000000300010c01000010000010d0001010c00001104;
rom_uints[572] = 1024'hf0003cc0000c000010111c00010000040000000c05c0304f000c3000fc0c30000c04c0000c7c3c000015c410100400000c40000cc503f0c43040c0000010000010ccc04c0c103050000000044c0000000100000400000400c0010010c00c0000040010000000f000000c040400100011300c000c0000f000003000c0c5400040;
rom_uints[573] = 1024'h100c113c3c0d0f0010300140c030040000044c10cc000400001000c0000c00050c001c404dcc310cc00013003ccc003030f0c01c004004040fc0000000003c301000d7c03c01c00470000000cc000f000c00c00030000c01000c30c010c0033400074c00100000000544000000000000000000d01000c00004c300000c0c4103;
rom_uints[574] = 1024'h100404100c40010400c0003000c0400400300c0000001000000c000331100040310410000c1c0c10003c400510300103c0370010004000f040030000041400c031101000010030004c010030000300337c0c3c000000340c00cc3cc011001c003400c31070000030030c040400c00000151010304c0c03000010100c01003007;
rom_uints[575] = 1024'hcc105000c700c0404134c0003cf040c03c443040f30000ccc3c0c013c0c00000dc4c40300444c0c00030f000c3c1004030c0041000104000c041c40c4d00c0000330cc540000cc00304440000000c0c0300cc0041000340c040400c1400440c0544000f100040000000000000c0000040000030300c00003300440004100404;
rom_uints[576] = 1024'h1c0d47f13cfc0451373c733ccc70007cd00043113d1c3c300373033d0474001f33cdc15c310c030043cc44310f77171c314f33cc01000c03011c3cc051003d1c10d01011375040015011c3013511cd140cc0dc040cc1c03303f330c7f03130033303c05f5f517340cc00dc4041f111c037c70301f05cccc3003c304131740c7c;
rom_uints[577] = 1024'hfc0030004f400001f13c007440430cc7000c40cc0ccf70c100c033c07510c13035f3c044074010000d1701400073c000c3c3004013c44fcc001304340f1c500c10414c50c5fcc35c434010c0f4c0c340d313000f0003c000400440c040013000f434015c0f1f44000fccf333f00d3000000100c0c1c40f040d1340c0f0c10000;
rom_uints[578] = 1024'hc0003c47104000000f000c0c0f0430d40003dd0c1c030c30cf3d00007004cd3071000c503014fcc0c005d0c04000041404d00000004105f000110c0c00d47034d405cc07303000df1c00d10c71100001c4c0710354040030c1d3040c4c30f34d333cc0dcdc000000037011c13c10500004f404cc04c47c3c0300c00c007c7c1;
rom_uints[579] = 1024'h1133d3371001003f1c0003c0550fc0c100140f13034c310c001431500c001100f47703c04000d033403303cc01c4000300350374f010c130405100f00310373001f100004c3f13043300000705000430c010c0030c0c330503d304431400011003030000d000ff000304341300000001011047f3f00000cc100103c10000;
rom_uints[580] = 1024'h100005c31031103c43337010f31007700015000003c4c030dc330c710300007d301035d44c3f300040d070000110503c10114030d5f34001731440401710cf0431031300003300d5003c3010300d011033103c0300c3000433100c05c00f03010077074407c5001030c000103f41c0c01fc003017003df40f300c3000c011f0;
rom_uints[581] = 1024'h310c040fddf0004d10f3c40f04c04150c015dc00dc110013c41733400c1000405370307d0f0dc000d0700d400330d700043c0f30010f013737710f1370001f047d34f114d0f40cc50d4c0c43030c40300cc4c004c40000033037c3c3f00f030477d4cc1501453007f40f37707cdc4000cc3504075c00040700f0cc3733007710;
rom_uints[582] = 1024'hcc00117000cc400343cf114710c3031003c130304000307000000d4d3007001510003131004fd4130450c00001c00044c1301cf00033c310000000303334470c0f03330030d013c1710c00004070433000c0030cc007c0c0c1c140d0700003d10701030011314030d00330c00310f0f377c0c7cc70c7c30f340100505074007;
rom_uints[583] = 1024'hc040c0017001dc51d4040f313c0f3c0c10c001747343f0c001c7c30c150014d30150c301303cc000043c41400f0dd00000000c44400130ffcc034d175430400341c3ccc400003c33344041133347000070c0f7100000cc1c311c030ccc7000f0003010700000010cf30400500443131005c0c0c3445dcf00033c0ccf0c0f0004;
rom_uints[584] = 1024'h71003500143cd0403c01441dc1d40d4003f0400307040c00d00040471003c04110073044000f33c00d03700cc340574cc00514f00513f0300c7d0410433000f00d0033f0f0414cc3444d0cd404c74dcc3f1000d0f4c0c15dfcd3ccc4c0c40001d001dc0c4304d0c00cc004d04f00000337c4f3330c14d0010403c101c0000c3;
rom_uints[585] = 1024'h10c00c0300033cccfcc3c113454400fc043c1000c4c4033f473c0c0d133d00000c04401303050cc031043000f44031d40430d073035f04340c04100000300cc5fc0c0c3c0f0d11041c0c0c003c34c43c3000340040004c130040073d03c3c4075c050c00010300043047c00f003c000070c707300c41443d3c0c103c000dc03d;
rom_uints[586] = 1024'h400cdfc340c00c01d004c0c00003333001704033c3744c1305010d00030c1300d0000330c4c150005f3f50c0c00157000000c40000df30310073300f30c3c0404000450cd140004c003000c1cf330000c1140d04100000c35354c00003ff05000000137c7d430005f7d00f0103d0c003c3140110d014710f3dc0c1cfccccf0d;
rom_uints[587] = 1024'h310c440cf175300c100f1000c004040044f0cc00c1040413cf1013440c4cc001100030cc1041100300ccc30c4c47440100400075c03cc3000401cf00c3f1fc00fd3c0545505400f1cf000c514030c07330cc01f030000000cccf0004c000c001001c0fc0ccf30000300f00030005000000414174400435c013034304c3130cd3;
rom_uints[588] = 1024'h43033ff0c103c447030043ff010d31d3041443003c101d3001300cf3000010537c07f750311f474010c0c3340001401341000107c031130d330fc5301103314dc7045310371300040000073df3d3f300c70030040100313000c43c4d00ff300df10c34104317300dd0310031033f0000c143000337c05d0ff10c300434304003;
rom_uints[589] = 1024'hc00043c000dc30d044cc31c00c0c100d00000100004c1374f3404444c030cc130c1103dc1c4070003d0cc0cc3074700c00330cc300c00001000d03331f403d01d0c30370c04c4f00cc17001074d00300c5f00c00333f3333f0003031c30fd0001344c30100311003cccf001300710f0000c0c001d3c40c0000000031cc010071;
rom_uints[590] = 1024'h315cc473cf3371dc00ccc1c03c4513c0144d3703cfdd033cc0004300c34cdc000000c0c70dc00741f45c000c000450300c0fd33c004c3310401c0ff700f00000f3400005544007001c001003130100d030034304c30133003cf37000cd003c0c0444045d000f30fcc0043d1440c000003f0c47104ff0003005f101334d040;
rom_uints[591] = 1024'hd00010fd10cc440f1370034073747103044050004f437050f5d0c033c100110c0cf730414100170053700cc331301010c751f0f03c3140c4c0d7700074003003c0314000101303405d000cc00c00c0403fc003c4c0530003310705cc300c00c1f1f343500f407334033143430c13100070c4c4d30cc3c4c3400070c3731f0053;
rom_uints[592] = 1024'h407043dcc35d3344f3f413c7c000f00000c000f0d7c3441c30400050d431c3040d504340ff40c0fcd400003100454000cc33030c0000c107d0c0c40c1013c04c13c0034041c40c03700001001c510fcf4cc00113c0cc04c05dc0fd40c4c4f1703541c0315f03c1cfc0400c03314fccf30100015301d0340034c40010f10040;
rom_uints[593] = 1024'hc070c01c73344c0100c1c310304373f0400c0cc03131d70040c0040413c0fc0c113f43130004c0c5fc7ccd1c03d11d00033c10354040cc73c0f03fd03cf170c00c0303c40dcdf0fc1305f14010700300fd00014f34000003cc4f34f11f44c0c410c13033c0131f433401004c05310c0000f1c4413130740043c404414ccc0cf3;
rom_uints[594] = 1024'h30c034df0dc0d13c003f50000d70034c01010330510d3c0100000111005d340c0300010c130c1300701c3100dc040731370100fc00f00c3400301f0c73301c00c00c40f044305001303c040cc41d11010c040070d1110300c077c0370c1101703707040c03c0003400f3303ffc43000c443434f00c4000c0003c113010340300;
rom_uints[595] = 1024'hfc01d40f3f3f40c01d3330cf30cc0c000000300000400c170c13c044dc40040c1300fccc130c0003c43cf003301cd5000000c00c40c3f17530300cf300354330313c314117000c30c00c0000134c000c7ff0410040c001fcf0c05044c000400cd3f03fc0c04103014c3300c311430c400005005513013cc4030003343f54c014;
rom_uints[596] = 1024'h700074fd153f140311c1c0030df03530030c0c04c331030c335c1311701054f1340c31f135c0403050c344c13d3c4c030031340310370c1300c0fc470c000c040503010c4300300c3534330057c00337dc000f5c0c0c0c007330004d3030f1300130cf343f1c3c00c1003331001f033c04703744003131400ccc0310f0050f5;
rom_uints[597] = 1024'h3070440f401000301100fc0cc30c3430f4303400cf3740400310700400011d001cfc303c4f00c500dcf00070c0001004c00040000000f0f31c300d50f01440c0f100f50050c030004070400340c0f410ccf034c000f4f00dfdf11f103030c0100c003130f4345c00340ff0ff00c000c050145010401c0310dc1010c0fc010101;
rom_uints[598] = 1024'hf000c00f13c40000c33345133500fc41cc300000003c030010341070d35403f0103c333c0054400c103d3c00305310f10c4f01c743d330011031c1c04c3c4d307c0170c41331010cc30000031030f1404010c44014400001cd4cc750ccc0cc0401103330fd4c530004c4f1133c0303030333c400331000000330100d0d100c50;
rom_uints[599] = 1024'h1030107d3040f40c14000c3000ff0c43c0000c0333331000010f10f33000144f33500400f04f1000010001000400d5010c343f30007cd00c001144004c403c1f451004cff51030504c70307f3344000031013310f004cc030505f3f0003703cf0f1f371050143103ff3f00410f304030c3f4c1d334c00f100003001000305140;
rom_uints[600] = 1024'h7d0043313444c000133c5003513d01c100174400c04000d0c01f00cf0001037c13c00370037c130f033d0c03cd13133101c340470001f000434131333040f0000701d34f13100140710c07ff1ff331030100000c77cc30310107431c7530cd03107ff4304d0cc3c30c1dc3030d03c000005744dc1333400c0340030d30d3307f;
rom_uints[601] = 1024'h300073c0d1dc0300c3cc1dc0f017c411303f0c40d030c03300033340001c70c70f0703c0d4107c004cc0cdd0c0330000403003dfc1113170c7f1c01f153cc17110f3300f43713133c0d440143fcd0000c10c0004ddd3c00000001340c1103403377f14f030f03c33ccc3c01530100000134f0340cc0373031303033100400000;
rom_uints[602] = 1024'hc014f1074300f00734435000dd4cc0c100cc00005d500330c0343000330003d134010c007010c57050103300003000cc00c10110030000c000500d03045340d1040c00d337011c503c14010443070030100040cf1000031000310f43c134001004c04001110f300fc0c00c040451334300c3c303443010000c0030c0013013c0;
rom_uints[603] = 1024'h430033043001c3400ccfdc05d4034c0c007f7100f1f4443303cd031c34000370c1017070440dcf0000d30d01d0d0073000f1f5c004003c0f44c00f333070003340007f3d00c3c07371050c3c00c0440c110cc04301f00330400300c140f4013103c3c00c4f4340330c30033001cd00d100f1311c010331f0cd0303df10c04fd3;
rom_uints[604] = 1024'h470f0c3103f35c3403d7011c0d0410013c00004d3fc3c0310001000f070417101c3f101304130400d0301010c30d3003330170310000000100031f0c0004304c0d00040710114f10007330cd31c03d0001300100000000c000350c013cf13704000d341c3000310035033400003000313d0430000133033303f40413040cf;
rom_uints[605] = 1024'h3003105103c0430300f0f0040df01030d300cc3c30301041c00cc03311344300013c13d0c03430040414400001f11c0300041341401cc13010c0c40c30000000000033035030f00fdf030d3040701007700005003c30c0c3050011fcd0701dc0c0c31cf3c04001c0011cdd100070dc00000054730430c53010040044033cc04;
rom_uints[606] = 1024'h303df3171c0310d03300cf40331d300305f0dc03104571301d0000704011fc0030033400530df031c704d3547004fff0c0510f044cd000ccf4fc0103d0c34030c034c30000f307d410000f403743330300d3403010000c013ccc07137c43700ff003c7c4f43340030c003cd0071400043ccc3000000f4131c0f000ff351d00c;
rom_uints[607] = 1024'h431d040fcfcfc341050c40104c310041700050004c30c0c000300404c010c4710401001cc40d0343017f31400704c40c31c3003cc0000000c04c000401c00343415fc001c434cc0c134c43c5c5c140304c7300013300300000500f3450c40ff301700c0041c0c0143ff3000131700000c303c3c5c1f00c341030000040044100;
rom_uints[608] = 1024'h340d70cf0ccf103000cc30c3304000350000fc401c3dc7f307377070c00f00f000041ff0f34cf00f44140000003371011c3d33cf514f344100013004050d1cd000c000003370400c00013f4100dd0d031c0100400c3c450000c40f4103cc0c007430030135100344c0cf30503041103d070cc3100cc4037510000c41c100c440;
rom_uints[609] = 1024'h4300100303744010d001c70337330d1000d0c0404043500400c13133d14cd13cc040537fc150d003dc71d001c0f0c04cf043030433004103007c040c00100041000040d1ddcfc04f0cc1c040314111cdf0c30130c140c330073300c04c0007000c000c0c0140c0003f0000c001c000c004d4111c11034010003300c370cc441;
rom_uints[610] = 1024'hc0344330c30000300300c000f0c7c00001c1c00001c133011343c0f000c003437c00310330c330c403c13000c70001cc14033040104000d001c3303d005c000c400141003333c001003300573000000300c001c0000000000c400044073dc0c340333107c00040001300014040000300400100474c00030000c00003034f01c;
rom_uints[611] = 1024'hff004c1100301300303400c0d3c4cc00304c03071040c0d0300fc00cf10410cf000010ccc000cc1000df0c101003430c3000037014300014300f044034001003cc0c004c0003c703cc31000010500000100c40000f1430c0ccc53340dc00cc70c53c34300f1c00f44c0003c50f4001401170305f400c034004300443c034c3c1;
rom_uints[612] = 1024'h300004d07d1dc0c000004d0c3f3cf00d4cc0c0c43d0007030c004344137c043f17cc4fc01c7cd040c50cc0cf0047f4113c30031f00130003300d00cdf0f00c00cc00f3040417cff0f5001130143111100c0c40c00c0c030cc4c04c0cc0404c5ccf50cc3101c710030c4f1cc000f1c010704f530f1d000f00004040c0c1001d35;
rom_uints[613] = 1024'h1430c31c00540000f140044c4070c0040c0004004d3000cc00700cc00300cc040dc1c053cc3010003c013c3000cc00400040344301001031cf00103f07071100d44000300dc01440473003fc0030000001d0300000010010d0c0300000013430fc051c40040000f004c00c0c00701c0c0c4433c10cc104cc0c0000c01c00103c;
rom_uints[614] = 1024'h103700cd443c10c0000070000c4014303f3c00f17103c31c54f30300d3300400c03000d70430c4313cc04101cf03440d3050f400114c1003344c40c040401030401c43f05400310fd4010503345cc0554c40000c500f100c0c5c014330004c3070fd5c04f0031c00f0303147c14010000f700004133c30001005700010040cc;
rom_uints[615] = 1024'hc1330d1f4104300401454c04305cc741007d11014c3033fcc41307c007040017d00c3c1310070001400c010c03c40c404c40dcf00cdf00040744c300410500300100300007c4400d40003003ff0c3cc00000040c0130f000c00d0000fc0c3104c0000040104c00300cd04103014c0000cc30f730130c0401c00d0700070c304;
rom_uints[616] = 1024'hd34c3d00fc0fd00340f034457c0030001d5005355cd0340cc030030f30144334cf1c533004c4c0340cc000c0100c00430470d10f711470001430f011013001c040cc0cf014054c43d1c0303d00300130300100030004700430300040c0000703013d144c5000411303c0000130000cf00c1c0cf0d4503cc03000343cf04c0;
rom_uints[617] = 1024'hc000f44c43f140c0f1003501104000010c00370303cc004d11f4300000c144c3344c00753c03c13c345d000c3c0cc714303c00cc5303101134100c30f4f450050c140c0031c4003404cc03100f50d0017000c3d4004010f1410000c700030c0001f33000045331140f43301c01c0f04c4c0c01370f041c000401000000300100;
rom_uints[618] = 1024'hc141f50c031f3000f40f1300d0c31d110000c0430f00fc003c00044530033c1c1040330c100c1400c010314100c0343103331c0c03031154340110cf770003c051dcc00134115000f0004004000d0cfc0c0000030300400340443334c31c0c0010c0f1000100003043cc3000c033000400303004f0011300f100f00503073134;
rom_uints[619] = 1024'h31003075344130131001133f10c07d17340df00507343c10c440c040300cc04c4c140035400c141c131cf0050133000305c004400d70c7c307301c000400030c0014104c0f00c030304100410003003000c047003003100c3cf443400504770f1041c4cf073133000070100f41000100343437014fc703110704400d1d0010c;
rom_uints[620] = 1024'hc1007c03c0140030cf044405c40d0c00003c3d00c4c133c310c340000c4303004f00003d03330313c440150340030c411030000400000d1ccc31030000cdd4040457c10c500000313d4c40c3031411c0100400010500010340000010430700005340010d71015f0c003000d04cc40030000300d0030f1c0303000005174f5000;
rom_uints[621] = 1024'hc30000000115100010cd0100003c330d03c0cf30c5003f0c0f150f4434000004037100c3c00510c101015d04111fc003400400040cc0cf0cc0ccdc4130c00cf05403000400000c03ff34d0707144400c000c007314c14cc100cf04003c05c5c070c07c0cf3004c0004040030304100d001d4c000010305004cf0010c4d410000;
rom_uints[622] = 1024'h3300004307c00300130d31c4c033003c030c0401f33104030000c01c040c13701300000504fc0f01c33c0400f0c0d300c340000d0314000c000df007430003030001000d530c000304034003000f4f000c0003100c0fd00700100003040c310104cd400d000147030c10001700030c300cfdc1cc0001f003433d010f4f100010;
rom_uints[623] = 1024'hc0000440c04f30c0f10c31405cc3c03003f00c0c0001004030003f0140033c05000f34014f013103c00ff0000cf00c000071003307cc00d33d1c030fcfc44000330ff300f0d00300010c00d00330c03f00f00300304f1d0fcc0400c30030400504003c00130c430045304000033003f0440433f13ccc100303f14004400003f;
rom_uints[624] = 1024'h5c074ccffc7330000cff0cc013f30c34c104c00f00cd34f0300403410c005c10410c35d300c453044dd003cc173140113c000f3033004530111073000043331d4f000007715c5001cdc04033fcf0433300000143300c300d03433301cf00c03d7013f10111c00000ccc015010f3003033c30000c30503000ff33330cd30004c;
rom_uints[625] = 1024'h3340031c1437dd334030f000c070041d003cf30c01c50c0dc400c01003cd00000d7013003304cc0c03d1074003033c1334c313571c4000c530c3003d7433d10c14d00450000300c40f73c0401d111000c1c0474000300401f43004c33050003377c3000fff1d5c3c404033774000003c0007031c0000440d003c0cd0ddf0f100;
rom_uints[626] = 1024'h4f00340040cd0010030c711c1c0d3030011740c0c0c310f00cc40034107104ccc30c0013c4f0300f404f700c70041470113000fd10c1733310307c01fcc04c1c70c040c4f413301cd3d030c0340070044031f050703000fc407dc000003cc1c1ccd11c301357d100c1f440c0c00104f0c0010044c40ccd30000340330c071d34;
rom_uints[627] = 1024'hdcc0130133cc3cc0c004100c0140011c03f1000030f70310341400cc3405f010401ff0c0033314043c5cf00004707c3d400140c17000d110fc1100cd30300c5d0330fcf3700030f000c0d4030cfc00cccc40cc7c3004001c0017377000c0d30410cc0dc11cf4007c00f00450cc03003747f3f031f07030140303001c5431133;
rom_uints[628] = 1024'h33dcd1040043000030fc030d53f5004f10c005f0433300300f0011fc040030f00c1f0cf1370005c3d500047f13dd0c3100033c5004f3030c00110c00d003c0070040c4f0f04d5c00003c00fc1f0cf1d041004c00c004cfd1007d03000740f347110d1f5300f04010301140c10030f0f44730c100303000300030310540c4;
rom_uints[629] = 1024'h70444301f013fc403c10140034c04c54c03f00f30d770030d014c0701130c0030c333c50007513311c00000000d1c003f044050300f140d3037304d0304f00434013433fc13073000070d0304d00331040c333fc0030c310c3d3c1d13c0071c0c010d0304f7f11c000cc000000d00300fc14d05d010c07134c01cd00cc0010c0;
rom_uints[630] = 1024'hc0c013014f100c333003040300030f0c00f00f0c4314013d0c00c400011331071c0c000f3057c530350f300340170103005c00004d0330000503300d03040d00cc0cc0103107d3003f331070000d0c7c31000000104303050c0c10140c00401031000f3f0f0d0c00403d033c00140f0f4c170305010d040d000d40010001f000;
rom_uints[631] = 1024'h405331d3304cc400113070334030f00400c430000414d1100c3033143d3500403c10d5030c0470fc33d35000c03110700034314cd0c074300047333c44001000000004311d454043330040cf00d7000010000000013400400000c00c00d0c03cccf177347310d0c004f0101c0000dc10c03000151c0071cf0000c00000005c04;
rom_uints[632] = 1024'h10dc33407100001c003400c070000700d030c0010513dc000c003030701000c0f0c0330070f30001c70403000110013004c0140003101c0000370f00013000f4c300ccc10000343000400000040030340400c044045003340f0041ff570101dc1d3054030010130f0c0000100100340011001010001310000043c4c33c0301;
rom_uints[633] = 1024'hf7cc0f000dc40c401007c003c007343000ccfc00330500100414500103c4d07f107c0c3f03ccd0000340000d03000c3d401c0fd0010f0074000d330f40c301003cc5000ddcc0340cff0cc0701c01300041c00c00cd0000cc0f03040d330107c447c0033cff0d0000cdc40c70c03d00311cc4d40140040f50130510050301c300;
rom_uints[634] = 1024'hd03000c70d74ccc401003d3c003c043d033c151c0d5043d00f000300330c104400331f0730410c34010dd504f0cf0c573c010077c344041f0c57cc30c7010000c413c170fd1c00711504000f401017c0c00300031000034cd0cf4c3d000c037cc300f411155c330f400400c000cd100c50334000341c437130030001ccf03c01;
rom_uints[635] = 1024'h4c3000d704410f300c04750010c40034003c03cf0df0113f0cc43c0000000c11c0034d13f7357d00f0d04f07f4dc01701330c770c013003c0c007730330f040107437f4d4f0c034cf4000003014c701c014c030c4030000dc347dc03c7c3400003014304011c1c0c41df00030d340430c34c7c0d000d010134cd010114000d05;
rom_uints[636] = 1024'h5d4031c31c30c143511000d0c334f00074300f100030c3f07c30003c3f33ddf1053c05005ccc5114d5c01010f4073000700d0cf00cf0330350303c344310d101c0304c33d3341034010c047c30c03c0cc7c0f30c03000000c433d3000d00430010d1c0d07030fc0c3c10c43110c000037c3c0301030c00000f0cc4d5001170;
rom_uints[637] = 1024'h1000c0710c103c0c17000d41c10454fc0c144000c0130430000000034cfc00050d000f4501c10d0cc3c00340c3f0d00000c04107004c4404c310003c3fd30cc1100017c44f10c01440031433f30fcfc03c00100304000031000003c040031c00f0001c07150301000417c0c00c3c03c3051450c300cc15f000c300003d000503;
rom_uints[638] = 1024'h307457cc07fc1f500f0fc0c33d04070ccc10d0f00030100dc3711d0cd000373314003004d040d0010fc44400010c143c0cf3173130cc0d000034cdc04c100c345d3c5f7010500d30d405344104fc7404fc130100303c1cc41dcc0c041c3ccc04c30dc1330035dd1f73f00454010c30300c300074f00c7000cd400c3cd1d3c00;
rom_uints[639] = 1024'hf05d35d4f050c0100703f5fc01400030c50f30fc00034011000010c0d00033cf0045f1ccf71c00cc300033070010403030f4cc11054f50ccc430dc000d00c713340d340003c331ff340c00400c0403f010f014cc40c003c71000c040011c0310143511300010003d4f3040304000400410034003c00003000c0c3303c04c1;
rom_uints[640] = 1024'h1c4007f13cff0c05000c333dcc7c0c7c100c50000c1dc070033350043041040c3701c55c010c430043cd44300c07c050010c3fcc01401f0000507f35404d3d1c01c310c1371c0c0d0c41403135000f07cc370c30cc0dc3f04f373c30c101400f3307005c13113000cdcc0d711030013500070711311c0c0034707c0cf1473340;
rom_uints[641] = 1024'h3100c0c40f050c010c300f3700734cc3c01c4c000ccf04f00003031774131030f403d047c100c10000030d000003000c00cc7401100000c0c05f30c1cc1c100c00414c5cc503004c407c01c0c40c13701000100300cfd0c040c044cc70053300f037310f331c05000fccc000030d14dc00f105dc01c40fc40d030303f0d030c0;
rom_uints[642] = 1024'h15443c7000400110cc000cc04c0400d004c0dd3c1cc04c303c3c000c7044fd3031440c503010c0f0d005c0047400001c00cc414c0c4000f400110f4c30d044040004cc13f4000cdf1c00cc3c700040c104f040304c40000404cf07c00000034d3c3cd1dc0cd0c03003700dcd3c10101434c433c034007c300000000c00004cc;
rom_uints[643] = 1024'h711731334030004ff4c03300f410f100000541f1f0300301c1113705c010401101473700040c0113f0003031c0014000340f50370001c11f0735d10c0431334300105c00030034704301000c3043037f10304c0000c0d3341030c07030000401300034000d400f074030035dc00000011f10034000c1000cc03000f3143c3;
rom_uints[644] = 1024'h4004cc3033d030030371001315037000c033037ff4d000dc30507507410431035005110c40330f401044000c001000c0c5400300c353014304404013c4c3c001c31f3111c010c500303000330c0017331033300c001404301c1f05d3034f00407317574301000334f100403f71dc0c0cf00330300fd343030c0f041074f34;
rom_uints[645] = 1024'h3dc0440fc100f00c0cc3c003c4c07c07c00400c1d0110d03c01434434fc0174c4f77307dc04dc410d0040d000337034004fc033130cc05c4077100d37000d3047d0001100c0007c00c4cc14f030d03004cf0c0c7c0c0d003f134c0d0303fd0c430070c01710003c3f000347c4fd00c10cf0404044f0404144f00c0043fc374cc;
rom_uints[646] = 1024'hccc0c10404cd30c33700cd10014c00f10c3f030334300c00431004c4177403c1100f17d70011cc0c3041c01004404c004c03010c4340fc7c033c004c4033030fcc0c03005f010d3014c0c00f04c0d400d03d330000144c0d300c004f00c30c7c1d70d0f0cd0714030d3c0c53c0341333037c0d31c0c03c303040100004000334;
rom_uints[647] = 1024'hd140c0414f35c0500404c00d003f0fc310d40c03430330000137034f3500d1040c5750014c3cc30c070c440000cc0010130fc0450c311ccfcc0f0c04d0c34c0f51d31c070d0c0303c10005430f40100043cc041430030c0d31dc300f1d304c3347f04000d103110033344340000f000330000103000d0ff3003f0c03133f0c04;
rom_uints[648] = 1024'h700074c004401040cc0174dc00d00d74c303400007074c03c0c00007c1030140d003030c003c34df7dcf300c030c0770c3010734141040037c7dccd0033f113c0c1cf333010c1cc3540c00d4d70040f03c0000c000ccc1410dc7c004c3d7000d10310c4d730013d03fc1041071c010f0c7c3f7700c000000c003c0411c01400;
rom_uints[649] = 1024'h471c0d03df4330ccf1c330c37407043d043cd0c0c4c713cc570c0101173c30405c0501134f053cc43d040c00044f01d43404107fc31304f43c15000000313004c3433f7c0c040135d000ccc010c303703c3143304c044400c040130c4c00c40450050c0511c303347347c01000fd003031f747f13c414531300c00310c0c04f1;
rom_uints[650] = 1024'h1414d1ff304c3030c00000010c00f0c3001435043c340701044c130ccd000003cdf000f00c7f01c005f3c1030c54c430500c0c40f03d30c31034301c37003c043004005031000004f104c10f0cc000043c5553004034040c01f5404c000cf15c0c10f007c314cc005f40c3f04f0d3c0c0c304010cc11431030103cd0ffcc34dc;
rom_uints[651] = 1024'hf10044cc0c703f30000f10c000c130000430fc000d340013c3501340cc100300430f00fc104d134317cfc70c0c443441010011750f3cf304000dc3fcc3c00c0001fff405514441c1ff400c0447cc0100c30045300000f000f3f30044f0000141031333c3ccf34300011000c34014c00000454144401045030f030040cf570cc0;
rom_uints[652] = 1024'h3173331c033c1c30f3f7f33510d310f401053003313dcf0010cc0c03cd300407c00f71041cc470054c013051cf10c0341003dd7fcf1100c33c34030001001401704101cf70c40141c00073df3d33710c73410001000010d00343c0c01cc300c7d0f071353103c0dd17dd73ccc3300c0c54300d3f3f05d00f53c30c474400003;
rom_uints[653] = 1024'hc03007cc00d03f1c04c10cc03c30004d003c0c400051dc34c3504074d3303c1fc00c430c03007000030d30c04074c70330f303c40dd03300045c0c070c433d300cc03040040041330c10131034000700013300c430030000300c3435dc0314001c45030c0c3cdc00010f30dc003030010310c005dcc40000c0304031fc004030;
rom_uints[654] = 1024'h3140c333c00070c0c1f1c1f03045d043007077000f010330f0000c00f34dd14c03c1cf0401000751f35c03cd000410300d0fdf3c744d331540c00cf740f0c00ff00c0370050404401c300030030000d33c00c30400313c0030f37030c00cfc00c4444110014330ff10c00c154003000c3c0003131cf0100005c101c04cc30;
rom_uints[655] = 1024'hd003d03d30fc70300000133033404143007c41045c414010f5d3c00fc110100c3cc73c41300c13005333cc007c040cd3c45100f00c715034ccd04010440c3003d73143400f0004415d30cfd00c01df70ffc000c0c043c400400740fc703f00c0f4c300d00c5c7337f0010304cdd3311340c4c01011c4f40300c040c0730fc053;
rom_uints[656] = 1024'h10400503cd03103044f3c340d7d1c0c44d003c04c0d0d045113300050cc041c33c0c500f7cf044c001100c000041c04c00d0001f0cc0c00103d0c5000040dcc04c131fc04000c1cc0c73000104535053c31cc00c1c1cc100cd51c1c05c10c4c071344ccf301f41c1c300100100010001c000c35743c4dc04c303d0541cf00d40;
rom_uints[657] = 1024'hc05c30c44000c0c0f30f00430cf000c1004f4005c50f4cc0040517c40c00007f00100047c0000d7fcd0c3f0100340c0c104140033f7cc0300300700040003f034cc30dc1404cd344c14503003001fc000d030470c003cc4f0001c3440c0543c17c30ccc1004004410c4c400c0c410001c431000135c34004373040cf03c0;
rom_uints[658] = 1024'h3cc0341f3c0001ff00031cc0d07000500171303001fd0c100000311503414710c7000d1c030dc30073dc40131f310031330dc33c5c3000017000130070301030c00c713040041330013fc40014cc41000d043030c0114040004701330c1c1c300333c30c4300c73100ff103300300111003100c5133500c0050700001c373304;
rom_uints[659] = 1024'hd30140fcc3cd000343fc00f30cc3000000130000c4113070c10c504d040040c171c000c00303470c430c10030130000000fd30c403f010004753f070dc143403c3cf14417000031c30cc0000f0000007fc410d000001003c0c003040c047000cc303f31f04403004d1300cc000313471000004543050d0033403c303f043cc4;
rom_uints[660] = 1024'hc0075f105fc34000435c13c0c00f50003400f00cf01031c3010430d301f44c1300350fd31c0100f50c0c0f1fc000c00000135000d03030310c0f040c30c0004c4c3004f70000fcdc534c71040d000c7cc000c41130c4000030c4c00303cf000713f33003f113f00c0040030030cc01c0775375400d070733c0c3010f001fc1;
rom_uints[661] = 1024'h3171510c0000007070f0fd4cf00cc001f0c400303034401c031c30444f31540c5ff0303c00c0c10010f03143fc401004c0000c41001cf4c410f03d5030d3000031f0f1335001fcc043400003303c30000df1010300f03001003510d44304d0100c1001f030305c13c043f03300000c0450154010431cc01c14d010c031003041;
rom_uints[662] = 1024'h3000c00f07c5700cc3f0551f0155fc010030300040700f04040550401354c330dc30300cc0040033443130300013c03c100001c400d33005043d0114100c0101300130c0c001300c0f007304100030433000c401d40070010d35d350fc303cc4c41cf37c3d3c0f0004c430030103034303c0c4300300050013000071c050010c;
rom_uints[663] = 1024'h5100d47000700441000c40334c0f00443010400033c310340103c1f77100d44c334104510043d400000301701000c0c01f703f010c30d000001030c070303013450110d33510104d4c00300333f000303101033000040000010030f00c0400cf00d3311c10100004ffff007003f33034f3c100d30430c3107403000430301000;
rom_uints[664] = 1024'h4053313004c30c033001304330f1c103104000f0400cc4300353cc0000037d03fc3c3c033c07035f31ff33f01710314000404700310104107105033c00f000f431034f131304407d0d07cf03f0f103f00700d073f0000530d707107130f0001c4cf7304d0f00333c0cc0030c03ccc0305737dc03d3544fd30c031030cc7143;
rom_uints[665] = 1024'hf10c73d100dc3000f00c0dc03310305d04330c001030c333cc030300d05c70c44f470cc100107c044fc000100c73c330044c03ccc1c53c700030c0001400c170dcf03303404c3f03dc140c1430c10c00c14c0c041c10040d00001040c10cf503377c003030f33c0301070014c000c1001343037000400300d3001330f000310c;
rom_uints[666] = 1024'hd00431000300000430571100dd5cc00100c000505157703c0f0030003304f3d131010f0f0010010040d13000403000cc50c00110c000c0c00311013004534c1014cc000033001d5000140004000303311c00000c1300330130c00f5000c4141000c041401133f10c00c0000005503003300300f3770c1000300000ccc03413f0;
rom_uints[667] = 1024'h301000c430753c400cdcdc04173040cc404f3c3001f7440307c500df74c00330d000707334fdcfc0f4d30150dcd00300733105c14000400f73004300407cd4cf105340f004c3103c71050030c001151c11c00003c1300003431301c140c030f0001cc03c43430033013400340d0d14d00cc0300c743330c031003ccc10c00c00;
rom_uints[668] = 1024'h130440c0c0100f040030fc0040cc00310003c0000310cc000f0c000300cf330c710403c40030400300000304c133301000300117c310000100d4c0f1f4c00041070401d000400300cd04000300041103130c1000500000001030cf400007c01f054d00d001c30003100350c001000303034310430403104003c300000130013c;
rom_uints[669] = 1024'h4fc4500700000000f0f0c50df01030000ccc0d3070144100ccc470d03443330d3010d003f0000d74c7003000fccc13cc03c3414cd00d3010c1000cfc34400407d003044ccdf0031c140d3030701047410000c4c00100c431c0cdc0d1c11dcdc0c310cfc4004103c0000d0301000470c0c04443443df0411c00c404003cd04;
rom_uints[670] = 1024'h3001f0431f43d0d1c30c0f40301004d0c1f0d00350457d000d3303400cd1f30130043004470d3035d300d0504303c3f0c7107f0010c43000f4cc014004f077f0c034000013c304c513001013330000c3c0c3500013401000ccd0470040433c0c3030d404353310f03d3003d007c300504f3c340000f341f0000050c3043d11c;
rom_uints[671] = 1024'h700004fcc34f1351004004007cf10c05000010113c30c4c30f30c430c704d37c444d01dc047c0300053f300003c704137103704cdfdc1f143140c00401f00370515f0030c440400c1301733104ff00034d3300c0033004004053c33410c103f30174001c40c0c0d03cf0001d414400c0030303f5f13c3c3410370300403411c4;
rom_uints[672] = 1024'hf00c70c00fcff33c44c00403c374003110d03c400d0dc7000333414033cc403030511cc0033c300c75144101c04f0031001d30cf100f054504013304011d130300d004c00000f100f0013f411c10010c1d0000001330043733341f5c340f0c3070770f0131133f40d0cf1c4000501c1c000c330d0c30033510001c41d0703340;
rom_uints[673] = 1024'h3311c3303474001103cf3c3473370d040dfc0013443405400d031f31040d13cd1044773c000d303dc751c0030f4047cc07fc0c433714404007cc01c0000cc013004031cd0c000434c00c000703100fd0410000cc1440000033700c04cc00700ccf0c0400544c4003f0000c000c00d031414dd111107400f000c010f70cc041;
rom_uints[674] = 1024'hcc33033d4f400030dc0c3c0001c30c0001c00100f1d70301000003050c00034340c4f50001330001030170300400c1c107030c5c0441c0d001df0040410c000000010003000c000130303504003400030c0000010500d00000000000000100c700030d000101410c0700c00343340300411c07034f0003004cc00303003f010;
rom_uints[675] = 1024'hcf107f00000cc30dcf0404c010f40c04001c3c031c07c010f000c31031070ccf00000cfc304fc3005013410000f3033c3030007007030007cf33c04034301003cccc004c300300000c310001c310000c003c70030f10c1040cf4404ccd00c00034300504031c00f04c3014f51f00105340700c5c40c0044d10000150d000c000;
rom_uints[676] = 1024'h3cc00700315c00c0503f710f3f3dc03d000301f43d0017140cc703441440c43317cc03c4037dd441f5f3c10000044ccccc304c1cf01c00330f0d400003c00c40c00fc4040403cff0c504d03c340000100ccc0c0fcc04330103cc4c0dc3004c1ccf5ccc3dc4c700031c5f01c1c3fd00007c4f1f0000500c0c04404cc0f1310131;
rom_uints[677] = 1024'h5304c00000540100317015001040c00000000400414443fc4c00c10140450f131ccc00535000d0c000c0303301c04000004100000000000c00f3103040370500104370f0fc3000100030100cf103f00004c400cc004dc010d01c700100410030cc000307004310cc77403c3c00000c3d00450031301010300040c10010c003c0;
rom_uints[678] = 1024'h300c7041d403c10c031c033c0cd1c0430033010f401cff00f10f000f0df0c0734c10310d01430340170d440003c00040d4040f531110f101330503041004000000c1c00fc5400314f14010500c41000144d53300d400f430c7c10014f30004c3403f11007c0d01c0133f04507c140504c0d0c30c400303101001037101000000;
rom_uints[679] = 1024'h430030ddc51000000f0c45f0cc05cc450030c100d5370f3cc31c3000d040400d7c00c3c10c007c035401d50000f3c4c440044cc3c0dd307f030c40010040104700000c030c4053c4d5c0100003c4c7c034000430c4c0404c7c43c00400dc03037c40c4040030cc43c0cc03d4001500040c0f0f770043cf401c730c4300000004;
rom_uints[680] = 1024'hdc30c3d73c003033074f03400400131000d4000357cd0040000d00f407c044375cc00500cc4f0c0040c0003c0c40c0000c743dd0c4d0440001434301c7d3001034c0c103005f17d4c13c00c300c03013000110300c10403c40030304cf30007030171154d03005000000003113c01f0f3131d0ff3c413000c30000330300c0;
rom_uints[681] = 1024'hd00cf7404330f0033c00c0c5031040c00c044400ffc3000d11f0300030010700f40c037030c00100355000000f00044400f0f0cc503313d004100c30c00450110c100c0c3005000374f000d13c7cd0014001c0300c1010f0410c00c400330c10c1300000035334d41f3300c0c03c401001c00c047f41d30004000c000134c030;
rom_uints[682] = 1024'hcd41f40c43103c01071c133c3c0300540c0cf31f7f0df300000407553403301c1440f0cc030c14fcf410c14c400404fd70331f0000f0f05434c1103040040c1c41d0f10030003000ff0c003000fc0df000000003003c0310140333c0cf10000051c5c000d13030301ccc007c10347370003104c5c0040004f0043c1403045034;
rom_uints[683] = 1024'h30050c1413571cc101410d73004f071100711f301073030130043c1403010004c7044c030700cd7401310f3001cf000340000444035000400340010130400430c0000134d000d01fd30413300d00fd0c000c4010030000c1c3d343c004404740f504d04031731304405401d304d0c31007434331040c7331007c433dc1cc3110;
rom_uints[684] = 1024'h31c7400310040c30cc00330404c1004010f0fd00c4ddf0031c304c033c0000030310003d03303317304451004c1303c1c10003050041411c300d0f03c0c11404405001fc000000c1fd300010131741c014401311051403034c00131730031100034404017d0c400c00034410401414d3000300131f00d0001000c040070f4400;
rom_uints[685] = 1024'hc304400000c5033013c101000c00c34d0003c030c5f3ff404f40000400100c30534000cf0005000c014c0044014c10c00000c1c400c1cf0c0113cd0140c3c00040cf000403000000ff040040407440000410004005400c0d0f1cc0000f04ccc501c0000fcf034f0005c40040c77000d030c4c040045004413001c0000c004001;
rom_uints[686] = 1024'h7000010300f103034f0d3c00cc00343cc0103400f33d0113010c00101430133cd0cc000510f000311330000400d030011300033c0704000d0701f4c300014330c0043d0117000c0334004013000013010c113313c0300003c0100047c0330101d301400d00400300cd1cc00703400000cc4d015c0701fc0cc00130cccf00c30f;
rom_uints[687] = 1024'hcf001040cc04f7cc0c40041414c130c000f0f0fc04f0100000000300543333d450c0f30044c000003c14ffc07003c0cc00041503c04cccc0f0ccc100fcfc44cdc304ff300f1c10f00000070c03d00cccc30340cc400400c03cc0400c0017c050404c0fccc1c013c00450340010000433340f033f0330d500043f04c004000d0f;
rom_uints[688] = 1024'h50c47cf3fc0030c07cff300100f00d000143c10f0c3dc30000d007400f405313550c01d010c010134c00c0c3003c05114c000f0033c3010051104331c00303010dc030c071511030c1cc44c0f0f04300ff0c01033000cc01404f3341cf30c3c0030331011104014cc30005c103f333703330304f30503f373c00c04f173030f;
rom_uints[689] = 1024'h3700331d0434d33370f3f400d073300c0035f3c0c01100011430f01073d100303c45d3300333c00037dd0300c003700304ff33171d00cfd43003cc004737111cc4d5c44070000004ff7000571c1013d0d1d340431011400c30c050f000110033773fd3c3ff1d1000104c10770c0001110034001d3004444c00cc0dd0dd30f003;
rom_uints[690] = 1024'h400034c140c10010000d3cdd5d3c703c00104fc000c013f001c50c34c03c14ccd7305c13d4f07100004c70f04034c4740031c1fd400d707c100c7d0030004c0c7cc070d73750701c13c331c00100700071710c007030403d7170c1dc5030c1c1fc10cc400f13d4001df05cccc030303400010440c40cc100300400400c070007;
rom_uints[691] = 1024'h3d3c7d13100cc33c701051030004010d030f10c0c7cf7300c73330cc030f030d44c1ff00300f013c13d50c0cd47430fd141045cfd740010000cc110010c0d035cc000f034303c4c3030c3000ffcfc040cdc4000003c304140c11034430100000c40d14d1cddf74000373c1500c000fdf747f3c030f40000540334001c5400100;
rom_uints[692] = 1024'h3004400510100040031301f4c0d53f50000100041c073330035cc0350f440330ff00010033cf40405c0c030c533001c10c10c00c05403f300dcc011fc1d0007c0030440140301015c3014cc0c001000cdd00030400ccc00f301400100c000400343d11c4013f4334010000c0f0100c0f00430300c003c00000004303c300307;
rom_uints[693] = 1024'h4f404c3001000040031417c004d44c57000f000ccf03300cc3000c4dc434f0030d3c3c4c01440000d00c47000000c03d3047d00300c543dffc7c07c074500113435f4f3300cd0040404000344c40cc1000d430fc0070d00030d4d4103c0040c4c1c1d00f4c7c01f040c1cc00401fc0003c07034d00c003c30701c50ccc11dc33;
rom_uints[694] = 1024'hf0c00053101cc0330304c000030f03403c003054150d300c05c005c04c0dc4c00c01c3005034000403043c0300304f0053c00c00000f30044033010c001d30003c301d010400300c3010000040000041001c0c015004c0c0701c44cc0d3300fc34004330410330101c0000d00040500c1710110d01c4000f0000050003034c;
rom_uints[695] = 1024'h4040011f3401f300103c401c0334c000000400047414c4003f0c3c003d401000dd130403cc34500000c70100304100c030330d40c3cc03030c34000c40000054140c040101050c40c3004003c0030004147000313404004001403071c00c40700c3d00474017d30031c404030030d0d4c17141110c0040c0000c30c013011034;
rom_uints[696] = 1024'h40c1d334030ccc400470410030000070100000001000ccc007c100f014410003303cc33cc70340100f70404345d13013070334400fc1700c014071303c1333cc7c0000c010000f03c07000c0c31c003c4140303400410c307cc4111f00311101f11c150c300031cc30c000013f1010400510011c0405013401000c4f330c30c;
rom_uints[697] = 1024'h30c0df30ccc00f701c04c703cc0030fc403cf30040310cd004d45c0503d0100f00703f33030cdfc41c31007c00000030400303c001000030000dc31c400c0d013c04c0ccd0c0000c3f0ccc401cc430000d000d00dc4c0000cc7304013301c4c007c7000cff4d0340c104004300000c011fc4c0114cd4000013c4c1c0000030dc;
rom_uints[698] = 1024'h4c004034c3403f400030d4c300c17c1001cc50c0d400310030c03004000d14510c0130330710c370d1cc4c4f0ffc054000c0c740304105fc014cc0cc0007050c410c140c0c000c004040000430444000c0c10cc00000c40c0fc4c4d003c0340c370c5101110330340070cf7040d004c0074300100dc430d30303c000fc10c31;
rom_uints[699] = 1024'h4c317d13044d0c00310035031cd40004007c000c0c3c13c003f00d00d3470c01c0034c1007757d007010000704cc3344c000c441141040000d0d3700337dc40d37437d410f3c0331c704c0031300300c004003307100c0c3c447dc0003f3030003314317310cdf0c01dc0c0751341300037c4c3d000d3d0d030d10011100f505;
rom_uints[700] = 1024'hc04c70f110cdf301401c7c0cd00731d0f4c3000c1000c000f74d3340300c30113145f000001c1c101714c44050f3c433cc33110cf0003707f450c040740300d401f0030cfcd0141030410c053d00033ccdf30cfcc30000f0c0c40310c00cc30005dc0007103030f34cf010457110f430033f3cc04dc0c34430000f00d0401073;
rom_uints[701] = 1024'h1030003d0fd0300010c4c14cc134040d03070c00c01f000000303f4300cc00017c0c000030c335d30fc5c34007301c0300c001d0330d440000c3000c03073300003707070f0001c0700301cc3c301f043c1010101030040100011003401fc01400130c43017300003014c0c000cf0003311010c30f301500310f00033d00f403;
rom_uints[702] = 1024'h10004550007f1005000f3c0c03c31170c00000000c0340c0cc0401100d30c0437d44c0034c300d0305c050010c11100704f0c173004cc0c010c70c1f04c10cc001d010304100050f4d7410440000d0007fd1000033f3dd0001dcfc0d0103c0f374c01003040441c0c33fc345700000403c4000074330f70011c300c0cc0d3cc4;
rom_uints[703] = 1024'h404001d30040cd3c0d00730c50001400030d40c00ff0050430d0c1c01c0dc4c3333c1cc313d3743031c03300c015011100c0107f0dd45035110040403d3c00307c7000cc01000030d3303cf1c00010400f31100040c031033c7100cc140710c40004731017cc31000cd4307dc3000001004070c0730dc00000000400333c0001;
rom_uints[704] = 1024'h1c0003c4400000000c4c000c0130010cc1010c003c5c0c30cc4000400440100cf400d11c4040430330cc030000040010000c304000044000301ccc0143c00130d0c0c40004400c0d004000f30503c000000000030301003010300007c1004500f430001c00100000cc40cd30000004000000431400000dc0003c040101470000;
rom_uints[705] = 1024'h34c0004030000000033403730c00035c000030003000001307004414101f040301000c13110001c00100003410c0030107c130040000000000000f4d04c000014d0c7000004c4003050330010003000400100000000000300400003100000403010c1f0c30000300c3000301100d400100133040d00400000000c4030000;
rom_uints[706] = 1024'h44000004001000cc0c3001cc0004000c0003010030c0c0000c011030030c400000000c001410013f4cc05c000040003000050003c0070c000c050c10000c00004c005c100c00003c01304d001000001c404100c014c30000410d004004040c00c0c00000c00013000004040000000000404c003c0041c4000003330001000000;
rom_uints[707] = 1024'h103c400404000c00003400340001103100301005c1003003000c4c3001c0000c300c0310103400c1000000040c40000000300000001f0c00001000000030040000004c00400040310c003f010300c00007400304000000000400c00000f0000f00000c00000d4c033c110c0004010d000c000c000303f0000c30f0310c04003;
rom_uints[708] = 1024'hc1004000000000000041400310c140c400000000c1100003030005144000314000400dcc4c0003000000004c000000f0100000030003040c0000431000030030043000c30044c5000030004000000440000403004000c4000000c00c00301000401004000100000003c00033010f0c0000000140030000400000000001300;
rom_uints[709] = 1024'hc014003000430400010000014c40c0000110404001c0100d003030300000000077001000000c00004c07d000704000000300340c13000d0004cc00401051014310001000000001000710040030010000cc00000000c00c0c103c000cd03100000140000400001000103003440000c00001000104100000003040400c7000000;
rom_uints[710] = 1024'hc0cc0304000dc000003000100c0000c3033f00300030d0034003000010343300000010103000cd00300130070503000003105c0c015df031400000000030000101003003074c0c03141001c0440cc400c04100cdc100000c01710000c0014100000c0030c04000010cf33000003314340040014000004c000000000044003001;
rom_uints[711] = 1024'h1400031000100400400000c00000000104000031033303001370344c10100000c000000000c000040001103300000d40040000400c00000000430000040510001d00073c000003000400043000300c0011004000003000001c030501001003000000000003511103334c310050301030100000031003300000000031c030c44;
rom_uints[712] = 1024'h3010000000f04400401001400c4004404c00004c4030000c300000000100040c00304000001040c4d10043003c0c04030c50000040c40000c400000000000100000003f1001c0f34000000000000000000000040001300000c3c0000404000100010070730010cc3300101000c007000000c0000c00000410040c10c0001c0;
rom_uints[713] = 1024'h73141c30300030000cc0040000000000c400001000003034301040113013001100030100034310001403000030000000004103003100001403100000034c300ff0f0030000001000000001000000433cc04000003004400c040c300003cc00040057c40014003004403000300c0133000c004010f0144041c40000000040f01;
rom_uints[714] = 1024'h404100c335cc00440000c0f0c00053f0004000003400000045000100c0c10031c041001031f010000c10000000000030d000050c501000500003010304000000400040000000000c0000000000000000000000c403000cd00310000c003015000300000000404014050000400000000000c1c1000415010f10c000000000003;
rom_uints[715] = 1024'hf10c000c0c440c0000000030000100d0300500fc0c000310035d00070000c330c0c000cc001dc000000c07000030005100400001004cc30400000303ccf0000003c0f001034000000c00c300040000003330410040004000c3074004c0000c40000703c00ccc0030410030000100c000004100404014410000000c00ccc30000;
rom_uints[716] = 1024'h440330340003103003003f0cc00c014030100013300c3000003f00330cc0000c3001070403ff030030d00305cf0c000010c070000d01140c0c00030000003350040014c30303044100c0000d030130030040000000c0010103050c0f0103050c3100731007d00c00cc01c0010f3f13030400000cc0c10c0011d3010030330000;
rom_uints[717] = 1024'hc000040c0301c000c40c000300000c0c00400c0000000300f01000040400010f04000c0c00033000c030f00000040030000000100000300003010c0c430000003cfc33001100000343130010040030000031030300030030003c00010c130000130100014c000000c000300303010030030404c000c40000000010000c003004;
rom_uints[718] = 1024'h3000000000c0c0c34000c000c000003000000000400030000030000000000001000000000331000005c345000000004000010301c04040c00040000000000c000000000000c0c05100000000c000000001100010000000030070c00030100000c00040400100c00003000000000030000300c000010000000100000000000140;
rom_uints[719] = 1024'h41c7034c0000400000000f04430430040104010407f000004c0d000111c000c000c30c01433005030000040d0030000400cc0400d000400c40050541100000330000001c0044c410000040000030033000013004004000000010440540000333c00540c403000c4f0000000c000000cc0c0100cd4000000c4000340104c10;
rom_uints[720] = 1024'h700fc003033c03c00004c0c0001000000100c0c300430000003000004c000000404c0cc400007000c0001000000414000403000010000014c00000001cc00c000f0d400004000c30030004000000c3000000030cc0000c0cc4f04000050404f00000000c0110c003000040010004000500443f07c500c0c0c4101430cc04;
rom_uints[721] = 1024'hc000f1040000004500043cc00003010c4000c04073001d000001000000c0cc03d0030000c044c0000101c0000f0100000040010040000040c03100010f03130000c100003c013103c004c04000c330011001000004004030c3010000000041000000300f0001000003030343000c1041c031c100000000001035300040010003;
rom_uints[722] = 1024'h4c00331c004d300000030100c000004000430000410cc0054c03f105d0c0040c07030cdc434140047700000013c000310301104c00000000300000000f330c40c04c00f04470dfcc1000c030c00001001d00000040100000c303c170d00000000000000003c333003ccc00000003111010010100c0477c000170000040040cc0;
rom_uints[723] = 1024'h1031003f03000c030c00c004c000400000103304001c00300000c10100cc0400710400000000040044000003010004000c04c000043001000413033c001000000303d0017004d350000000040400100400010c030c10033000300c000004000c00033000141040000000010000300000040004000000000303000003013c010;
rom_uints[724] = 1024'hcfc0440c101f03000003100330000040cc3000300cc31c30c30400011310014c00303010101c1000010d4f00000000c000001000010000c000f00f0003300100000c3014000000f000100040400000000c0000040030c400433c0001047000c3040cc03000040000001c0100000000f100030331400cc00000c00c300c000c00;
rom_uints[725] = 1024'h3000100000cc000000f000400033003034040c000004010000000c00400050104030300030030104100130000000000000300000001c31341cc000500010000030000100400000000c030013000004000001000000000000507030104000100040033030000000000000000010c3400001000000000003001000000100000001;
rom_uints[726] = 1024'h430c0c000034140c00100c001c00d000000100030c3300700004303c4000d1c0440001041040004110401000040000040000014c34100440c04000000000104f00150000c30000c00004400004c3734000040040000003034d300cc00000c04c034010d00030400c4010440000000003c300c001014000711004cc57c110c;
rom_uints[727] = 1024'h10003000c00100000000000030c000400000004000d0104300000004000000400040000000040005004c11400000c00000300310003407000013010000c0000400000000000000c00c0000300330040000c0033300040c0000010000000707c040000d00000c00000000004040c00004040400000000010000c0040000001000;
rom_uints[728] = 1024'h3040103000000000103141000070000100c140400000f0100350501c03000330000001400040c0c010000000c01304c000000030003031001100405030000000f034c04004105040010c0400400030c0000400c030c0c001300400007000000000003430410030007000c0300f000000730307d000100010031c001030d0c140;
rom_uints[729] = 1024'h1c44d0c00c001000010003301110010000000000300f0403000440cc0000001000c100001c000003011c10c10340100400000010c400400401001c100c0000c0f0000000000030101030140000000000000030000004300000c000030000000400000d000003001000001400000000c300004100400000030000400d000100;
rom_uints[730] = 1024'hcc00c000340c40103000d00cc10000c00030000c4d033c00000000c00030001000000300c010003043310700c00000040000010f700010000300000004000d0000000f0004000140401000000c400c000c0c00001f0000010c0000400004000001c05c4000300000100030000040000000c3cc300400100140cccc3030040300;
rom_uints[731] = 1024'h400013000000d00000030000c0000003000334030033400dc4401030004400000f43101000d001000000000000001041000000070100c0000404c003000134c0117001000704010403000001010010100000003010013000c40000300040010000040000000043003000c000c0000000010c30000000000f043c004c0;
rom_uints[732] = 1024'hc01400cc00000c040001400050010c013003010000430f00c30c00000040c00d0004030000000000044c0000cc0c0000300001070000050000c0003000000c0104c00000000150000d04000f0c3c0c000c0c040000000400f0000000cc04040007c010c0010c13100303001000000000dc000000030403300c001000010011f3;
rom_uints[733] = 1024'h310400300cd004f03cc03300c0c1000330d110030d0753f0cc400000c4f005100c0134000000c44040c1001c000030d3030010000c1c0c00000000c340001040300075f000c0c1c044d001cc0300400c0c3d40000000401000f00100c0c013000500f0000100004000d0c00040470000000005030c0400000000400001c0;
rom_uints[734] = 1024'h1130040c40c40cc0110c4c00c30110c00000000074400cc040040470c5c00000007430041dc0050000d440300c00cc00004c0000c01cc000000000c4004104c030000000cc00040000000340c00f4c00c0000c0000c010300c43000444300c017010c0143f000cc4340c001000004000f0050034004c00001000c0000400c;
rom_uints[735] = 1024'hc400000104010010c3c00043c3c00030c0110001cc1f00400000101c00c0c700030000410041000c0303d4000c10cc701037001c00000000000000030000000401000040c0c4c001001400c0407030c033c003c33040c044c0c00000001050430004f0300c010000030000c0040040000000034000c00000c01000040fc0400;
rom_uints[736] = 1024'hc3000000f030000000003cc003105000000000000030403004110300004000c0001000040000301c1450000030c010c143c00000c040000010300000010000000404000c0000c00050c0400040c03540c00300c000000000013030c0000003c0301003d13330c100010300000111000000f0000000c004f00170100004004;
rom_uints[737] = 1024'h54000c0040400300000001f30030000f000d0000030047000001400300030100c11cc0040000cc000cc31d10000c4003c300000c404303404000000100440001dc00100cc00000040300000043cc1400d30000000105410000017001040000000000c00000000c0033700000000dc000000040c010003000000000c3c4010043;
rom_uints[738] = 1024'h10074000000003300c000d30c1000000003000033300001000000070000000004000111000305300000040003000000000300000000004c001100030c10c0030010000104000103100004003c013107c005000000000c00000403134d03001c300301100100040000100300330001001000003303040c3004c30300000040c1;
rom_uints[739] = 1024'h3000cc0000430000005000003000001404000030c0c0000c0c03310c0030010000040000540d300401cf0001343c030000c00000000100300cf0040003300000003100c00000000c000000d00000000000300000350c0c400040040c0000c00000004000c003040000010c1000000434031004c0cc4004c000045031000c0c0;
rom_uints[740] = 1024'h30010003010040110000310301000001107d00c01033d31014013103000000000000011300010340000000000c0040000f000c0003000001010031400040030400000300010530000000000010000003100c00404000c00030000000c003000d31c037000300000001033c0000003003400000330010000000000001f1;
rom_uints[741] = 1024'h4000100000000c301c000c00c300c000010000dc00440000040040cd0004000000c000440010c0c0103040cc000040030c0000c03004000104000000000000000000f004401010000000cc0010c14004c44c03000000d0c0c00cc004000100fc0d0344000400c0c00400300c0c0000004000304000c00c400400001c43cc34;
rom_uints[742] = 1024'h330000000001001c00cc0c0000c40140104005001704300f000f400c0005007f0d03010000400000040c07000301000300040000c1003000000704400d05030c00013400010c0014040000100000c3050000000c0000c40000040141f00cc00013cf150473004110c00f0010001404040301000c0000c00304000000050c0303;
rom_uints[743] = 1024'h37001c113c000003131c001040c0400311500c531cf3cd3030370004310301c30c30d03347c00440110000103c3d403d10c030101c00000000001350000301000003003030301d53013310315f010001000c100c003505300000103c003030c00050400000303300073043c15c04010030373c0030f001000004000010c44;
rom_uints[744] = 1024'h3000f00f1c00003c00030300131431000005c43013300d3010030000c0000030377cc1110cc00fc01c43030c000103050400040010003044040104030104d33033070010c00000130101300030340300030c00030000504003400400000c00004034041d0000000010000c00300330000cc00000000040730303033303007000;
rom_uints[745] = 1024'h4007000003003c000000000c7000100000004f00003303c0c03011301000003140c0001c307c000041101000000043c3003003c500000c00001010430034cc00c000333000300303500005000c30100300c00300c000c010c00030000000000100401010000c000330311000000100300333303000000000000400010000100;
rom_uints[746] = 1024'h1c40c000000004c10130030c30c0033430c400f33c0000004005d0000001d00430100000000000400400013004030033c100000c000400000dc004000000040c0000000000003001100000100c0000c00000003000300004030000000cc004010030c00000000c04d0000400c010030c00000000400030000000004041004;
rom_uints[747] = 1024'hc030004004000000001011004000410000c00000000400000000000004c004007043000400f01300304c004010c0003404300000000004000300000400c400040c10c0310c0c00c100300334c40f0c0303cc0000f000000030100cc500c0000f700c00c04301000000100003300001c0000004040cc0000043c430004100004;
rom_uints[748] = 1024'h34730000040c3400c00000c00101300000f0000000c0c310004000400000004000003100040010c0c004c00040000000004000d04001103000007000c0d000100000310cc0030031700040003010001010300c0000d0031000000000001100733000c03101030c0043000000000013000000004000c40040001400000c0000;
rom_uints[749] = 1024'h1c000040c1044000d4c1c00000cc00000000c100d30c0c403c00003400c000040f400000000401000040100000031000044000340c010000c010cc0040000001300ccc05c3c050c0c100301334c0030c300c0400c0400400f10c0400104000cc40c0c30cd0004300710040400430000000c0c0400410000340d300000c000000;
rom_uints[750] = 1024'hc0c1007003030000c003030f0c000001000c044007d704300c0c040c430100000101004c30ccc41070c0000003033001003000c00c0000c43013c0000000000d3004100040000033404000040100010010400404100000310033030d370510103013700000303000d010004400310030001010013000c000001000000301000;
rom_uints[751] = 1024'h304040c030000000000400040000000030c00000f000300f00000040c300045001030450c03000cc01cc004000c00000000500004000cc0000300000f000000003cc00000c00300000000c10000000030000000000000000c0000000000004004004c0310000000440000c0003000f0000000010000000000000004410310c;
rom_uints[752] = 1024'hc00000000c00ccc300300000c0000030103303100000404030003054000000c0113003440004000c1c0340300000003100000000000401f00013000004c0c0c3403000010f001c010c4000410000000000030000000134330010cc0000c0043040011030100000000c40330033000000000000000300000000f0000440;
rom_uints[753] = 1024'h140001000040000003c00000040c311347400300004c000030300000000000c0c74100010000030400c000000c00000004000001c0000003000001c407040014400000003c00400c040000310f000c0000c0c000000440c0444000100000000770d00000100100000130074300cc0000000000c00004400030000000c000000;
rom_uints[754] = 1024'h4cc004000001c0c0010c700300cf303000000cc0c0c4100000c5c034000004c00400000300003000047c4c004040c0c40000c0000000300c100d3d00c0004cc0704c01140440001c0010300000c0000d0101c3c030c3004041010000003000000c0c0c01c004c0000300000c040040c01001010404000000000040000c040000;
rom_uints[755] = 1024'h30004c0000cc0003001101f0011400011013000140007040330000000300030000000300031c010303311f00000010100401010f043301500301010000001000c000c01c000001400040c0403000c00041000000cf000400c34400410000000000c044c011000000cc0300000c00c00000c03f400040003050c00001013000c0;
rom_uints[756] = 1024'h301000000004f0410040401d130000001000010343330000000010c1c00f300000103000c300054fc070003000d3001100040001c0f00000f0c00d10004300000000103000005000c00000000300001001000101000000cc010000304c40304f00100000f000004070013300003000041030000c30000c00043040c04301;
rom_uints[757] = 1024'hd030000d01c300410310000c1c00004000401010000300000300100001000000cd03300000070c00100c440c0001c30400030c034001000000040c30400000030100030001c0000015440044000000c00dc00000000410c010c0c00001000cc30cf0000000400000000c03004010000000c3c3300c34030c0007050c00100140;
rom_uints[758] = 1024'h7c03341000033001c03000030c014c01714c00004f03400000400010030001001130010140000000030110000401300003000000004000300c0030000c00003300000d401030007000030103043000041003010304000000000400004f130001c300000030c0010001140dfc0030000003004404150d3400c0000007cc4100c;
rom_uints[759] = 1024'h340c0300030010303730c0000d543000100000300c10c03004000c173f1000cc00411000040c03343003d3300030000334000c00100030300000000c30150000010000003000c010100cd00030103000f00003030014f000cc400010110003cc30303500103c003c100c00c03c4c001000100c10001030010010303040303;
rom_uints[760] = 1024'hc33000010300307000100000c4030000c0100151500c007c1033d0011c0000f3d41300450030003304030f10000130450041000000001000c00003c00000c313005ccc30c3c00003c00000000000c500300341004000d0d34101004c01410f000000c31300c0000030c010f0003100714000f300010010010100000c0000;
rom_uints[761] = 1024'hc0c0cf40c1c70330cc040003c04000304003f000000003d300c0000000c0000f0370cd30c00ddf011000050c000000f0400000000100f0300c01300070004100fc01c00cc0c3004330000040c000010000000030c04000000c3010c0000c000040c000c0307c000000000070c00300010c00000c001000004001100300c03010;
rom_uints[762] = 1024'h100040300400000c01001cd40d000c1100010004003c00000730431001c030041000400c0001000400003f00040c0000340000100f0010cc0c00000001c0040c3c3000000c1504000000000000300c000040044c0c000c400000c400003c000d11111330004040000000000000004033003000430c00000c0001001100;
rom_uints[763] = 1024'h40003310040030003c00000301000003007d0000103f1f004000300310010f00d00c0c0030003c0034003104000d4c0300c010411000000c000c0400313c0400000030310000300104000040003cc3000100000040004110c1440c00000003000c00400000000c0c0010000000001031100c000c4001400c0101000014000000;
rom_uints[764] = 1024'hf0003cc0010d034d001c7100004403000000000051c0c000c40c005f330c000000440033000d004104c100500003003c0040004c0000340400000003001000404000001c00300310031031440010000011c000000000040000070000000cc03004c04303000003040100004440103400403d0c000000003000300c0010330140;
rom_uints[765] = 1024'hd033000000cc0000c00031004000000100000c00001cc000c00fc000000c400003300340f00000004001cd030000c00100c0401000c300d0530c4400034010c0000040c0000001000303c007c00000010d01dcccdc00c00101c0c05103c40000344340000003f0c70c130000000040030010d000cc00100001c0c3010140c000;
rom_uints[766] = 1024'h10040110004d03001000003000f00033013400c500035100c3510300000104407034c00000110c003400137103100300c1300100000130c01010003104d033c0001310004c007400000400341000c01310dc00300df3c30c10030030400011013430030740444030030c300700000000001d100040303030000001000000f110;
rom_uints[767] = 1024'h5c14017c070c0000c0030000003140c000c1400c30050c0000c0c00003c000000301010401030000c070000030d0c100000044000150040000000000000c00031400311c00c00c0110000010011013040f0f0c3100c0000f430000c0500170000004000100c3d0010443c0000c00030400040f3000040304703400000cc3c00;
rom_uints[768] = 1024'h40000000030000003000000000400000300140000000410000c0300000000000000031000000c300000001d0c0000003000000c000000000300000001000c1c0003000c1000000004000301000010000010000000000000000330000000000000030000000100000c040001000000000c100000000000000000000c000000010;
rom_uints[769] = 1024'hd0000003000010000001000000000000000033c00000130004c3400310000300c70000010001000000430041400000030001000000007000004331000000f00004300300300003400000000100004000033001000000010300c00001411344c000000000000000001000000000000000401001004c013003300001000;
rom_uints[770] = 1024'hc000c000c1000400000000003c00000040c0c030d100000110030300c50000000300300403014000c034c0013000000000000040000000c000000000c1c000040404c00400003100c300030000c00000004000c10040010541000300000300000001100000000000004070000000030004000300004c000050000300000100c;
rom_uints[771] = 1024'h44000000040430000000440000000030000704400c1104003000000044040040040c4c0430007413000004003fc000c000c00000001000000401c0000044000000044430450000403400f0cc030000c70c04d00000000000c034c000000000100c1034000000070000cc00c000000100000000cc047013000040000000000034;
rom_uints[772] = 1024'h30014000004043000c0000340003003c050c001403510c040c000341c000c43c040000034700000000370000000003000c010004031c00000033000074040000004040010004411c000000107f404044340cc0004c000010000000000000000010000700000140103f40000000410401000100000300000c11311000000c000;
rom_uints[773] = 1024'h4040000000400001000040004003010000004000410000c000000000014300030003c300000000000304c000000300000100000000400000000000010000000000410000000000c00000040000000040c1c000014303400000000000430000000001000000000000030000000100000000000001000000c0400000000001400;
rom_uints[774] = 1024'h300000104c00300000000000000003000000000000000000000000010000400000c000000000000c0000000000000000c0000c0040000000000000000000000040001000000000c00010000100c000000010000000000000400001000040000c40000000000000000000000000000000000000000000000000000000040000;
rom_uints[775] = 1024'h1c0000f0700000000000401300000000000010003430c0007000340c00c030001010f031000000001051000000000010300000c040000000003000103030000010104010f000300d10c1000040004040040000300010000000000000010130503030c000004000000000004001d0000000000000c030001300303010001000;
rom_uints[776] = 1024'h3000000d040300030010530300050c400300001007040c0cc00100170c0f030300010400000000030cc0000c010c1c000c041400071f0000013100000300001030c03403015003040000000000340c0c0c000003000c03000c0000000400300003000d0050300f00040000103300000000f000400017c30c000c000301000f0;
rom_uints[777] = 1024'h40c0004000000300000000000c00c041000104000000400000000000c04c000004000001000000004c000000000000c100404044034400040000c14104000000000000040004c10000000000c14000000400000c4000c040000000c04304400340000000400440c3000041000000000000000cc30400000000c400000000;
rom_uints[778] = 1024'h3400c00000c00103100000c4000000000c004040000000000013300000000000c000000100c34000000030c00000100c0000c000045101004000000000000000400000c0000000000000000410000000000c4000000000003071001000000c0004000c3000c00401c000000400000000000000dc00000503050303cc00000100;
rom_uints[779] = 1024'hc10104331c00c301003000000010c1c30c001005130c3100001000000100000304310340541d000c0500c000030403000c0c000000000034000100000044000003300003c00000000001c301000301c03f040000c0000000030000040100300001400005c0000700034100010c00000000000043004d1c030000000000000d04;
rom_uints[780] = 1024'h330030000030c000000000c010040c003004000003ccc00040c00c300c300004c00c4400c03000000000700000d000003c000c401000000000c0000000040001444c7030300c10c000401010f04c004070000110003030c0001000000040000010c00000040000000000100003000c00003000300300100040000c0040c0040;
rom_uints[781] = 1024'hcc0030000030000000c00000400c00000000000c70400300f00004543c00007404c003000000030000000c300044003c000030000000c00000000030d0003040000000300040700000000400440d0300000000000c000030003410040040000000c0000000c0300001100300000000000010000000004000100010000c100000;
rom_uints[782] = 1024'hc0000000000000000030000000000000300000000000000000000403500000100000300000000000100000000100000000000030010000000010000000010030000000300000000030000000000030003000000000000000000000000010000000d000101001100000010000000000000003000000000000001000;
rom_uints[783] = 1024'h3103c100000000000c00c3c14030003010000010c400700c000000004000c0000004004000300003000000100000c000000c04100c301000c010000014dc00c0003001303004043000005000c0f030c01000401c700000d0000000000000100000300004140050100004000514c000000005c00003101030104003000c300;
rom_uints[784] = 1024'h10100000300000000000003400000c3000300010040110004030c0000034503440304c40c0fc1000000014c030c310000001300000d0400000103000000040100010100050000c00000000303000400000003000c000000010003000005000c0003000100040d000303c00000000004000001030001300000010003000300000;
rom_uints[785] = 1024'h30000000000030000004310003000300107000070c0c1000004101000001000000000030000c01010c0100000000001030000010000300040133000030133000100001000400000004000100010000c400310100000400000300000000000000010f0000000000c00c000001000011000000000003c0003c00000003040c03;
rom_uints[786] = 1024'h4003c3010000000300000001003050005300000400c0000030010000c00000030300001c34003040030000c0000000c00100000045000040010000c040100300000000c000c0040100000000140000000000000000001000000001c0000300c00000400030004040000000000000c000000000000003103000000000001030;
rom_uints[787] = 1024'hcc3c040000c0003000003300305440704015031043c0c070010000c0c0f000400050c3010300300000000c00040000401000000001c340c0004c000000c0400000c0c10030000030f0000c1000000300000000c50040000001000000c00340001000c3510001100100004000000f00c00040000703034500404c000040000040;
rom_uints[788] = 1024'h4000000000000000003000c000000040040000000000300c000c000000001040400000000000300040000c00000000030000c0d000c00030000c000000000004040030000000140000000c4c000040000004c00000000000c000040000000000000000004c0000000000400000000000000040c0c00000c000000000c000;
rom_uints[789] = 1024'h300010100000300010c00030c010c000700000300003c0c4c0004030003000c4f04014004c000000f030100000041000f000700c401300001010000c0300040000344000030000100004f010001000300040004000000000c00000000c0000300c0000000400000400c4f000303030cc707000000430000c000000c00010c;
rom_uints[790] = 1024'h3000001030000000040400000c330c000300100c0c0004c1003000303c0031004300300cc400000011000000000c0030000000100000040c04c00c03050010000000300010c0000c000c44014000000000000403000000000000000000000c04c000100c00000f0000011c14000034003030000404c0c0000040d4000c0c;
rom_uints[791] = 1024'h3004040300000000000c03000000300c300c1303000c00000031004c04030400001000000100450000000000000000000c0d10000400000000000000340104000500333c0000004c00000004010100040100000001000000000314001000000c00004000000000404c0000000000000040000c000000000400000000;
rom_uints[792] = 1024'hc100000000004004c001000000100000cc00000003000000c7000000000000c400004000010007c000c0c0c000000043000c04c003f00040c003030007000040400c0003c4c0000010004040c04c000000004000000700cc000000c040004000010140c000c000004c03c00c000303cc0300004c03000000c1d04000;
rom_uints[793] = 1024'hc0030300c00c00000000d000cc0000d101000001d000030003014040000000c0c04003c0000000400003c000004303c00000000301000070030000030103030001000000c4000100c0010043000000030000400100c0000000000040000000040040030000010101c3400040400000030341030000000004004004000003000;
rom_uints[794] = 1024'hc0000000c0f0c00000400000400000000030000100c0c0000040d03000c000404000c000000000007040000000d000000000000030c0010000c100000000004000c000000040c100c00000000000c0c0f0c00030c040001004030000c0003000400040000000000000300000004040000030c0400000c000000000004000000;
rom_uints[795] = 1024'hc004004010011000003010073040c0000440000000140010000000d0711030340000040000100030000030000000001000100c000000c00030c0040000040030000404c010100004000000000100d000000000001010400000001c1000003000303000c30030000010300000000044443000010000000000000000000c00000;
rom_uints[796] = 1024'hc0001000030000100000000000400000d0d000c304300000340c1040c37000030000c30013c010c003000000c00401013000030401000000000000000000003000d00c00000004c0c0c030c0000040000040000000000001d0000400000000514100004140c0c00000000000c00300c300c04004000000c000003;
rom_uints[797] = 1024'h10000000000000d40000043501400330004c000000d000004000030c05000c0030000001304000003001103000000000005c00040010000030c003004000c003101410540300003c000004700c30c0100c033070130000c0007000030000004410f0000000103100010000030003000001f0143000004030d000000000030330;
rom_uints[798] = 1024'h1001440000c00030000010c4000040000003000004041100000004000c0c0400440304000001000000000000004000000c0000000300040cc40000000004300400041c3c05040f400400000004400c00000400000000001001000000040400004000000000000007040c00000000000004c0013300000104000000003003000;
rom_uints[799] = 1024'h40001003400000f00300c00004000000100110000d3001304000101300000c71000000d0730000335100030c0000000000000c3000400001000000000003040001031c0000001000404073000410000c00400c304170300000c000000400000440c000304000000007007000000000000003010030300000c00003300000;
rom_uints[800] = 1024'hc0d0004000000000400010700000000004c00000c000304003000000013010040fc00000010040301041000300004000c00000c000010000c000031000c0400c01000000300040040000000401434000000000003000000040000000000040000300000310100040700300300010030030c0000001000000000040004000c00;
rom_uints[801] = 1024'h11300003000000c00040c103000000cc00c011010c404000c340037300c10000c0000f000000004000f3c000000300400000000000004003000040000000000000c301c0000000000000000c40004040c040000040c3c00000c140051c0000000000c1c001040300c3440000c000003c00000030000000c30c000dc7f0003040;
rom_uints[802] = 1024'h30000010000000000401000300000000100110030003300c0c00030000043001033c0000010103000c00000c00000000000000001000000011000113000301000d000105000c000430000000003c0003010005000000000000000003000f000003000000010100000030030000000300000030000400000001000000103001;
rom_uints[803] = 1024'h3000414040c00000300000c0000003400003007140000000040041430004030131000001000300000000010000c000430c000c00000001c00400c000010000000004000100000000031140010140000001000000c040030044000000c0001340000000000010c0000340c3000300000000c00000400010c300000400030;
rom_uints[804] = 1024'h10300030000000000010000030300000040000001010300000301030501000003000003000100030f000000c3000000000001000000000000c00000000000003000030003000010400003000000c10041000001000001000c0001030000030300110003004000030000000000000000000000000000030100000003000c030;
rom_uints[805] = 1024'h110100100130033100000000000000030030c10070310000004f00010300003300000034040033100000011100000000000303010000031100010000000403131000000000000000000300010101d000000000100000100700010000000033003300040003030000000000c1300000400301000307000301000100000403;
rom_uints[806] = 1024'h310cc00000011000c0015043000000c00000000100003000c113000000100000c01004000c0001000100000301000000000403003cc000000004300310c10000101000000000100400043cc0f0003000d70000001000000000000000010004400003010000000003000400000430004000100000000000003000000311f0c;
rom_uints[807] = 1024'hc0000000000003001104004000c0000001030100f0c001000100000010140100433300001000000000000000000000700c00000001c00c03c0000c440010000000001300000000c30030010000400000000c00000000000000000000000003030303c004000000000100031000430000000000000030000000040000010;
rom_uints[808] = 1024'h7000000c00100000000010c0000000000004004003000c00010040004004c004007000004c00004303c030c0000000000010cc0010400040000c047070fc000034000400000030000c000c4ccc0000c00000400c0400c000000c4000000000003000300400c4000000000c4000000000c000c00030c00010300c000040d000;
rom_uints[809] = 1024'hc0c00000000004c00003000c1070c3010000040000000000000c00000000c400000004100c40c40000000000400c04010000000f0007000000000c0401000000c0c30443c405000300c0400c0070c000000000040300c00004004c41c0d0004c1d00040004000c0040003000003c00000000003500000f40c0000c0140040700;
rom_uints[810] = 1024'hc000c0000000000010040010c34000000000001043400030403011000000141000000000c0404000c000000000000000000000000040c0000000c000001000400000c000d010000000000000404000000000400c00000000000000301030000000000000000000000000000000c0c0c00000c0410000000000001cd0003030;
rom_uints[811] = 1024'h40010000000c4010310101301000310000000000333330000040000140030030000004003c0100300c53300c0f00030001010000130100003301004741000000011000c000300000400c3333010000400005140030001013003100c301300000341d03300300000c04300000100003f001000c130000410000300c0000000c;
rom_uints[812] = 1024'hc0c00000010000cc0000000040c14000000000c00c00c000000304000004c0004f0c004004000400cc40c40040444000003c4cc000000c000001000000c0000000000400400040c100c000cc4000040444040000000000004000040040cc0000c0400001000c00000400400c00000c000000004000000c0c0000004040000000;
rom_uints[813] = 1024'h4030000004000003100330000010000000100c000000001004f04000001410100000000000000034000030000000400c00000000000000001000000c04004000d00010100000000c000c3c0c4040000000c00000c0001010000000000000031000300004100003000000000030400040c000000000c000c000003;
rom_uints[814] = 1024'h40400001400000000000040030000000000000c040000000cc0000004c000000c000000000000000000000000400000000000000000000cc000000100000000000000c000000000000400000400000c0000000c0000100c000000100000000000000000000000000000000004040000000000000000000;
rom_uints[815] = 1024'h4000c300c0000000100130000010010000100300000030000000004001000000000000000040000003000000000003030000000000000000000001030000001003000000003000c0030000000700000000040000070000000000000000000010000040000000300010000000000000000000000;
rom_uints[816] = 1024'hc4c0000000000000000c01000000000000000000000000000300000000000001000000040000000c0000000000430400000000000040000000c40040000000010000040c00000000000000004000000000000000000000000000030000000000000000c0000000040000000000000000000000000004000000000c000d000140;
rom_uints[817] = 1024'h40cc10c00000000300d00030c000d00040c0440030c3000000000cc0000c004c0000c000000100000044000073033000000040001300004000000c000000004400040000c00000f0041004c3004000300100400000400001000300040000000440000040c04300000040044010000c0000100c01003000100c100f000c0000;
rom_uints[818] = 1024'h300c14004d0d40c00000004000000043c004000401c1030000c30000004c00440304400000400000000000000004000c0000100100000000000c00100000000001000100010000000cc0100411000001000000000000004000014c043000000000000000000010000303000100040000000000000000010400000c0000000000;
rom_uints[819] = 1024'h1400001000000c00c000000c00c0103003100000003000003000000000000000c00410010000000c0010003000000000000000030000000c30001c14d00c00001000c0100000000000003400300000000c00c0003000000c000000c000000000300010100010000340000000000430303000000000000c0000300000000010;
rom_uints[820] = 1024'hd301030000441000010010000000001c0003000000c04003000370300000000004034cc00000c100000000c00004000003001000003030000070040100310100003000000540000003000c00010000000003000010000030100000000000040001c00400c0100000003010030003000300400000c000300c001000300;
rom_uints[821] = 1024'h3000040001000100000c400000400300000003c04c011301c01040010c01030000c10000404330c00004030300000001030000000000000007030300004c0cc00cfd001d010040010400074000000300000040c04000000000304040c003c04003c1c0000003c000410300040003000001d140d400034301000000c00103c00;
rom_uints[822] = 1024'hd00c0140030000c001c31300000330000000c010003400000c050304100031534000004000040030c070cc0030330030000000c00c010000c000030000c04304c0c0c000010103c313030000011cc0c040000401c400000000000417000400040000cc000f4c004000004c00000040301030054100000400000000001c040d00;
rom_uints[823] = 1024'h3000000000000000000000101030000001100cc010000000000000c000710000000000100000000100300400f0f0000300000010000003000000000100303000004000131000100000100000c0110000001000c00000000c040000003001100000000000400040100010003000000030003000301040000000000130300;
rom_uints[824] = 1024'h34000000000f0010140c0c11340400310c0c401c0c000c70441c00040010040000c000400c3000f40c0000040004000404400050344000c000000410cc000ccc10440000041c1c0000003400043000004000410000000c0100140c0c30400cc0100000000c00741c044c001004040c3000040c0044340c04003430140c0c;
rom_uints[825] = 1024'hc00000030000000030000070000000010001300003c00004030040c00000003101400000c0c00030000000030000003000044000000000040000300000c100000000c000000040400040000c000001c010000000000000000000000c0004000000000c00500000000c001000000000c4c400000000000004000000000400;
rom_uints[826] = 1024'h30c4000000000c04040003004cc00400c00000000000000000c300c00000c0000cc00000000700c0400144c000430000000000000000000c0000000cc3040000c4400040c0000000040400c00c0000004000000000000000c0000c400000c0000003010400000000004000040401000000c3034000000f004000000001000000;
rom_uints[827] = 1024'h13c00000000040010040000000000000c04001304000000040000000000f3010c3044530000000030000c00c0300400001001000f10040000c043000010000010100014030004001000c00000000c000000100000c000310000000c00140c300000c001300c10040400cc0000000c000000000010040c0040d1c000000;
rom_uints[828] = 1024'hc00c0000000c00400010100000000000000c00044000fc000000004c00000404004cc0c0000c00000c04000000c0000c0c4c000000c40004000000000c0000001000000040000c000000000430000c00100c00000000040000043000040cc0c004041c0000000400000000004040000400c00000000c00000000000c01000400;
rom_uints[829] = 1024'h3c00000000010000000300c040c00000005000000044000000c0000300004043000c4000000cc00000d0003000404000c303c0000000010000000000000000100010030000004040000000014000c00000000400300000071130000000003000000d00400000c4030000c00000000000000000000000000000c00000004000;
rom_uints[830] = 1024'hc0000100000000000003f31400000300c310d04343010000c300000300c0c3430040c1000000d1000300110000000001030000404501c000300000000300c0c000c00001c3030300d1400040c000000000000051030000000000c30000c0000040000003400010030103004043400300c1c0c3c140000001300000031000110;
rom_uints[831] = 1024'h401030f004f0cc50000000000004c00c00000450c3000c100cdcc0c3c400003ccc400030c050dc0040005030c0f030003110000c00404040003cc0000030cc4054044100c400004000000010c00c0040c07004f0c0c030400003c0005010300000f030304400000100c0001050300000000000c00c00103350300030000c4c3;
rom_uints[832] = 1024'h3c043f040f003004000f00c014033000100404131104100004000010403050000013100400000104cc004d033030000000000c031000001000030000040cc0000c4030017c000404001c40131c10c10f104003000003000000f0303000000030030501300010000c0000c400101100d0007c001010400000700130c00340000;
rom_uints[833] = 1024'h3003000000030010410c0401c4000070000300c000c70c03010303040c400000100f4401004001000cf3c0000300404000000000000430000370c003000c313300003040000300c34000000000034001030100030000000307000050c0103000d0400030700400000c000310000000400400014010000043d10100300010030;
rom_uints[834] = 1024'h4fc04c4000000000000004f000cc000c0cd4f000c0000c0010430f4000cc1c04000c0c005c000c005ccc0000000c04300040c0040000000000c300c01000404050004040000dcc0000c000000000007004010d0000004001000300100304c4001100c0c000c030040001d000000c34404000000030c404304000c1000300;
rom_uints[835] = 1024'h3700000000050c3400337533001014041f0004534f5c1311300c000c30040d07714cc0070c0c34100c07c40130c031041c3000f41310000c00043000100100003034350301040000000000131c0013143030c004340c00000134100c1c101010000004000010043cfc100000001f04003c003001000c13001013110450011030;
rom_uints[836] = 1024'h33c030000033030030000100c013007001040053444400001c004341cc011430300545070000300400c700c34005040000100000140000510343004000031f1000000030c3434004100130104300000030c0000c0c00c0003c1000440300000c117437470440c110330004d0334000001030f40030001040c100004c03fc000;
rom_uints[837] = 1024'h100000000000c0010000013c000300400413000001000130c0c00100c0c00400340000d0030dc0000004100003c000000000000003401040c0c000c0000030000c40100000400100040004c13100c300000000400003000000403fc003004004010000141010030040000444000000400c000f0430c003c0400303000000000;
rom_uints[838] = 1024'hc000004000f000c000000004540000000000000000011040c0000c00000000004000010040f30000f31cc00000c0c00000000cc000c004000000000030000400c000c00004130000000000004000000d00000400c3000300c40001000043400004c000000000040000030000004000c0000cc00c30043000014043031004c04;
rom_uints[839] = 1024'h413041c045c0000004c00100004c0010c3c0533cf031c000743f0c0100d4404010030d0100000cd4005100403004c01000404100703c44c310000050c3c00000d300001100c0c0c040f040400000014000003300f00cd00010303f040040f050001110100041003c04005440131051013000005010c001000c01300c031c03;
rom_uints[840] = 1024'h10000c01033000d40c300030d4303c1400307040000f1c13000010f000cc004040100331c0330003000010c134000000034c4073003014d010503341000000337fc0c5c40c7003c000004c04c033c0c00130000030c0d10f1070000300000101003440010c3300c41403300000c00f03c003c17030c000000130d50030;
rom_uints[841] = 1024'h4d00430000000c0300400044430d000000000005cc304341040d03c1c00c0c000000000001001004000000030040c00d4044000300040300070c0c4003c000000c413c01c0040ccc000001000040fc40401030c003000050400c00c0430403031c00000000073000cc03000000000300400000004700000000000100c001;
rom_uints[842] = 1024'h100c300000001c040100303430000c134004303300c000104c4cc00c00000130003030f00004010030000000110100c40c03300000000c0103003003000030410017011000040003300053000c00000d5004000c0110303d130000003000c440c033000000001070c034030c0000400010dc0300000400043410c00c0110;
rom_uints[843] = 1024'hf1000070304d0000000010044000c0c300700035cc000003045f040041cc330c133030000000100c3004310300070333000000310410000430f0c0000000c0000031313011000030c3000f0000000100c0010000140c04000100101401cc30500043073700000304401c3000300001040c4d00330c0004771f01133044104113;
rom_uints[844] = 1024'h300000c0003c10c0004030c003100cf03073c000d1c0000010ccd000c0000407c10f400000c030403c1030100010000030000040100000d0010cf0000000c010704030507430c00000011310c00c30003040100040c00000004000cc0c0000d3003040003100c000c0000000c0f1003c440400033040100000704c3014c0000;
rom_uints[845] = 1024'hc10040cf0cf0000000c0030001000000033000030405f30f04000403c000051310c033c0010045030001f000044313c1c3f40d3001c0074000040c010043004c0cfc03000000374cc000010700303003010300030700040c0304005104c10000000cc0000004000f04c00c01030cc00d000c035000040d000004c4101010001;
rom_uints[846] = 1024'h350001d040c0001000300010033331003000003070000100000000401000001000003000d04000c00000410030000004f030000040c03000c001cc0030000000000000100000004000010040000000003004000000400000c00300100030000330f05030300010300300c0001140000000000000013000000030c00013003000;
rom_uints[847] = 1024'hcc07d010400100030c30c0033044031f000040045d0d3c01340003c04100000c01c4cc7c400303011040d7000000011c005000c04045033400cf0000444001001333c300111333004c030014434010000cc000000010c0c030c40001001000c1f4fc41003c417000c30d000400500010c3c4c0100cc00500000c000300000300;
rom_uints[848] = 1024'h10000300c030400004c004030400c0f33040d00dc00000300003f04140c451c0043c10000404440010010c0030f35000000c003310fcc0c00314f0030d000001004000005044041110000000300000c00000f00103300000030007c03001c0004c731000405c1400f0000f000301000130300000000fc1300404400301300003;
rom_uints[849] = 1024'h100050000c4030000c170100040343c00130040400310000014430110040000010c40100135c00c41400d0000000031000000c14ff0cf0040300317cc000030c0031007000001400300cf50004304c10000040004000003c0cf040440100c040cc14000c01c00400704300cc0000001503c00301000040000000c300c0d0f03;
rom_uints[850] = 1024'h3000c3c031030130400010c04000c053c07000330dc5c1000000411130010400c3040003c30043330313c30000c00300f0300300010030400135000cc03101030000034014c50001f0000000c101000011100104000000110003010000000000030003000305c000430033f00040000000303041c3034040c040000103010340;
rom_uints[851] = 1024'hf070000343301030f00030c400004c0040d140d00030f003003040f0c000c05c5300330103cc3340110001303051440010c00030100f01c500c0000450c140c0c0f001c00040c0c0004cc0131000c00000c030104400100331000300013040000340004100c01310000304100f030000703000000300000040000004c0000000;
rom_uints[852] = 1024'h30c30050301000000d03004010c3034c00030003c00d51f0300c0f3d5400305300410010500cc0c000d071000003000000000000c0c004c00004400000001cc04304300301001000044000300000c40300000000c1030cc00000c0c0400c030c03100030530100000c00003040c000c3000000c040ccc30030c3000000000401;
rom_uints[853] = 1024'h3500140040000d3000003743f30c0530000730000001000d030d00100000000010430430400433c0103330710c0c1f4000c0100400100000030030000004410030c0c004100cc0400034000001c1050c3000040300000f0ccd03000001300710401003003033430300440c030000000310141410001d030c1000000033c00400;
rom_uints[854] = 1024'hcc0004c040040000c00c4400044c0000000403000000c53000140c40104000c1000003c0300c000051000000000c10c0407000c30104000c003d10034f00f100030343d03000100c0400000d000c000004000000040000000c00004cc0c01c0400c0000001001c0003c40c050050300034c0c70c10040000000c0c0c00504c0f;
rom_uints[855] = 1024'h43030140010130000130f344000000040000004d0c13c01040000044f0040300f0003010000d045041403010000140300000cc001300071000001000000c50503150030000f400f4f030030004505c000c00000000100c0310007040f0c1030000c030000000303704c013000100101c470040f00000004c1f0001400;
rom_uints[856] = 1024'h50413c0313470cc1f007004350cc0010003c0400000041c33133100d0000001c3c00131000c40001001073050031c3510400003c0c1000003c10141000f000c040d03435300000cc0c00c0f40314503c04f0000700000010c470f0fc444010c00ff4fc00d00030073c003c34c0f00003403030003030000c30c000130d07000;
rom_uints[857] = 1024'h3c303300110c00f0003c4d131c04041100c30d0c1df11c00000c000030700f333004dd3d00001c340000c00400000100000c00c3000130470c3011001410303000f033007c0000000c3000044c0000000d0001101f003001000013410c3c04040700300c0c0f0403c0000c04000d004c0c03030f003004070000000030003010;
rom_uints[858] = 1024'h300004c000030c0000104030304003000101c0030f00000010d00013011300031040010013000000031033000000300000f00030000040c00300404300101300013330000110000000000000c300c3000040000000100700300000040100303300004310004043f0000000000000003000000001333000c400000000030;
rom_uints[859] = 1024'h330000400d0c040301007700cc00c04300c30cc05100000001cd430d4343c331cc401001000000000c0000c100000001030100030104003d00040104100f301d4040d3c000404c0000c00001cc00c000c0000c0dc000401000c100010004c0c7174c70700000000040c300c300010304000c04043030d30400c000c70003;
rom_uints[860] = 1024'h1000c33000c030000004c300c041001001c0410001d0100c354100c0000000170000700340001004c00033000030c001030011f0303000000140c0007003c4100030c140c0d01c0000030001c30100303041004000434003c0c00010000c0004040140001000400c400003304000f001310004000000000030030400c000300;
rom_uints[861] = 1024'hf0040d400100c0031c100310d000300000d00c71310c0304070000cf003110000700d05031031000301034000030404000040000010030300330c0030000013c0100001310000c1c53000030c0000000303300010000000004001d3001700400000050030c5c0000d170100000301000fc0400c43031c401000000c00030c70;
rom_uints[862] = 1024'h1331010040001003c1f00040f0c500003100011014100013000014001c47c04070400000100000000100403400cc4040000c34003004cc4c0110000034000c000003104300000100003004070000740000400c030000001000003070000c000400001000000003000000070100c4000c005334c050130c00400000300000;
rom_uints[863] = 1024'h1c1001030403c00c0000034c03300031300d10010c00000003c1010100d3103d000110004ccc030001401103000001007103000000c304310000000001304030500310c100000000031d3001c400000010330004030c303330030303001410330100040071000c01300300013d3000010303030001c3300100000c0043044130;
rom_uints[864] = 1024'hf0d30c0000f000c00010c0015000401004000000d031f070400700300000000070c00000400301041000000007004010cc4000c01030444400040030c0dc0000cd000000c00010c000c0401031001001c0000500c040000030400400010050000030c0131000004c300000c0001303004000f40000300003700000cc04fc4c0;
rom_uints[865] = 1024'h300000000f54f030400c030070400d0001c0015047c341144000400301cd00c01000330303c100c107dd004f00000001400c3014304104c0c000030101500000004000100001c40000000004140140d01000003010000040c0400c1000c0300003f0c0f004030000000043c010000cc30000041000000340014c0034000000;
rom_uints[866] = 1024'h3300031000000000000003001001000003000010030030040c0c00000004030400430000c10003004c0700000000000000000000100c00000d0403101000007c4000000404000000040c040040400000010000000004000c040000003010000403030000000000000300040010000414c00c34000000000410000130040001;
rom_uints[867] = 1024'hc0044000003010000030c400c40c00340004034404141010c0c03450000300004000100c0000300170000000001c000003c0003410f010000000004f301000000003000040400000003400001c14c4001103000330040000003000401000010030303c0000101c010d100000004000300d30305c0000310000000110c05c3010;
rom_uints[868] = 1024'hc0c000010c40000000d0000010010c0000c33000011003f0c040001c044c000004cc00303040c00400c0c0001003003c00c0000fcc4c0000330dc0c033c00c50c0c30440000010050030103010000f00c000400000000010c0c0400df0d11140cc00c130f0000000004000cc0001000c1050034000104c000010d01cc010c0c4;
rom_uints[869] = 1024'h301100401004001030000300000000301f331000c010300000c70313c4000301001003713010315100031000d0000100403000110030c0100011000000007131000300d00000133033f010000071304430104110304c0c3300140c00330033c40000000030f0330000330000100003303c0000030004101000000010000;
rom_uints[870] = 1024'h4400c0000000300c00d010000010743d0c00100010300c304fc04400100004c0003100100001100010010000000010000300c00c00400040041430c0000000110000000001040010143000333030000100500030000c0000300030403000000000001040cc001c70000000040050000f30300000301030000000040c00001c0;
rom_uints[871] = 1024'hc003000f00300105000000110040c70001001000400000c0010c000014000d041100000050000100110001000f000f0143000c303010000c400000000141000000300144c4000140500000000040000c3000000000000000c0000300000c0c0001004300000c000c30000000c44000000330004101004000000000000400000;
rom_uints[872] = 1024'h400010000000003000030400040c3c00c104000000000c00000300144c7400040c1314030c000044c31000dc00000000c0000cc043010033403c004441000040400c03c0000304c40000000c010f001c70000000003000003100001c10000000c00101000104000300cc005000004100cc00c000050000104c000003004400;
rom_uints[873] = 1024'hc0000c000000c40003f071d07ccc31040000000003000c030d0000000104000000c410300cc1003000cc3c030c000000070c030c13c10c01c1c13000004000c4d3c003c4c00d0333c0000c000300000c4400014000000100004fc000c0004c0d034700000000000003c00000000030410007f0c0374303010410004c01c070;
rom_uints[874] = 1024'hc00000000400000341c00c01cc343000030007000003cc0c0004011000000010040301000001000010071f0003c0400003000303300000001c050000434000070c00030041000000000000010007000503000000c000010400000c4300030c31000000041004030000000004034cc0000000001300403303300001010044030;
rom_uints[875] = 1024'h710040c044301141c3c7c00040037300401330101340cc0000010011f7dc004c331140303330c07c07c03000c0fc0f430cd0c400417340cd0003000700c103411000040fc03701c07041f00001105301cdc044000c13540f030011f030047403100100004040f000c30040304d10c0000440c0003dc30005c00000c001c030c;
rom_uints[876] = 1024'hc000000000000000000000000005000c044001c00004c4030003000040030cd003004301000c0004cd40c00040404001003050c3000000000001000000c500040c000000c0000cc5cc004c00431404001000004500000000404003004000010003400101004000000403400003c00000000000000c00c00000040000000040c0;
rom_uints[877] = 1024'hc0130041000500000c000000000c00000030000001c0300c0000000000000c7400400000000400c300004100000c0004000000040c000f00000440010000100070300004d0000001cc00f070004500001007043000000cc0000c000d0000d0c041f00000300000300400c04c0441000000c0c000040c000000001000000c0000;
rom_uints[878] = 1024'h11c000c10000400000c000000000001000000000000000000c4000400040000003000031000000301000000300030000c000040000000000000000430000000400000c000040400000000c03430000100000000000c000001000300001c0c00100004140c000c011000000100000000000030000c4000000103007003000;
rom_uints[879] = 1024'h40034c00000000351351030f4000030000003300300000c1000004001400000000100170000c4000000cc000000100000003000f01ccc3000c00c0000031410300000301000c0003d0004000001130000000000003000305c00007040040050f00030c0000400000101440030003f03000d1c04000c03401014100400;
rom_uints[880] = 1024'h440cc030030100ccc00001c000c00001000000100003c000030500c0001170400000c00c0100c500c5000c43000003000000003c0040c000000f000003010000000c3005c50003000100400000c004f00000300000000000330040f0030c00c100c4100c0c000001000000f3000003000000000100004c0000000100000c;
rom_uints[881] = 1024'hc000c1130000000000000004c040000cc000c04070c0c0310410000c00000c000d470c00000000004000440000000000040c0007000000040000000013d0010000c0c00001000000cd000c443c004c004000404000000030c404000000100040470cc100000c4003000000445040400000c0000c0000430c000c010c00cc7010;
rom_uints[882] = 1024'h400004c07c0100c010c001c00dc0fc4000004cc00000033000c00000007d0004c4044043c0304010400c03cc0000100c00000000000c0000034c000000f34010004040100500000003c000c000400c01700000407c4003004341c0c0300310c00110043c03c3010000c300c0c00000001c01004400c000041003000000000000;
rom_uints[883] = 1024'hc0004000000c300000c0011100540305001c00c00c0070000000437c000010dd4000f010010c1d001004dc00004000000000003c4303105000c0005c13000c0000f00000300001c010400100001c3001c0c00003000c0011300400403c03c00000f30100c00c0100004003400c000003003c30030c0300000000410011431140;
rom_uints[884] = 1024'hc043100000300040440131d00010000000c30c073000000040040c000504f0cc000000004000000c440000000cc00c000c0001000c0300c0301c3303000c0040000040000014003000c0030c01000000000cc0000100010000004000000033001c000000000004400c000010001003000011000cc0c0003000010000030;
rom_uints[885] = 1024'h1c000c3000140c003c00d434c0c40074000c303004001cf0c00007031ccc0c400c430c0c0005d0000000000000f70c300000000430c10033100c3400305cc00043100031dc000050307410700c00003c40d0000cc4000cc413c3c00400000dc5000c1030500f00303400007440000000c00c101c3c10050c300c1c001000100f;
rom_uints[886] = 1024'h130103031400c701f0c400000000310001000003030c31030003d400000033c300040f0007c500c40c0c1000070100000003140c4000010000c01d0000000400c00004c1300c000c000340011c00005d00104c100340000001400400d314040030000c304100000400000d00000000100404051000000c0001303103030001;
rom_uints[887] = 1024'h40004003000000000330040100430003000100c4c5030c030000400300001301c100000103000003410303401030000000000000300000014041000d00000000000103000000000003dd030431001000000000c00040010cc04130c303000dc0000305070c0003c0330001000000000f03000f03010000c0000004400003;
rom_uints[888] = 1024'h3c030c000300000c00000700001030070031000c40000c003c03044000000004000c00c00c7000300030040000150700010300300000300d040000100004100000fc047c11100000d030003c04c1100034040400700f0010003d30140c1030400c34c500000c100d030c0000034400041c40300003100000000040040c540330;
rom_uints[889] = 1024'hc0cc000000c00c000004c040c000000c00000c304100c4100015010100f0000c00400d0c00c0c0000c003dc004003003000000114000004034300c0c00000cc00c30c010c0c0000c0c001040110000000cc00040cc0040000c3c04000700371440340c0c00004043c0000040003c00c0000010c00c040000000404043300000c;
rom_uints[890] = 1024'h4003000300c04000000400000c0c0004c0040311010cc4c3c0000000000003040001400300cc31d0000c030000000000030070004040c0010000000000000044000400cc000000400c000000140000400400043000000c000000d0c00c00000f00100c410300043c00004040d00400cf7030c34004f0000c0c0000c000000;
rom_uints[891] = 1024'h400001133070c1000010351014000004c00c00c000310f000c310040100c0c11100f00d40401410301c03300030c10000034000c030000004040070c034c0000c340000c00450040000fc0c01c0c0000000d00000100c44c0007010c0003c30103c010c0010c130f0103400300c50400400c0c0d0353c1cc0000030c13033d01;
rom_uints[892] = 1024'hcc0c0c00000c30004000100010d0004000000004140cfcc0c040000c300c001c0030ccfc00401d111000000000f004c00000000034c0c004c0d0000c3c0000100c0cf0000c10c0c0033001340c300c00401000c70c0cc01000140000000cc400040111c0103044000cc0400400403000000c000c000000c004c000cc01c01000;
rom_uints[893] = 1024'h4000c0000000000003500000000000004000030004010000000030000c400000c00c40000000c00c0003000001000003c000003030000403c000010000000413030000100c0003033001f0000000000000004000000000000c00000003000030430c004f000000330300f000000000c000100000000400c0c3040c010c074c;
rom_uints[894] = 1024'hc0f44033c00000c01000f313d040c3010f10c4303035d100c3010003000037701071c404013c100043c700c031f0017153f0010304f0c3403d340c005c00c000c1d0d371d0033000d040f071c03d0014401031113c00c0c00300003111c01030731010331000100c31f300443f003301c0000030010c7c00cc1010000403031;
rom_uints[895] = 1024'h4003030004400000d034004c40c054c003035100c0c3010040c0000fcc00d0c70cc3035310c000f000034500004c1017003000300c0004334013400cc00444c3004130d4410300345100c0c0c00003410044004c3100034000700040c100c4c030c0330304d300000001003d0400c0000000001cc1c3c0000d043140400f0000;
rom_uints[896] = 1024'h10003100f00004000003000040030c00010055000010000000300033030101403030000000030340c100130033c000000000c0010100003000300000403c000004100037c000104011040100003c130134f000000c30c000030330000000003100401000010000d100004101010c3103c303f1010000004000030000000040;
rom_uints[897] = 1024'hc0004000000000000030074004000040000000c07f000f0000004c305c400400000004cc0030000040000303c0010340c007000001004000030000400000000300100003010400c010030000000300000301000c0c0000c0030000c0c007c001007000303000000130c0001000000d000300010003300d00110000000103030;
rom_uints[898] = 1024'h10034c000100010300c0000004f1000c015d01c03010000c40371040104c40c00000000040005c000c00400c00100000013c0344c004000c00001003000c004000455c004100100dc10030c01300000100044000000000045001300000004034c0000000c000000000000000c0c000003440400300403503010000000d400000;
rom_uints[899] = 1024'h343c0400000010c007007c04000c0034001004470c5f4f10000c301f31010007710300030c30301c0d073410000100441c000030031034003004000c14110000343401d0410c30105017ccc3130337343004c00430330c300c30103c5c0c1011f330000000501000cf000003c40f04003c01300000701034001cd000000c0000;
rom_uints[900] = 1024'h30f03000007013c00f007100001333000004031300414c301030000503011430c4100500004c00000c0300c000000000c00040011450005103404043c030030000100001c00000c43000301030000000300c0100000c04044010435300000000107703544000c110003000d00340100c00c00000300010030000000000300cc;
rom_uints[901] = 1024'h40100000000c0001000000ff40000040011000000100010c00c00103c0000700340100c0c3c003000004100003000100000000000340004000030030004c00000340100c0000400c04c004013001c004c000000001400f0000004f3000c0000400430010111000000000040400010000000c0307c00043c041000300030400c;
rom_uints[902] = 1024'hdc000004000c0d00000000000100000c00010300001c10f44d3001001400030c30001510330cf0031c00c000000110040030000c101c0340030c0c00033000000040300004004c0c00c0700004000c00c430000c0c000030314000030100400c0c0f0000000040400c00000010000400000c0c0010c04c000404340000030004;
rom_uints[903] = 1024'h14040010075000004043031c0070c300013d003330031c00133000f00d01404000003110000cc0cc40c5530303f000000d075740140004003100c0040c300001300104301000c10104007433000c0004000000400003cc0010030330000003040011110101301003304134540c00010003000004010003105fcc00003000030;
rom_uints[904] = 1024'h340c004c407000000001103035000014303cd000007c7000000c10000010fc300c034004d054c3c0f01c17000010cc3400003000404c34003017c00040434d040000007cc001c0004004c01000004400ccc0c03000000c00c0c040010c00c04000013c0034404c3c0000000450305010c00000f010f1700c010000c13dd05003;
rom_uints[905] = 1024'h341000000000300070110000740000000000400040041434100c1000100400003310040c030c00c040c40c0000040c00101430703004403040500c34003c0000030400d000007030c0003010000413f05400340000000004003c30c0000040303cc0000010c034044c00300000101000040000c00470004000c0000c0c00d;
rom_uints[906] = 1024'hc01033300300001034000000000c3000000105007340d000500c0f000011c3013c4d0301cf1c04410030000010040000070003303000140c000011c0033c003d040000010000044030c000000c00000400430340000c00c101130000433010c4400330c0c004041f000430044c0000000c00c0000c00030007f4003040301c;
rom_uints[907] = 1024'hc1400000000d0030007310c34150000700331c00d3c030103453d43040cc300013f4301c40101033004731c33007300c41101431000030140130c000c0013030303101311c4070301f00030043000c003341010017c0000101f000070d00014101330430310c030140c03033000000c00c0101030000303003c00300403330d3;
rom_uints[908] = 1024'h3c000000007010013030f7c0030000c001003040d0c030c010c01000c00007c3c00c4104c0c03054c0103010fdd014407003cc4010c0100c0140c000000010004041701070000170000110dc000000403040003c5000c00103430cc0007000d3100040003104000000000000c030004c000001f030401000004000c300c000c;
rom_uints[909] = 1024'hc0c400c0c0c00f000004330000000003000000033440f71f000007700003040401f333c0010000c3010dc0c007504f3107f45c000d0007500303117d0c030040ccfd03400050030c00c00100003733c000034040003004030c00074103c00001c01dccc0d304c00347c00d000f03000d00000340c00040000401c0030040000;
rom_uints[910] = 1024'h100000c000001003cc000053001000000000400301300010100000c00000000000000040030001003500000000700000103040c004003000c0100000430003c000000000000300000041000000c0000000000030030000330305100000130130100000040000003000500110000100c00000013000001330000003000040;
rom_uints[911] = 1024'hc307c040403000030000c0000045040000014c0400004c000500030c4100100c0100037d4000c7c11070c0030004c000004040f3414100c4000cc000070000030003030300c000704c00f0037300000000c400000010000000c4001040c00000c0cc10000001000003cc00000010001033f0001003f13500000c000304007010;
rom_uints[912] = 1024'h300701d0330000f0000300041dc0f3000dd000c00313400c03c334000440c015fc004000c044c150000c00fc07000000c30030110000000010f0330000010030010c015004000dd000000070000001c4400c0c00f30000000c30c00000c4000c3301c040401400f000000100c40415f0300303c0430003c001000001003c04;
rom_uints[913] = 1024'h100000f4030c000130000c40000000013000300050cc0c0503001001100000c34310010400cc010c0cc0010000c4000001f043030f43000000000030000cc0000c14c00c010cc00cc04000000400000000003400000ccf0fc40000000d040c013c03001000500711300c0040034000cc040000400000030101700c0c0003;
rom_uints[914] = 1024'h3040c3c00103c003000c00c05000c353304c004001d0ccc0000c0104300130c313000000034d030340100303000000c1c00103330130000501014300037005c30300007007001000f040c000d1c0030010040103000000000313400000033130c343c3010001d030403000030040011503003001c3034310004310001400f040;
rom_uints[915] = 1024'hc0300043003000003400000300043000400100010000c000c03000300000004c53100ccc00003040004000300000000000030030100370000c00000310013000c03001300030f0d100000053000000001c00fc0030100000001703d000004000034010410101100530300000300013033000f000000000004340003003000000;
rom_uints[916] = 1024'hc00040004000c000000300c0030340000300c010c04130c0011f0d50c001030040001300100000050c7000000c000c000010c0c000c0c300c000500000d00040400004000000001000c0000130c03040000000c000c0030034c010750003000010c700400470c000000044400000c0410000c0000dc0000000300007005001;
rom_uints[917] = 1024'h10050010040003000003070303c040c00c740073c050100030101004300130150030130000500c01330c3310100130c030d0004001000001c00010000c000044330f004530100f300340000000001033000000330c0001c0c0000000100d010400303f100374703f04000730000010110100400041003001dc5004c3c00070c;
rom_uints[918] = 1024'hc000030044c47010030c00000450c01003040300445100300404034c1004040001000700010cc700500100300000f0f0007000c00017000033fd1c000c4f31c0000703100000cc0c1400000c1330030034000033c40000140034044c0000dc00c0c00700cc001001c33000010040000000d00000003000c0c00c0c001440d003;
rom_uints[919] = 1024'h305040001000300007c00100c004c0cc0000c300000c0c10330040000c04c034004000000d10401c741c01400000030040c300000cc00300170104000000000c1100000c0003100000043d40000004101000001040000011000000c040c0010c004300c0040000103004c030c0404140100c4440030007000000000401000;
rom_uints[920] = 1024'h34005030300033cc0c0300003001010113000100c01f00000313740fc00313010300443103c040001000040340171f010013003700313d0410f10100300c31c13401c000130c000301c00fcc413c400305430340730003010004030c004001cf00c033f10d013730430010300dc030000313031103030040c30c004030c03540;
rom_uints[921] = 1024'h3c30430c0ccc0430103c1d137c11101100000c000cf110300c1fc430300000000f040c0100011c340c00000000000000000c030000000c03c000010004143d000c0c7c003c0000400c3004170c000000014011100c10071c00401001003c04000740000c110003031d0c0014100d00000c030f0cc03004040004000001301413;
rom_uints[922] = 1024'h3c0000000001001401040003040004000010003030000000c13000300430004c00000c4403000000000300043c00c0100303030400040c070300004040000000100003001c00000000000f3f011000000000000004000ccf04003000000337010004000003003f0000001000000000003003c010070030000001010400;
rom_uints[923] = 1024'hc00000000073c000003000c0300cc30c04403c001cc40000000000d03c13334cfcc30430301001304c700040000000000010c0030c00c30000d0000c000000000103030d4c000344000430c000cc000d0c50003c00c00000000030d00010404030710037070003030000003000000c100004400401000300005040403c00300;
rom_uints[924] = 1024'hd0440300c000040000000000df00300000f00000ccc110000000700003c005d310400c00000003035010704040000030003001300d00300000d000003000d11041c0c500001000d00040003000c0003003010001c00000c00300f0000040000140000030100040000100007040000030003000104001000c334000031301403;
rom_uints[925] = 1024'hc407010001c0c03311000c0010c0000000100130fc0c1700030403304430500040f400500103510100103000c0303c000013000005033c330c0333033041000330c000130000000010301030040c0400000c0c050000303404000d3c013c1004330100031c5c10000570d000003000303c001010304df000300000d00030031;
rom_uints[926] = 1024'h30533001c00c3010cc0c3000010cc500100000011040000000040000011304034030000030d300004430000030000c0003040c34000c00004001030000440730c010430000000001000000000c00cf0400700000000000000c0000000043000304000c101f010c4c0000010300000440000050000c1c003000404000000000;
rom_uints[927] = 1024'h1cdc04000003300d003043400330dc000001001130f10c004cc0010c00031c71c005040000f00c140534510300cc00004103000000c000350c3504c005313070404300f0103c40300011333104341000107300000300043370503330c0d000330100441041305c0c30100011010400c0000c0cc5010c34040cf3700143040c00;
rom_uints[928] = 1024'hc003100170f000004c00c00300100010303000001c00303c000400344c00000700c10000000000371000000004f00010c00011f04000504400130000f0dd004cc00030c0000000c040c0300100010000d00000c0c3434003704007c031304000007010101100304100307300101000c04000c4100000c040401030c000c0405;
rom_uints[929] = 1024'hf00000c04c403c00400033c40470cc0040c00113447740004f03400000c0d0c000f0304300ccc00dc71000404003030040ccc01500004500c40000cc0110c0c0c040300c000100030fc01107f70c00d0c003300000403050c0004040c0fc3000c3f0000c05430430000000c0000005c33000c1c10000030000000004000000;
rom_uints[930] = 1024'hc10330041000400400000000001c00d00303c1d0005330300030c00010000000f4030f0004c43000004000000c3330000000000000100c0030dd040310d100004c41000045300000100400004343403040010000010030040c000000c0000000030f1010c0400000000000000003501004010c40040030c0c400000104000001;
rom_uints[931] = 1024'h30030000301000303004000400000700001304101700000000134000000c040400100000100001000000300000000f0300c03100000000c000041330100000000000307000300000000001000c0410510000000014c0c00030004011033cc000303c000040003001000000040030500c30005c40000000000c010000400000;
rom_uints[932] = 1024'h30344c0014000c030c00100d0303000000000c0415003c0c3330000005c000000c003300140c00001f3c0c0004300300011003f035033030001003030000000c3f0c443400010d500f0c03c0003030000004c033300001030c0400133001040cc00003134040c00004000c1007100100140034030011c0000501000c0100000;
rom_uints[933] = 1024'h100300011300c30040f1031310003101010000f730340c000341000f40001c000030d1001337030d00010303400001010c000103330000030dd10001000000300703030003010103004030000100d10303c3000003000004c0c330300000003000413311013003030331010000f0000000000300010040003000000500010040;
rom_uints[934] = 1024'h100000440030d0f0c030100c1074000000043050f0fcf040c00400140c04c0d10003100000000010304000004000300000c4404010107010003001c0100011cc4000010000001c14300040300003004105000000300000300000503000000040c15004dc004c70000400440040300c000000140000000030c004100014000;
rom_uints[935] = 1024'h30d0041c100001c11037c0f10000000045c4030c0311f010110000c04d30c40100040010401100cc003000c0000401c030f0c03014c071303c0410000c0000001c001104340d10000000d00c00001000c000000000f000c0001c0000001100c44100ccc3c0c010003004000030030304c000c000f01003001000c040;
rom_uints[936] = 1024'h1410000040c00010001000400040c00cc000400040ccdc300030f00070c0414c00003050000000044cc11400f0001c00300040d3030000107c00c0c00040000100c000400004004040000000f0003000000000c003c00030d0dfc0000000c0000001001000001000000004000000300003d0cc00001000c003f0d0300070000;
rom_uints[937] = 1024'hc0c00000700000f00c07f1410041c0f5000c0000030f000140cc0c00000104000000d4530340c01071030000030c000000040f004013010c00d10031c1004010c400c003f0030043040000000300c000c0040c0c40000c010144030000000c40cc034700c00040000003c0000033000040000001c0000300000050010401c130;
rom_uints[938] = 1024'h300004300040c043000c103cdcc0404430300000000040d4000400010010c001c540701004001440001071300000003c00c0c03000004000c00014043000401043c03000f00400c33000c03040c04c0c0d0000c00000c014000330007f0000c01000303050300030000c004041300000400000057100cc00030c0000d4041030;
rom_uints[939] = 1024'h75400541d007140347c340dc01107dc05104cc00c0c00011f3d000407000000c440cd34c0300f040003030400c14311041ff53d104c01cc045c000400410c03f007401c041400000c154cf0000301040c05300000f0041f0300430000041004300000000c04000704d00c010040401017d007000040770c0010331c;
rom_uints[940] = 1024'hd0c3c000000040cc000c00700c44000040431c00000030300c7000030000000031040010000c3000050dd0c40400300003300cc1040411000c1000700c500000c000000c000000530000c00400000c010000010000400000c00040403c00104030000017d010000044000d0000400c4400000040c00d30000000000000040c1;
rom_uints[941] = 1024'h1011000500c01100c0030000000000000004013d35000000c00000100c3450443100030400030000500000cf003040c0040540cc0f400c30001d0c30000003000305d00000000c01f0440004300045030100c0000000031c00cc300103c000c003000043040005c100400501004001c0c040540c000000030300000f400c;
rom_uints[942] = 1024'h4000110000c000004010000300d0000c004400000000000c00c00000000c1003300003340000000010c0000300c0041c00000000130000000000000030000300000000010c00014740000000cd10030000100000000300c0c004000030000101f00100000000c0000000000300000000000100000000c000000110330330c000;
rom_uints[943] = 1024'h300037d00000003001040030fc0010000001370040c00cc01300301c010c300300343010400c00c000c0c000400000000004400000103c04003d1c00000307033c7300c0000000103d303400c0001740000000030000c070300004704cc07314c00000c0d010000001000400040073030001100000c00000c00400000c;
rom_uints[944] = 1024'h10c0040c00000301c0c1c400000303c44010000030101300003c0300000501117000000000000100c4c3c0000c43000003000000004c0000c011000003000300000010100540c1000300c100000c030000f0000030000000000030030000010040003000001040000041400000f3000000040100000000000000000000000000;
rom_uints[945] = 1024'hc040c000c00040000400cc000000c00c0033c0044c01c00c00403000c00c01040c4403c00000c0c00013040000700000030c0004500000400c0500030010c10000c0c740c0000000cc000044c00000c011c0400000000c33c40300000000004c4700c0c0000000030c433044404001100004c00cc0004000000d000000000410;
rom_uints[946] = 1024'h700115c03001000011cc41c011fccc0130004cc00130530000000003104100d4c4334c1300f00100014c30c000000400c04000f000004300004f000400c0001c0c000000c11000304fc00cc700cc0c014040300000700000704000f0000310c004104d404303c50000c30000c40000001ccd000400003014cc0300000040d0c1;
rom_uints[947] = 1024'hc4c0400ccc50c00d0000000140401001000c000034c40004c043c00000001401cc010017c010040400c0003700130d00010ff1703004400f11377ccc0c00000000c03c3f00100c00c0047340c3000c00100030340000100d003c00c030c40040f0110cd0040030003c0000cc00000c03f00f30010000000c0000411000043;
rom_uints[948] = 1024'h3000300010400030000c340130000c00000000001cc74000303f00040c300130000004000300400000c010000000ccc100040000f100303000f0301c0000c10000000000400c00140000400000c000000000000000cc01000103000000c0300000001c04000000000400000000100000005000000030301000004301c0003f0;
rom_uints[949] = 1024'h1c000000010030100c0c340500c40f44000c000004001c00c300040300000c0cd1400c4c100400010c00500000c00c000000001030000000107c3400404000000f1c0030ccc000530070c0700f0400cc00d0000c040000c400d0c0040c0000c0000c1d004c4cc00c0410000470000000c000c04c4c10000c0000050010001030;
rom_uints[950] = 1024'hc410c54303000014010004000c300c7000413010401000c100c0401000400100001000030003c10004fc1c03000440c0c00303101c73000000c00c0000011001d0c00003d1340001000000700000000311100300000000001d10000400c300000030000001400000000c000c000010004fc40001000fc3300340040000000000;
rom_uints[951] = 1024'h30000c0300030100000347000000000300c704000004c00001030c0043030301c30100030001000040c04100034000400000000000c0003000014301000c0000403000004300000403000f0100000d0004010000000000000001000d00000330c10003000104000000c30300c00000000003000003c0010140000301c3034003;
rom_uints[952] = 1024'h300000c00400c0c300c00100010000700c0130c403d3c3c3c4040501070d0000000c0c31c443030103734000014c03400000071001c34300007041000101c000c0c300c0c0000cc1f300c000101003034040400700f001c030c7017cc0c37400cf40107c3c01c0c370c30000300001000703cd0030c0c03103400040c140030;
rom_uints[953] = 1024'hc4c0d000c0c000c01c30c000c04000000001004c300000000014000000f000000070010000c0c0001c707cc004000010300000d4400c035000303c0c70000d00c030000010c0000c0f00c0400c00300031c0c004d10000000c3004005000300440040c000000004300c40040000c00000003c000400004000034000070000010;
rom_uints[954] = 1024'h4003040c03c0400c0300000000030001c04000000f0cc00000000004010000d04000400700cc01000c43000000000000030030044100c0010c00c43c000000400004040c000c00004c0c0000000400400400040000c00c0c00c000000000c00000000c000000340c00004000c000000c3000c04cc4c000034c000c0000000;
rom_uints[955] = 1024'h70000110030000000d00351010003304c00c0001000103000031000c530c4f01100300100005310300c34330371000040000150c030004f500003300030d0000c000300d00410301000c00001c0070c00300c4000d3300000003c04c4003c30100c00307010c0300d103000700050300000c00010340010c0300000110030500;
rom_uints[956] = 1024'hc00c50c0000c000000100000d0c30c04c030000444c0c0003040004030000051004cf0f0000c1c000400000000f0c00cc0cc000c0000c404c0c000000f3000100000f03000d0d0c0004140040000cc305cd0000ccc00001000440010000cc0c0140c0cc000347000000000440110c030000c0c000ccccc0c0000000014000000;
rom_uints[957] = 1024'h3003100050000400000c0000400000101010000101004100400033000c00030050004c040f010001030000c040103003400413c001010000000000c7400340000310000000f00000000001101000000000000001000000100000f043000003300000000701c1000000000310100c0100c40000c001003000f310;
rom_uints[958] = 1024'h4c0c41103c0c0000c0100c3401f0010304010c00c3071c00003001147c4f00470004dc0000133c113030400300103300c5003010304c0034030300c004c40c000c1d0cc01d0c00000c440c070c1300003301030c03030c000000c10f111c01c0073001003500410413030034440000000c000cc33013c7f300011100c0100030;
rom_uints[959] = 1024'h41035300010c00000303404c11c75400000c5000c0c0c50540c00c3f1c0d00c33f0fc1100c00300000037d00c34c0c14003100400c04100c01134c430c303034cc4030f04c00c0f05000c0c0030c10400004c00f713000440c7c413c010404c4300033471403400c0415000cd0c400f00100000c00f3004300f4010003300300;
rom_uints[960] = 1024'h1000000000101000001000000000100000c4d010000410040000000c0040400c00000000000c0c04000000003000f00000004000000c0ccc0000ccc0000c10000000000410000010000004040c0c0400000004000c00c400000000000000000c0c1004100d000034000000000c1000003000000000100000000000000;
rom_uints[961] = 1024'h303001000000001f00000400000030003ffc0000000000400400000000340c0d00000000030000303000070c0400c000400003003300000000040030000010301010000000040c000000003030100000131000313000103c0130001003000000300000000100000000000000300014010000004000000400000000;
rom_uints[962] = 1024'h10170c13010000100004000c03c10000000c0000001004001d040000005010000c013000040c15004c034c000c07000c010003010c0700f0040000000000000001540100100400040000003103010c1040010400100c3c0010010c0000000d00000c1c0300000330030000000010000c004c0030104400003000000000000001;
rom_uints[963] = 1024'h400000000000004301004c000100000100000000010c30004403003f0000000f0000140400070000c00044030000040000000c010cc00003011300000010000f4040000400001000004c0c00f301004c4300c300000000000301cc050101000c00c14004501100003400000d00300133000300100301000300c0c3050c0043c;
rom_uints[964] = 1024'h330c0404050330000001000000000300cc14434004c4040000d000300000000c500000401c040c01000000000404003000c15400040c040043300000004300000000000000000050000010c104010400031c00040000000000030430000c0c0001144003030400000c00c001c1400404000c0c00000c00000400010040030700;
rom_uints[965] = 1024'h4000c000000000010031c100c00000000000010000000001c000000143040300000010c33040030003010000000100000000000340100000c00300000000000300100000000100000044c000000000000000004000c00003010303000000c40000000040000000000000000030000001c00300c0000000000043030003010;
rom_uints[966] = 1024'h311000c0c000003001343c000030000c00000430500400c000000013003c000c40403c000c0000030004c0000000000034c0310000300010c00000000014040000000004300c40040cf0100c000000000000000000040000c0004014000c000000000040300030d000cc0000000004c4003000103c041c0000004010000;
rom_uints[967] = 1024'hc00000000400000d00c0000000000003000300030030000301d000030c00111003010c000000000000000000030040400030000010000030001010000000030001003000c14000000000000040000400000000030c000000000000004000011000001010004003000000010000000000700000000000000000030000;
rom_uints[968] = 1024'h10000403030300000000000300f001400000001003100030013531040c0c100000000000000000001000000005000030000000100410100000000000003000101013003000000030000001000c0000000000300010000010000000000400000000000c034300300c00300d004000040000000c0000100000001000000104003;
rom_uints[969] = 1024'h304003000c0000000100040014400d00400040004000c0c04c0c0fc000000101400000f3000000000000c00c000300000003010001c340040c000000040000c040000301030140c000000400034000400000000c00c0c00c00030c4c0000000003000cc003c00000000000000030000000400000000400c000;
rom_uints[970] = 1024'h100c0c10000000030c0001c431000c100c00000000000010000000000104000000000103010300c47403c0000c00000000000440000500000001000f0000000100100100000f00030004004000000c00000c00400c0010410000014300c0040000c4010104451004c004000c0100000c001c400c000034000000c000c003;
rom_uints[971] = 1024'h100004c00000000000010040c00c013003300011c000000040c044300c0c30f133c3000011c000007000100030400cd4c0040000010f30000c003100c4000400f0400000c0000400001c300300000c40f3000000000300400c0400441303c000170153000300000030000100000c3030000000300100c00004000000000050c;
rom_uints[972] = 1024'h3004300000300000010030000030f0000000300c10c0000000300000c03030c10000700000000000c01030100010c0043000c0001000000003c000c00000000040013001f00400c00340c010f00000003000000000001000c00000c00030000051000000000000010000001000013000000000f000000000100000000001000;
rom_uints[973] = 1024'h3c000000004000100030103000c00100c043001030440300f04000400000000001c0003c30100000c0310000400000301033000030d000340301300310103000c0c0000000010043000001d040c040000000040000030000003000000030c000c00000c00c004cc0c010000000000000000000f03000000010000f00f0d04000;
rom_uints[974] = 1024'h3000c00000000000000000000040000000000040403000000000001000303000001000300030000040d000000003000000000000000000004000c04000000000d3000000000000403000000000300c00000000100000100000001000000000000000003000000040000000000040000000000000100000000300000000000000;
rom_uints[975] = 1024'h3000040000007100007000014000300000c0440704300c00300000004000001000c0c00040300003000000000010310010000000000c000f0c00000000d300300000103c0c04040003c14000c00040c000000000000000004010400030001c40103000000001001030414040000000000000000c400000000000000004000;
rom_uints[976] = 1024'hc00031000000000000c0030000d0050c40000400000c0301000403100401001000400000000c0c000000007000000000100000000d0cc000001300030000c015000000d0000000000000c0cc400000000000c00030cc030400005c4000430c01140000000000000000000000000000000000400c000c000003000c0;
rom_uints[977] = 1024'h1000011c400100000000000000000000000003000010100c0014000000c030000c0000000004c0000111000c0001000000000100400c03000001c0013f30100000004100fc00010303000000000000310431000000c00000000c0000101000010300300c000000400000040300000004000d01000000040000010d000c00000f;
rom_uints[978] = 1024'hc000400000300000c000000010000003000300c0c1010000010000c0f03003030110000143030000030000000000000100000301400000000000c0000000c000c0000000000300000004c000c000c003000301404000c0130140c0000000030343100001000041c03003000000c04000004100000000000304004000c040;
rom_uints[979] = 1024'hc03000300c3000330004c00440000400001100004000c03030000003000c0c5040000000003030403030c000001000305100500000030c010030000000d00000f3000000300440d0c0000000400030000000c000300030000000401000c044410044000104000040000000000010000000000400003040000040400000100000;
rom_uints[980] = 1024'h1300000000000f0000000000000004040c001104001403000000000000040c000441000001000000000030010003000c101400c000000000300c000c00000000000c040c1000000000300c0000000030c000c0000000c00c04000000040000000000440000000c00000300000000000040000000000c0c0c03040300;
rom_uints[981] = 1024'h310010010000030000010000000c000000030000000101010000000100001000130000000301000010300300000000010003000000100100000101000000000004000003100100000000000300000000000000030000000000000000000000010000000100000000000100030000000000000000030000001000030000000700;
rom_uints[982] = 1024'h103000ccc014000c40d000c40400000c0c50000004013000000400400004001033103301017c14000400000000f00000000000c000d00000300010c0000000100000000000000010000c000c0430000000000c40040001000004000000000000000400001c000000003000010c100000c030003000000000000000000400110c;
rom_uints[983] = 1024'h70000000300030c0000000000000000003300000000000000000000000000040000000000010f0000300000000003030000000000000130000000000000000100011000c004000000000000000000000000000c0000010000000700004c00010000000000000000000030000400000000040000010000000000100000;
rom_uints[984] = 1024'h50c0c014300000c00000400d00000000c000c01000000000401000004030103030f0c0404000003044f0001000c04000000400013000000000500000f0c0004005400040400031c00000400000700340c000400000000040c3d030c000d000c04000410170000300400000c0f040300300c043c00000c000000030c0c040;
rom_uints[985] = 1024'h300c0000000400000150001000010010000001c00000030004040000f0000030cc0000000c0030000c00000400300010000010100000c0c0000000d430000c00000030303000000010043000100000100010100000000c00001003300000000400000000000010300000000100100000003c003000000000403041001100;
rom_uints[986] = 1024'hc0030000000000000000000041000000004000c010c0c040cc400000003300400000c000000040004000000000000000000000c0010000c000c00000c040c04000c0c00000000014c00000300000c1c000000040c000000000000040c000000000000000003000000030000000c0c0c010000f4000010000000000004040004;
rom_uints[987] = 1024'h1000000010001000000c3430003000000400100000040000005000d00c1030000000c0f050dc00404031000000000c00000000000c0000000100000001340000000400000000040010004c00003000010000100000c000000000000000c0300000410430003010000000000000300dc01030000000100000300000000c00400;
rom_uints[988] = 1024'hc000000c0c00040004c4000c000c040104000000000c0c000c0004000c00030d0004040c000f400400301000000000c0004400000cd00c00040f000000300c01100c0c04000000000c04000c000c3404000004000004000000000c0c000400000001400c050c400c00c0041004010000300c000c400000000330000001000103;
rom_uints[989] = 1024'h400000000c33010000100300330400100000cd0c004003003c0004000310500010130100000000100000000000700000010001c000c0103030300010001001000010000000c100000000100000300003000130000000040003004c0c100000500000430010000004c0c00000000000000010037100413000000040000c0;
rom_uints[990] = 1024'h100000000c0040000100000100c0000400004c0070000000044000cc0013040040340041004c01007000000000000010040000000040000000000000004043000400c000c013010000000040c0c047004000c0000000000000000040400000100000d400c0000043000000000000000000100000000000000c000000004c;
rom_uints[991] = 1024'h4000044c00010c000050000003000000100400c530000c0c000c0c10003400001000001000000030400c00000c0c001030003407030000013000040400030003000040004c01100000043c0010000030003000000c304c40000000000000300000000004400000000000350000300c004030010cc0000cc3000040300000;
rom_uints[992] = 1024'hc0000070700000c00000c0000000000000c0c000000030400000003000c000404000000000000000130000000000c000c0100000000040000000041030004040000000000000c0c000004000000000000000000000000000000000000000000000400000c000000000007000004000004000c0410000c000400000004000400;
rom_uints[993] = 1024'h1000c4400004030000001c3000000000101c001404040400040c043c0c1c000c00000000000c0400133c000400c00400000400004c00000001000c0000000c000c311c3000000000003000043030001c0c000310100400000cd4001004003000001c0c001030000c300000010010440c00000c3c04000c000400033c0000100;
rom_uints[994] = 1024'hc000000000040000000000100c0100000000000010033000000000030000010000004000000405030140000000000000000000004013004c0001000100000003000000000100010f100000000c40300000010000000000000005000300000000000311010001000000030000000000000000000c000400030300000000000301;
rom_uints[995] = 1024'h30000000003000000000300000000000000000000000001000004430300000000000000400000030000000000000000300000000001c00000000000000400000000000470000c0000010000000000040000000000000000000304000003c000430000000001000000400000000104000300040000030000000011000430000;
rom_uints[996] = 1024'hd030310000000000000000003130010000500001100000000000d000100300003000000000100010004000030000000000003c00c0c000130f0030c00000000000003010000000440000300000000040000000000000100000c0000000000031005000000000c030003031004000000000300040000c300000003000100000;
rom_uints[997] = 1024'h10300c3404300001004003100000000000c00400003004073000000c00103c0010403000c10c000000000007040f0001303013403c101000000c0c03010001000400000c0000000030000c00300c00000030000c010c740000000010003010305c1004300c07000030000c000004100000000c0000000000103404003;
rom_uints[998] = 1024'h4000000000000c0f000100040300000104000130010f000c000c0540014c000f00000000000c1100410c000000030004c00f0000030001040300030000000f0005000000003101000003000000000c01000103000000011400110300cc005300040030300000000300004001030000030000000003000303000000000003;
rom_uints[999] = 1024'hcd00400301000300013c01000304100000000100010003300f00000000004030400300010331000c400010000030c0010013000c00013000c000f0000110004003005000403033040510000003001000000300000003000000000000030000000001010000000000000103000001c0030300033300000000c0000c7300001000;
rom_uints[1000] = 1024'h40cc00c0000040004003c000040cc003050400000c100300000c00c0000000c00d00c4cc100c4003c0010c0000030c0000c70005040c0003d000000001c04000440100cc00c400000000000c410c00c100004000004c0000000000cc031000000000c03001c401c043cc0c00f00003000000c0c0040003004c0c0000c00f0c;
rom_uints[1001] = 1024'hc00400000f0300c4000304000370c00100000300000cc00d000c4040c004c400000010000c0cc40001c00000043c400cc0430f034000010000c101000c000010c407000304000003c00c044c000001040047000044004001000400000010040c4c0c34400100000000030101400000000004030d000040400000000c00010100;
rom_uints[1002] = 1024'h4dc000000040000000001000c0c700140040000000004000300000000000001cc000410c00005040c403000300000000000c103c000300000100000730000010400040010100000c0100403400000000010000c0430100d0434000d000100000000003004000300030000c0000000000300000d0400103c0c000000010105030;
rom_uints[1003] = 1024'h1000004000000505010500c4050000000004d004044000403cc001003400000c003c40c0400400430400c000044001001004c3c0000c4cc100000041000001000c30c0010c00140000000043000000c0400001c0000300000c1031c0c0403000f00040000000f000004410cc0000c0c000100340000300040000004000;
rom_uints[1004] = 1024'hc00c0440000c000c00f0c0040005400000400000c000c00000004000000000004000430100100000004cc000404000004000c0c04000000000c00000000400000000c4000000000000000000444000c000000000100000004001100000c01000c000050400400000000c00c000004013000c0040000000000000c04000004100;
rom_uints[1005] = 1024'h110300c0000010401000101cc00000040c001010c700004040000c0c000400004010f0000000000000000300000c0000000017000004000033000003f40c0c1c00000d00040000c00044300000004010704000001010000000000000010c00401000c0000400000000044470000400cc0c0104110000003cf10030c00c040;
rom_uints[1006] = 1024'h100000000000303c3000000c000000000030301010000031000000001000000000000000000000000000103000000000c00010000000033000000000000000000000100000000000300010033030000300300001303000000000010000000000000310000000100000003000300000001000;
rom_uints[1007] = 1024'h3000c000000400000004300000000000343000000000301000000000003010000000000000103000100000001000000000000030003c0030000000000000000000101000300000000000000000000000000000000030000000000000000000c03000000000000000000030300000003000103000300000103410000c;
rom_uints[1008] = 1024'h400000000000cc00c4c00000400040000000c0000c000003000000c444c0000000000c000000f00030004000004000c000000000000000000400000300c000040000410000c00000000040004000003000000000c00000c00c00010010000004c000000000004000000000c0000000400000000000c000000000c0c00040;
rom_uints[1009] = 1024'h304c00004000430010100000000000dc104400040004303000000040001010000004000000c000c0010c000000404000c00000030000c00000000000d400c0000000000000000000c000000400000000000040004000c4000004003000dcc0004000000040000100000470004033010000c3000c000004000000000c00c07010;
rom_uints[1010] = 1024'h30000000000100c000004c0000000000000000c000f0000000c00000104d001004000c0000000000040000004000c04000000000000000000041004000c040000040010001000000000003c010030c01000000c04140000040414000003000000450010003c0c50000000000c00000000000010400010000000c000000000003;
rom_uints[1011] = 1024'hc010000030cc00000000c1003000d03110000030000c3000c00000403000000000000000700cd0100000300000400010001001000004000000c0f03000003000000030100000001000000040000000000010000000000000003400403000000004007100c000000001c010000000003000000030400000301000003000003300;
rom_uints[1012] = 1024'h1040000c00000000000000000000400010004000000000c00000003000000400400c00330000000003100000000400000140003300000000300000033000000000f00014400000000000000000000000000000000000000000000010000000000300000004000000000000000000030000000000000040000000000;
rom_uints[1013] = 1024'hc00000c00040010001000100d04000f0000000040001000c0300000000000400000000104040000000c1000000000000c071000000000000030000000000c000c00000003c30000004000403c0030000cc00400000000001c000400001c0004000c50003000003004013000040c000000c0c0ff400004300400000c000c0000;
rom_uints[1014] = 1024'hc4000430000000c400000000000c4003001000000cc0c400000000c0001c00104000000000030000104300000000d000003000004c004000c0c70001000c4000f0000010001000cc0000040c000000c0003000c1000010003000001000c30000014000001040001030000000113000000000004000000040001c004040003303;
rom_uints[1015] = 1024'h10003000100000c00004003070004400c13011000c0c1030000400000030000000c0005c0000000030700000300030003030300040100000c010000000000000c0111000f001000010000c100030c000000000000000000000dc0050100c0c4c10000004000c00004c1000100000301000300030100c1034000000000030003;
rom_uints[1016] = 1024'hc1c00001005000c300c0000c00030000030001c10111c000070044c10040000030c0400007410001033100000000000000000010010003010040010000000100c000070100003000003003001000000010400030103301003c000100c1c30003c040000d0043000750c3030301000003030000700000000003000040010103c;
rom_uints[1017] = 1024'hf000c00030c0300310003000000000300000c0404001040000d0000000c000000040007000dc0001003070000000000000001014004c00000000004030000000303000c0c0c000000f0000400000000000000004000000000040100000000110000030300000400001010040000300000010d0c000d000000000000030000300;
rom_uints[1018] = 1024'h400000000000400000000000000000000000000c00000000000000443c0100000400003030c0003004400000000000000c0000000c00c0000c0000000000000000000000000000404000300000000400040000000000000000c000000c00000000003000000004c0000040410000c00cc0040040000000000000000000000;
rom_uints[1019] = 1024'h40000040010040c04001030000c004c00000000140400000000050000003010070c00040000c40410c410000c101000300c000000000000030000000c00040000c00c000000301004000000003000000c000000103010000000000004003000c13000000000000c10300300000c000000c0010000000c00000400150004004;
rom_uints[1020] = 1024'h3000c0c0000c000000000000000000c0000000044030c0300100000000c00000004000c00003004c3000010000c0300cc000000d000000040000000000c00000410000100000000104000000030000000100000c000000000004000004400000500040c00400000010000000500c0400000000000100000c04034000000010c0;
rom_uints[1021] = 1024'h307c300c0000000000000000040000003130100000001000000007030000040c3000300000000010000004100c340000000030010010000000000030001030300010013000003c3000001000003d00300c0c0030000000000c00100f00001014000c300c04000c0030340030000c000000003c00000000030000003;
rom_uints[1022] = 1024'h1d041c13000d301000c00c300330003000300c00000c100013300000703c003430070c0000010c00303c1004030303001000001000000003331003000030030010100c005c0300310d14300400030001101c30331030030000000030100101000430010000004034300330070001000003100c30010300c00000000000000103;
rom_uints[1023] = 1024'h400000301000001c3050543001004c0c3031400c000c00100c0000c000000003c3003140011440000003000000300d0000103000001000c0310410001070000f44034000003c00011000001030003400004c004000c0000304000003001c30031c3430314430c001fc100010500030c0003400c000100030100010f4c0031c0;
end

reg [1023:0] outputReg;
assign out = outputReg;
always @(posedge clock)
begin
  outputReg <= rom_uints[readAddr];
end
endmodule
