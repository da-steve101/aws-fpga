module MuxLayer(
  input         clock,
  input         reset,
  output        io_dataIn_ready,
  input         io_dataIn_valid,
  input  [15:0] io_dataIn_bits_0,
  input  [15:0] io_dataIn_bits_1,
  input  [15:0] io_dataIn_bits_2,
  input  [15:0] io_dataIn_bits_3,
  input  [15:0] io_dataIn_bits_4,
  input  [15:0] io_dataIn_bits_5,
  input  [15:0] io_dataIn_bits_6,
  input  [15:0] io_dataIn_bits_7,
  input  [15:0] io_dataIn_bits_8,
  input  [15:0] io_dataIn_bits_9,
  input  [15:0] io_dataIn_bits_10,
  input  [15:0] io_dataIn_bits_11,
  input  [15:0] io_dataIn_bits_12,
  input  [15:0] io_dataIn_bits_13,
  input  [15:0] io_dataIn_bits_14,
  input  [15:0] io_dataIn_bits_15,
  input  [15:0] io_dataIn_bits_16,
  input  [15:0] io_dataIn_bits_17,
  input  [15:0] io_dataIn_bits_18,
  input  [15:0] io_dataIn_bits_19,
  input  [15:0] io_dataIn_bits_20,
  input  [15:0] io_dataIn_bits_21,
  input  [15:0] io_dataIn_bits_22,
  input  [15:0] io_dataIn_bits_23,
  input  [15:0] io_dataIn_bits_24,
  input  [15:0] io_dataIn_bits_25,
  input  [15:0] io_dataIn_bits_26,
  input  [15:0] io_dataIn_bits_27,
  input  [15:0] io_dataIn_bits_28,
  input  [15:0] io_dataIn_bits_29,
  input  [15:0] io_dataIn_bits_30,
  input  [15:0] io_dataIn_bits_31,
  input  [15:0] io_dataIn_bits_32,
  input  [15:0] io_dataIn_bits_33,
  input  [15:0] io_dataIn_bits_34,
  input  [15:0] io_dataIn_bits_35,
  input  [15:0] io_dataIn_bits_36,
  input  [15:0] io_dataIn_bits_37,
  input  [15:0] io_dataIn_bits_38,
  input  [15:0] io_dataIn_bits_39,
  input  [15:0] io_dataIn_bits_40,
  input  [15:0] io_dataIn_bits_41,
  input  [15:0] io_dataIn_bits_42,
  input  [15:0] io_dataIn_bits_43,
  input  [15:0] io_dataIn_bits_44,
  input  [15:0] io_dataIn_bits_45,
  input  [15:0] io_dataIn_bits_46,
  input  [15:0] io_dataIn_bits_47,
  input  [15:0] io_dataIn_bits_48,
  input  [15:0] io_dataIn_bits_49,
  input  [15:0] io_dataIn_bits_50,
  input  [15:0] io_dataIn_bits_51,
  input  [15:0] io_dataIn_bits_52,
  input  [15:0] io_dataIn_bits_53,
  input  [15:0] io_dataIn_bits_54,
  input  [15:0] io_dataIn_bits_55,
  input  [15:0] io_dataIn_bits_56,
  input  [15:0] io_dataIn_bits_57,
  input  [15:0] io_dataIn_bits_58,
  input  [15:0] io_dataIn_bits_59,
  input  [15:0] io_dataIn_bits_60,
  input  [15:0] io_dataIn_bits_61,
  input  [15:0] io_dataIn_bits_62,
  input  [15:0] io_dataIn_bits_63,
  input  [15:0] io_dataIn_bits_64,
  input  [15:0] io_dataIn_bits_65,
  input  [15:0] io_dataIn_bits_66,
  input  [15:0] io_dataIn_bits_67,
  input  [15:0] io_dataIn_bits_68,
  input  [15:0] io_dataIn_bits_69,
  input  [15:0] io_dataIn_bits_70,
  input  [15:0] io_dataIn_bits_71,
  input  [15:0] io_dataIn_bits_72,
  input  [15:0] io_dataIn_bits_73,
  input  [15:0] io_dataIn_bits_74,
  input  [15:0] io_dataIn_bits_75,
  input  [15:0] io_dataIn_bits_76,
  input  [15:0] io_dataIn_bits_77,
  input  [15:0] io_dataIn_bits_78,
  input  [15:0] io_dataIn_bits_79,
  input  [15:0] io_dataIn_bits_80,
  input  [15:0] io_dataIn_bits_81,
  input  [15:0] io_dataIn_bits_82,
  input  [15:0] io_dataIn_bits_83,
  input  [15:0] io_dataIn_bits_84,
  input  [15:0] io_dataIn_bits_85,
  input  [15:0] io_dataIn_bits_86,
  input  [15:0] io_dataIn_bits_87,
  input  [15:0] io_dataIn_bits_88,
  input  [15:0] io_dataIn_bits_89,
  input  [15:0] io_dataIn_bits_90,
  input  [15:0] io_dataIn_bits_91,
  input  [15:0] io_dataIn_bits_92,
  input  [15:0] io_dataIn_bits_93,
  input  [15:0] io_dataIn_bits_94,
  input  [15:0] io_dataIn_bits_95,
  input  [15:0] io_dataIn_bits_96,
  input  [15:0] io_dataIn_bits_97,
  input  [15:0] io_dataIn_bits_98,
  input  [15:0] io_dataIn_bits_99,
  input  [15:0] io_dataIn_bits_100,
  input  [15:0] io_dataIn_bits_101,
  input  [15:0] io_dataIn_bits_102,
  input  [15:0] io_dataIn_bits_103,
  input  [15:0] io_dataIn_bits_104,
  input  [15:0] io_dataIn_bits_105,
  input  [15:0] io_dataIn_bits_106,
  input  [15:0] io_dataIn_bits_107,
  input  [15:0] io_dataIn_bits_108,
  input  [15:0] io_dataIn_bits_109,
  input  [15:0] io_dataIn_bits_110,
  input  [15:0] io_dataIn_bits_111,
  input  [15:0] io_dataIn_bits_112,
  input  [15:0] io_dataIn_bits_113,
  input  [15:0] io_dataIn_bits_114,
  input  [15:0] io_dataIn_bits_115,
  input  [15:0] io_dataIn_bits_116,
  input  [15:0] io_dataIn_bits_117,
  input  [15:0] io_dataIn_bits_118,
  input  [15:0] io_dataIn_bits_119,
  input  [15:0] io_dataIn_bits_120,
  input  [15:0] io_dataIn_bits_121,
  input  [15:0] io_dataIn_bits_122,
  input  [15:0] io_dataIn_bits_123,
  input  [15:0] io_dataIn_bits_124,
  input  [15:0] io_dataIn_bits_125,
  input  [15:0] io_dataIn_bits_126,
  input  [15:0] io_dataIn_bits_127,
  input  [15:0] io_dataIn_bits_128,
  input  [15:0] io_dataIn_bits_129,
  input  [15:0] io_dataIn_bits_130,
  input  [15:0] io_dataIn_bits_131,
  input  [15:0] io_dataIn_bits_132,
  input  [15:0] io_dataIn_bits_133,
  input  [15:0] io_dataIn_bits_134,
  input  [15:0] io_dataIn_bits_135,
  input  [15:0] io_dataIn_bits_136,
  input  [15:0] io_dataIn_bits_137,
  input  [15:0] io_dataIn_bits_138,
  input  [15:0] io_dataIn_bits_139,
  input  [15:0] io_dataIn_bits_140,
  input  [15:0] io_dataIn_bits_141,
  input  [15:0] io_dataIn_bits_142,
  input  [15:0] io_dataIn_bits_143,
  input  [15:0] io_dataIn_bits_144,
  input  [15:0] io_dataIn_bits_145,
  input  [15:0] io_dataIn_bits_146,
  input  [15:0] io_dataIn_bits_147,
  input  [15:0] io_dataIn_bits_148,
  input  [15:0] io_dataIn_bits_149,
  input  [15:0] io_dataIn_bits_150,
  input  [15:0] io_dataIn_bits_151,
  input  [15:0] io_dataIn_bits_152,
  input  [15:0] io_dataIn_bits_153,
  input  [15:0] io_dataIn_bits_154,
  input  [15:0] io_dataIn_bits_155,
  input  [15:0] io_dataIn_bits_156,
  input  [15:0] io_dataIn_bits_157,
  input  [15:0] io_dataIn_bits_158,
  input  [15:0] io_dataIn_bits_159,
  input  [15:0] io_dataIn_bits_160,
  input  [15:0] io_dataIn_bits_161,
  input  [15:0] io_dataIn_bits_162,
  input  [15:0] io_dataIn_bits_163,
  input  [15:0] io_dataIn_bits_164,
  input  [15:0] io_dataIn_bits_165,
  input  [15:0] io_dataIn_bits_166,
  input  [15:0] io_dataIn_bits_167,
  input  [15:0] io_dataIn_bits_168,
  input  [15:0] io_dataIn_bits_169,
  input  [15:0] io_dataIn_bits_170,
  input  [15:0] io_dataIn_bits_171,
  input  [15:0] io_dataIn_bits_172,
  input  [15:0] io_dataIn_bits_173,
  input  [15:0] io_dataIn_bits_174,
  input  [15:0] io_dataIn_bits_175,
  input  [15:0] io_dataIn_bits_176,
  input  [15:0] io_dataIn_bits_177,
  input  [15:0] io_dataIn_bits_178,
  input  [15:0] io_dataIn_bits_179,
  input  [15:0] io_dataIn_bits_180,
  input  [15:0] io_dataIn_bits_181,
  input  [15:0] io_dataIn_bits_182,
  input  [15:0] io_dataIn_bits_183,
  input  [15:0] io_dataIn_bits_184,
  input  [15:0] io_dataIn_bits_185,
  input  [15:0] io_dataIn_bits_186,
  input  [15:0] io_dataIn_bits_187,
  input  [15:0] io_dataIn_bits_188,
  input  [15:0] io_dataIn_bits_189,
  input  [15:0] io_dataIn_bits_190,
  input  [15:0] io_dataIn_bits_191,
  input  [15:0] io_dataIn_bits_192,
  input  [15:0] io_dataIn_bits_193,
  input  [15:0] io_dataIn_bits_194,
  input  [15:0] io_dataIn_bits_195,
  input  [15:0] io_dataIn_bits_196,
  input  [15:0] io_dataIn_bits_197,
  input  [15:0] io_dataIn_bits_198,
  input  [15:0] io_dataIn_bits_199,
  input  [15:0] io_dataIn_bits_200,
  input  [15:0] io_dataIn_bits_201,
  input  [15:0] io_dataIn_bits_202,
  input  [15:0] io_dataIn_bits_203,
  input  [15:0] io_dataIn_bits_204,
  input  [15:0] io_dataIn_bits_205,
  input  [15:0] io_dataIn_bits_206,
  input  [15:0] io_dataIn_bits_207,
  input  [15:0] io_dataIn_bits_208,
  input  [15:0] io_dataIn_bits_209,
  input  [15:0] io_dataIn_bits_210,
  input  [15:0] io_dataIn_bits_211,
  input  [15:0] io_dataIn_bits_212,
  input  [15:0] io_dataIn_bits_213,
  input  [15:0] io_dataIn_bits_214,
  input  [15:0] io_dataIn_bits_215,
  input  [15:0] io_dataIn_bits_216,
  input  [15:0] io_dataIn_bits_217,
  input  [15:0] io_dataIn_bits_218,
  input  [15:0] io_dataIn_bits_219,
  input  [15:0] io_dataIn_bits_220,
  input  [15:0] io_dataIn_bits_221,
  input  [15:0] io_dataIn_bits_222,
  input  [15:0] io_dataIn_bits_223,
  input  [15:0] io_dataIn_bits_224,
  input  [15:0] io_dataIn_bits_225,
  input  [15:0] io_dataIn_bits_226,
  input  [15:0] io_dataIn_bits_227,
  input  [15:0] io_dataIn_bits_228,
  input  [15:0] io_dataIn_bits_229,
  input  [15:0] io_dataIn_bits_230,
  input  [15:0] io_dataIn_bits_231,
  input  [15:0] io_dataIn_bits_232,
  input  [15:0] io_dataIn_bits_233,
  input  [15:0] io_dataIn_bits_234,
  input  [15:0] io_dataIn_bits_235,
  input  [15:0] io_dataIn_bits_236,
  input  [15:0] io_dataIn_bits_237,
  input  [15:0] io_dataIn_bits_238,
  input  [15:0] io_dataIn_bits_239,
  input  [15:0] io_dataIn_bits_240,
  input  [15:0] io_dataIn_bits_241,
  input  [15:0] io_dataIn_bits_242,
  input  [15:0] io_dataIn_bits_243,
  input  [15:0] io_dataIn_bits_244,
  input  [15:0] io_dataIn_bits_245,
  input  [15:0] io_dataIn_bits_246,
  input  [15:0] io_dataIn_bits_247,
  input  [15:0] io_dataIn_bits_248,
  input  [15:0] io_dataIn_bits_249,
  input  [15:0] io_dataIn_bits_250,
  input  [15:0] io_dataIn_bits_251,
  input  [15:0] io_dataIn_bits_252,
  input  [15:0] io_dataIn_bits_253,
  input  [15:0] io_dataIn_bits_254,
  input  [15:0] io_dataIn_bits_255,
  output        io_dataOut_valid,
  output [15:0] io_dataOut_bits_0,
  output [15:0] io_dataOut_bits_1,
  output [15:0] io_dataOut_bits_2,
  output [15:0] io_dataOut_bits_3
);
  reg  rdyReg; // @[MuxLayer.scala 14:23]
  reg [31:0] _RAND_0;
  reg [5:0] cntr; // @[MuxLayer.scala 17:21]
  reg [31:0] _RAND_1;
  reg [15:0] buffers_0_0_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_2;
  reg [15:0] buffers_0_0_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_3;
  reg [15:0] buffers_0_0_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_4;
  reg [15:0] buffers_0_0_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_5;
  reg [15:0] buffers_0_1_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_6;
  reg [15:0] buffers_0_1_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_7;
  reg [15:0] buffers_0_1_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_8;
  reg [15:0] buffers_0_1_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_9;
  reg [15:0] buffers_0_2_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_10;
  reg [15:0] buffers_0_2_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_11;
  reg [15:0] buffers_0_2_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_12;
  reg [15:0] buffers_0_2_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_13;
  reg [15:0] buffers_0_3_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_14;
  reg [15:0] buffers_0_3_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_15;
  reg [15:0] buffers_0_3_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_16;
  reg [15:0] buffers_0_3_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_17;
  reg [15:0] buffers_0_4_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_18;
  reg [15:0] buffers_0_4_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_19;
  reg [15:0] buffers_0_4_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_20;
  reg [15:0] buffers_0_4_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_21;
  reg [15:0] buffers_0_5_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_22;
  reg [15:0] buffers_0_5_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_23;
  reg [15:0] buffers_0_5_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_24;
  reg [15:0] buffers_0_5_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_25;
  reg [15:0] buffers_0_6_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_26;
  reg [15:0] buffers_0_6_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_27;
  reg [15:0] buffers_0_6_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_28;
  reg [15:0] buffers_0_6_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_29;
  reg [15:0] buffers_0_7_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_30;
  reg [15:0] buffers_0_7_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_31;
  reg [15:0] buffers_0_7_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_32;
  reg [15:0] buffers_0_7_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_33;
  reg [15:0] buffers_0_8_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_34;
  reg [15:0] buffers_0_8_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_35;
  reg [15:0] buffers_0_8_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_36;
  reg [15:0] buffers_0_8_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_37;
  reg [15:0] buffers_0_9_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_38;
  reg [15:0] buffers_0_9_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_39;
  reg [15:0] buffers_0_9_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_40;
  reg [15:0] buffers_0_9_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_41;
  reg [15:0] buffers_0_10_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_42;
  reg [15:0] buffers_0_10_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_43;
  reg [15:0] buffers_0_10_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_44;
  reg [15:0] buffers_0_10_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_45;
  reg [15:0] buffers_0_11_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_46;
  reg [15:0] buffers_0_11_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_47;
  reg [15:0] buffers_0_11_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_48;
  reg [15:0] buffers_0_11_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_49;
  reg [15:0] buffers_0_12_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_50;
  reg [15:0] buffers_0_12_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_51;
  reg [15:0] buffers_0_12_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_52;
  reg [15:0] buffers_0_12_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_53;
  reg [15:0] buffers_0_13_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_54;
  reg [15:0] buffers_0_13_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_55;
  reg [15:0] buffers_0_13_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_56;
  reg [15:0] buffers_0_13_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_57;
  reg [15:0] buffers_0_14_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_58;
  reg [15:0] buffers_0_14_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_59;
  reg [15:0] buffers_0_14_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_60;
  reg [15:0] buffers_0_14_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_61;
  reg [15:0] buffers_0_15_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_62;
  reg [15:0] buffers_0_15_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_63;
  reg [15:0] buffers_0_15_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_64;
  reg [15:0] buffers_0_15_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_65;
  reg [15:0] buffers_0_16_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_66;
  reg [15:0] buffers_0_16_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_67;
  reg [15:0] buffers_0_16_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_68;
  reg [15:0] buffers_0_16_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_69;
  reg [15:0] buffers_0_17_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_70;
  reg [15:0] buffers_0_17_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_71;
  reg [15:0] buffers_0_17_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_72;
  reg [15:0] buffers_0_17_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_73;
  reg [15:0] buffers_0_18_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_74;
  reg [15:0] buffers_0_18_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_75;
  reg [15:0] buffers_0_18_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_76;
  reg [15:0] buffers_0_18_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_77;
  reg [15:0] buffers_0_19_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_78;
  reg [15:0] buffers_0_19_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_79;
  reg [15:0] buffers_0_19_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_80;
  reg [15:0] buffers_0_19_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_81;
  reg [15:0] buffers_0_20_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_82;
  reg [15:0] buffers_0_20_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_83;
  reg [15:0] buffers_0_20_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_84;
  reg [15:0] buffers_0_20_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_85;
  reg [15:0] buffers_0_21_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_86;
  reg [15:0] buffers_0_21_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_87;
  reg [15:0] buffers_0_21_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_88;
  reg [15:0] buffers_0_21_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_89;
  reg [15:0] buffers_0_22_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_90;
  reg [15:0] buffers_0_22_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_91;
  reg [15:0] buffers_0_22_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_92;
  reg [15:0] buffers_0_22_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_93;
  reg [15:0] buffers_0_23_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_94;
  reg [15:0] buffers_0_23_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_95;
  reg [15:0] buffers_0_23_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_96;
  reg [15:0] buffers_0_23_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_97;
  reg [15:0] buffers_0_24_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_98;
  reg [15:0] buffers_0_24_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_99;
  reg [15:0] buffers_0_24_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_100;
  reg [15:0] buffers_0_24_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_101;
  reg [15:0] buffers_0_25_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_102;
  reg [15:0] buffers_0_25_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_103;
  reg [15:0] buffers_0_25_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_104;
  reg [15:0] buffers_0_25_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_105;
  reg [15:0] buffers_0_26_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_106;
  reg [15:0] buffers_0_26_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_107;
  reg [15:0] buffers_0_26_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_108;
  reg [15:0] buffers_0_26_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_109;
  reg [15:0] buffers_0_27_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_110;
  reg [15:0] buffers_0_27_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_111;
  reg [15:0] buffers_0_27_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_112;
  reg [15:0] buffers_0_27_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_113;
  reg [15:0] buffers_0_28_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_114;
  reg [15:0] buffers_0_28_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_115;
  reg [15:0] buffers_0_28_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_116;
  reg [15:0] buffers_0_28_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_117;
  reg [15:0] buffers_0_29_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_118;
  reg [15:0] buffers_0_29_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_119;
  reg [15:0] buffers_0_29_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_120;
  reg [15:0] buffers_0_29_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_121;
  reg [15:0] buffers_0_30_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_122;
  reg [15:0] buffers_0_30_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_123;
  reg [15:0] buffers_0_30_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_124;
  reg [15:0] buffers_0_30_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_125;
  reg [15:0] buffers_0_31_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_126;
  reg [15:0] buffers_0_31_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_127;
  reg [15:0] buffers_0_31_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_128;
  reg [15:0] buffers_0_31_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_129;
  reg [15:0] buffers_0_32_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_130;
  reg [15:0] buffers_0_32_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_131;
  reg [15:0] buffers_0_32_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_132;
  reg [15:0] buffers_0_32_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_133;
  reg [15:0] buffers_0_33_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_134;
  reg [15:0] buffers_0_33_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_135;
  reg [15:0] buffers_0_33_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_136;
  reg [15:0] buffers_0_33_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_137;
  reg [15:0] buffers_0_34_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_138;
  reg [15:0] buffers_0_34_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_139;
  reg [15:0] buffers_0_34_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_140;
  reg [15:0] buffers_0_34_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_141;
  reg [15:0] buffers_0_35_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_142;
  reg [15:0] buffers_0_35_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_143;
  reg [15:0] buffers_0_35_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_144;
  reg [15:0] buffers_0_35_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_145;
  reg [15:0] buffers_0_36_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_146;
  reg [15:0] buffers_0_36_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_147;
  reg [15:0] buffers_0_36_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_148;
  reg [15:0] buffers_0_36_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_149;
  reg [15:0] buffers_0_37_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_150;
  reg [15:0] buffers_0_37_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_151;
  reg [15:0] buffers_0_37_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_152;
  reg [15:0] buffers_0_37_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_153;
  reg [15:0] buffers_0_38_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_154;
  reg [15:0] buffers_0_38_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_155;
  reg [15:0] buffers_0_38_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_156;
  reg [15:0] buffers_0_38_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_157;
  reg [15:0] buffers_0_39_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_158;
  reg [15:0] buffers_0_39_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_159;
  reg [15:0] buffers_0_39_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_160;
  reg [15:0] buffers_0_39_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_161;
  reg [15:0] buffers_0_40_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_162;
  reg [15:0] buffers_0_40_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_163;
  reg [15:0] buffers_0_40_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_164;
  reg [15:0] buffers_0_40_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_165;
  reg [15:0] buffers_0_41_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_166;
  reg [15:0] buffers_0_41_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_167;
  reg [15:0] buffers_0_41_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_168;
  reg [15:0] buffers_0_41_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_169;
  reg [15:0] buffers_0_42_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_170;
  reg [15:0] buffers_0_42_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_171;
  reg [15:0] buffers_0_42_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_172;
  reg [15:0] buffers_0_42_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_173;
  reg [15:0] buffers_0_43_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_174;
  reg [15:0] buffers_0_43_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_175;
  reg [15:0] buffers_0_43_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_176;
  reg [15:0] buffers_0_43_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_177;
  reg [15:0] buffers_0_44_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_178;
  reg [15:0] buffers_0_44_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_179;
  reg [15:0] buffers_0_44_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_180;
  reg [15:0] buffers_0_44_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_181;
  reg [15:0] buffers_0_45_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_182;
  reg [15:0] buffers_0_45_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_183;
  reg [15:0] buffers_0_45_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_184;
  reg [15:0] buffers_0_45_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_185;
  reg [15:0] buffers_0_46_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_186;
  reg [15:0] buffers_0_46_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_187;
  reg [15:0] buffers_0_46_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_188;
  reg [15:0] buffers_0_46_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_189;
  reg [15:0] buffers_0_47_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_190;
  reg [15:0] buffers_0_47_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_191;
  reg [15:0] buffers_0_47_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_192;
  reg [15:0] buffers_0_47_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_193;
  reg [15:0] buffers_0_48_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_194;
  reg [15:0] buffers_0_48_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_195;
  reg [15:0] buffers_0_48_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_196;
  reg [15:0] buffers_0_48_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_197;
  reg [15:0] buffers_0_49_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_198;
  reg [15:0] buffers_0_49_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_199;
  reg [15:0] buffers_0_49_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_200;
  reg [15:0] buffers_0_49_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_201;
  reg [15:0] buffers_0_50_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_202;
  reg [15:0] buffers_0_50_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_203;
  reg [15:0] buffers_0_50_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_204;
  reg [15:0] buffers_0_50_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_205;
  reg [15:0] buffers_0_51_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_206;
  reg [15:0] buffers_0_51_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_207;
  reg [15:0] buffers_0_51_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_208;
  reg [15:0] buffers_0_51_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_209;
  reg [15:0] buffers_0_52_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_210;
  reg [15:0] buffers_0_52_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_211;
  reg [15:0] buffers_0_52_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_212;
  reg [15:0] buffers_0_52_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_213;
  reg [15:0] buffers_0_53_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_214;
  reg [15:0] buffers_0_53_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_215;
  reg [15:0] buffers_0_53_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_216;
  reg [15:0] buffers_0_53_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_217;
  reg [15:0] buffers_0_54_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_218;
  reg [15:0] buffers_0_54_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_219;
  reg [15:0] buffers_0_54_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_220;
  reg [15:0] buffers_0_54_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_221;
  reg [15:0] buffers_0_55_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_222;
  reg [15:0] buffers_0_55_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_223;
  reg [15:0] buffers_0_55_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_224;
  reg [15:0] buffers_0_55_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_225;
  reg [15:0] buffers_0_56_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_226;
  reg [15:0] buffers_0_56_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_227;
  reg [15:0] buffers_0_56_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_228;
  reg [15:0] buffers_0_56_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_229;
  reg [15:0] buffers_0_57_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_230;
  reg [15:0] buffers_0_57_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_231;
  reg [15:0] buffers_0_57_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_232;
  reg [15:0] buffers_0_57_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_233;
  reg [15:0] buffers_0_58_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_234;
  reg [15:0] buffers_0_58_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_235;
  reg [15:0] buffers_0_58_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_236;
  reg [15:0] buffers_0_58_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_237;
  reg [15:0] buffers_0_59_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_238;
  reg [15:0] buffers_0_59_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_239;
  reg [15:0] buffers_0_59_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_240;
  reg [15:0] buffers_0_59_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_241;
  reg [15:0] buffers_0_60_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_242;
  reg [15:0] buffers_0_60_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_243;
  reg [15:0] buffers_0_60_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_244;
  reg [15:0] buffers_0_60_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_245;
  reg [15:0] buffers_0_61_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_246;
  reg [15:0] buffers_0_61_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_247;
  reg [15:0] buffers_0_61_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_248;
  reg [15:0] buffers_0_61_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_249;
  reg [15:0] buffers_0_62_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_250;
  reg [15:0] buffers_0_62_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_251;
  reg [15:0] buffers_0_62_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_252;
  reg [15:0] buffers_0_62_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_253;
  reg [15:0] buffers_0_63_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_254;
  reg [15:0] buffers_0_63_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_255;
  reg [15:0] buffers_0_63_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_256;
  reg [15:0] buffers_0_63_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_257;
  reg [1:0] cntrs_0; // @[Reg.scala 11:16]
  reg [31:0] _RAND_258;
  reg [1:0] _T_1071; // @[Reg.scala 11:16]
  reg [31:0] _RAND_259;
  reg [1:0] cntrs_1; // @[Reg.scala 11:16]
  reg [31:0] _RAND_260;
  reg [1:0] _T_1076; // @[Reg.scala 11:16]
  reg [31:0] _RAND_261;
  reg [1:0] _T_1078; // @[Reg.scala 11:16]
  reg [31:0] _RAND_262;
  reg [1:0] cntrs_2; // @[Reg.scala 11:16]
  reg [31:0] _RAND_263;
  reg [15:0] buffers_1_0_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_264;
  reg [15:0] buffers_1_0_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_265;
  reg [15:0] buffers_1_0_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_266;
  reg [15:0] buffers_1_0_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_267;
  reg [15:0] buffers_1_1_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_268;
  reg [15:0] buffers_1_1_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_269;
  reg [15:0] buffers_1_1_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_270;
  reg [15:0] buffers_1_1_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_271;
  reg [15:0] buffers_1_2_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_272;
  reg [15:0] buffers_1_2_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_273;
  reg [15:0] buffers_1_2_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_274;
  reg [15:0] buffers_1_2_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_275;
  reg [15:0] buffers_1_3_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_276;
  reg [15:0] buffers_1_3_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_277;
  reg [15:0] buffers_1_3_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_278;
  reg [15:0] buffers_1_3_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_279;
  reg [15:0] buffers_1_4_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_280;
  reg [15:0] buffers_1_4_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_281;
  reg [15:0] buffers_1_4_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_282;
  reg [15:0] buffers_1_4_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_283;
  reg [15:0] buffers_1_5_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_284;
  reg [15:0] buffers_1_5_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_285;
  reg [15:0] buffers_1_5_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_286;
  reg [15:0] buffers_1_5_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_287;
  reg [15:0] buffers_1_6_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_288;
  reg [15:0] buffers_1_6_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_289;
  reg [15:0] buffers_1_6_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_290;
  reg [15:0] buffers_1_6_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_291;
  reg [15:0] buffers_1_7_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_292;
  reg [15:0] buffers_1_7_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_293;
  reg [15:0] buffers_1_7_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_294;
  reg [15:0] buffers_1_7_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_295;
  reg [15:0] buffers_1_8_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_296;
  reg [15:0] buffers_1_8_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_297;
  reg [15:0] buffers_1_8_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_298;
  reg [15:0] buffers_1_8_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_299;
  reg [15:0] buffers_1_9_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_300;
  reg [15:0] buffers_1_9_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_301;
  reg [15:0] buffers_1_9_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_302;
  reg [15:0] buffers_1_9_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_303;
  reg [15:0] buffers_1_10_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_304;
  reg [15:0] buffers_1_10_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_305;
  reg [15:0] buffers_1_10_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_306;
  reg [15:0] buffers_1_10_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_307;
  reg [15:0] buffers_1_11_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_308;
  reg [15:0] buffers_1_11_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_309;
  reg [15:0] buffers_1_11_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_310;
  reg [15:0] buffers_1_11_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_311;
  reg [15:0] buffers_1_12_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_312;
  reg [15:0] buffers_1_12_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_313;
  reg [15:0] buffers_1_12_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_314;
  reg [15:0] buffers_1_12_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_315;
  reg [15:0] buffers_1_13_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_316;
  reg [15:0] buffers_1_13_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_317;
  reg [15:0] buffers_1_13_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_318;
  reg [15:0] buffers_1_13_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_319;
  reg [15:0] buffers_1_14_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_320;
  reg [15:0] buffers_1_14_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_321;
  reg [15:0] buffers_1_14_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_322;
  reg [15:0] buffers_1_14_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_323;
  reg [15:0] buffers_1_15_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_324;
  reg [15:0] buffers_1_15_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_325;
  reg [15:0] buffers_1_15_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_326;
  reg [15:0] buffers_1_15_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_327;
  reg [15:0] buffers_2_0_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_328;
  reg [15:0] buffers_2_0_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_329;
  reg [15:0] buffers_2_0_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_330;
  reg [15:0] buffers_2_0_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_331;
  reg [15:0] buffers_2_1_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_332;
  reg [15:0] buffers_2_1_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_333;
  reg [15:0] buffers_2_1_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_334;
  reg [15:0] buffers_2_1_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_335;
  reg [15:0] buffers_2_2_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_336;
  reg [15:0] buffers_2_2_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_337;
  reg [15:0] buffers_2_2_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_338;
  reg [15:0] buffers_2_2_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_339;
  reg [15:0] buffers_2_3_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_340;
  reg [15:0] buffers_2_3_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_341;
  reg [15:0] buffers_2_3_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_342;
  reg [15:0] buffers_2_3_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_343;
  reg [15:0] buffers_3_0_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_344;
  reg [15:0] buffers_3_0_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_345;
  reg [15:0] buffers_3_0_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_346;
  reg [15:0] buffers_3_0_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_347;
  reg  _T_1988; // @[Reg.scala 19:20]
  reg [31:0] _RAND_348;
  reg  _T_1990; // @[Reg.scala 19:20]
  reg [31:0] _RAND_349;
  reg  vld; // @[Reg.scala 19:20]
  reg [31:0] _RAND_350;
  reg  lastVld; // @[MuxLayer.scala 66:24]
  reg [31:0] _RAND_351;
  wire  _T_1052; // @[MuxLayer.scala 19:15]
  wire [6:0] _T_1054; // @[MuxLayer.scala 20:18]
  wire [5:0] _T_1055; // @[MuxLayer.scala 20:18]
  wire [5:0] _GEN_0; // @[MuxLayer.scala 19:23]
  wire  _T_1057; // @[MuxLayer.scala 22:34]
  wire  _T_1058; // @[MuxLayer.scala 22:26]
  wire [5:0] _GEN_1; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_2; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_3; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_4; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_5; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_6; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_7; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_8; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_9; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_10; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_11; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_12; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_13; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_14; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_15; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_16; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_17; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_18; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_19; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_20; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_21; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_22; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_23; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_24; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_25; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_26; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_27; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_28; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_29; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_30; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_31; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_32; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_33; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_34; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_35; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_36; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_37; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_38; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_39; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_40; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_41; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_42; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_43; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_44; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_45; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_46; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_47; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_48; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_49; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_50; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_51; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_52; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_53; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_54; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_55; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_56; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_57; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_58; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_59; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_60; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_61; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_62; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_63; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_64; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_65; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_66; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_67; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_68; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_69; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_70; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_71; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_72; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_73; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_74; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_75; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_76; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_77; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_78; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_79; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_80; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_81; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_82; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_83; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_84; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_85; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_86; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_87; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_88; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_89; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_90; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_91; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_92; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_93; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_94; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_95; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_96; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_97; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_98; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_99; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_100; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_101; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_102; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_103; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_104; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_105; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_106; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_107; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_108; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_109; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_110; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_111; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_112; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_113; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_114; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_115; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_116; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_117; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_118; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_119; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_120; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_121; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_122; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_123; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_124; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_125; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_126; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_127; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_128; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_129; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_130; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_131; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_132; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_133; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_134; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_135; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_136; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_137; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_138; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_139; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_140; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_141; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_142; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_143; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_144; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_145; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_146; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_147; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_148; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_149; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_150; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_151; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_152; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_153; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_154; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_155; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_156; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_157; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_158; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_159; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_160; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_161; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_162; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_163; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_164; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_165; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_166; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_167; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_168; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_169; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_170; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_171; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_172; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_173; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_174; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_175; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_176; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_177; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_178; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_179; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_180; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_181; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_182; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_183; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_184; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_185; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_186; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_187; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_188; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_189; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_190; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_191; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_192; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_193; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_194; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_195; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_196; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_197; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_198; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_199; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_200; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_201; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_202; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_203; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_204; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_205; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_206; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_207; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_208; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_209; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_210; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_211; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_212; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_213; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_214; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_215; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_216; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_217; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_218; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_219; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_220; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_221; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_222; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_223; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_224; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_225; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_226; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_227; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_228; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_229; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_230; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_231; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_232; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_233; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_234; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_235; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_236; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_237; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_238; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_239; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_240; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_241; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_242; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_243; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_244; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_245; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_246; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_247; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_248; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_249; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_250; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_251; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_252; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_253; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_254; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_255; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_256; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_257; // @[MuxLayer.scala 22:44]
  wire  _T_1061; // @[MuxLayer.scala 29:15]
  wire  _GEN_258; // @[MuxLayer.scala 29:36]
  wire  _T_1063; // @[MuxLayer.scala 32:26]
  wire  _GEN_259; // @[MuxLayer.scala 32:38]
  wire [1:0] _T_1065; // @[MuxLayer.scala 45:19]
  wire [1:0] _T_1068; // @[MuxLayer.scala 45:19]
  wire [1:0] _T_1073; // @[MuxLayer.scala 45:19]
  wire  _T_1090; // @[MuxLayer.scala 55:25]
  wire [15:0] _GEN_266; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_267; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_268; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_269; // @[MuxLayer.scala 55:35]
  wire  _T_1092; // @[MuxLayer.scala 55:25]
  wire [15:0] _GEN_270; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_271; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_272; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_273; // @[MuxLayer.scala 55:35]
  wire  _T_1094; // @[MuxLayer.scala 55:25]
  wire [15:0] _GEN_274; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_275; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_276; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_277; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_278; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_279; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_280; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_281; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_282; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_283; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_284; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_285; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_286; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_287; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_288; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_289; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_290; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_291; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_292; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_293; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_294; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_295; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_296; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_297; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_298; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_299; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_300; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_301; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_302; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_303; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_304; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_305; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_306; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_307; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_308; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_309; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_310; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_311; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_312; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_313; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_314; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_315; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_316; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_317; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_318; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_319; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_320; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_321; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_322; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_323; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_324; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_325; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_326; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_327; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_328; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_329; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_330; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_331; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_332; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_333; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_334; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_335; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_336; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_337; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_338; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_339; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_340; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_341; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_342; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_343; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_344; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_345; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_346; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_347; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_348; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_349; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_350; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_351; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_352; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_353; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_354; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_355; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_356; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_357; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_358; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_359; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_360; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_361; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_362; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_363; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_364; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_365; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_366; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_367; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_368; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_369; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_370; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_371; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_372; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_373; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_374; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_375; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_376; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_377; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_378; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_379; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_380; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_381; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_382; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_383; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_384; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_385; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_386; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_387; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_388; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_389; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_390; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_391; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_392; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_393; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_394; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_395; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_396; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_397; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_398; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_399; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_400; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_401; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_402; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_403; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_404; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_405; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_406; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_407; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_408; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_409; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_410; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_411; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_412; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_413; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_414; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_415; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_416; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_417; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_418; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_419; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_420; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_421; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_422; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_423; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_424; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_425; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_426; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_427; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_428; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_429; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_430; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_431; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_432; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_433; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_434; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_435; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_436; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_437; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_438; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_439; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_440; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_441; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_442; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_443; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_444; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_445; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_446; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_447; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_448; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_449; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_450; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_451; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_452; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_453; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_454; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_455; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_456; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_457; // @[MuxLayer.scala 55:35]
  wire  _T_1778; // @[MuxLayer.scala 55:25]
  wire [15:0] _GEN_458; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_459; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_460; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_461; // @[MuxLayer.scala 55:35]
  wire  _T_1780; // @[MuxLayer.scala 55:25]
  wire [15:0] _GEN_462; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_463; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_464; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_465; // @[MuxLayer.scala 55:35]
  wire  _T_1782; // @[MuxLayer.scala 55:25]
  wire [15:0] _GEN_466; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_467; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_468; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_469; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_470; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_471; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_472; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_473; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_474; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_475; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_476; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_477; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_478; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_479; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_480; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_481; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_482; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_483; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_484; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_485; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_486; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_487; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_488; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_489; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_490; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_491; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_492; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_493; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_494; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_495; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_496; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_497; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_498; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_499; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_500; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_501; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_502; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_503; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_504; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_505; // @[MuxLayer.scala 55:35]
  wire  _T_1950; // @[MuxLayer.scala 55:25]
  wire [15:0] _GEN_506; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_507; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_508; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_509; // @[MuxLayer.scala 55:35]
  wire  _T_1952; // @[MuxLayer.scala 55:25]
  wire [15:0] _GEN_510; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_511; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_512; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_513; // @[MuxLayer.scala 55:35]
  wire  _T_1954; // @[MuxLayer.scala 55:25]
  wire [15:0] _GEN_514; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_515; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_516; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_517; // @[MuxLayer.scala 55:35]
  wire  _T_1994; // @[MuxLayer.scala 68:27]
  assign _T_1052 = cntr > 6'h0; // @[MuxLayer.scala 19:15]
  assign _T_1054 = cntr + 6'h1; // @[MuxLayer.scala 20:18]
  assign _T_1055 = _T_1054[5:0]; // @[MuxLayer.scala 20:18]
  assign _GEN_0 = _T_1052 ? _T_1055 : cntr; // @[MuxLayer.scala 19:23]
  assign _T_1057 = cntr == 6'h0; // @[MuxLayer.scala 22:34]
  assign _T_1058 = io_dataIn_valid & _T_1057; // @[MuxLayer.scala 22:26]
  assign _GEN_1 = _T_1058 ? 6'h1 : _GEN_0; // @[MuxLayer.scala 22:44]
  assign _GEN_2 = _T_1058 ? $signed(io_dataIn_bits_0) : $signed(buffers_0_0_0); // @[MuxLayer.scala 22:44]
  assign _GEN_3 = _T_1058 ? $signed(io_dataIn_bits_1) : $signed(buffers_0_0_1); // @[MuxLayer.scala 22:44]
  assign _GEN_4 = _T_1058 ? $signed(io_dataIn_bits_2) : $signed(buffers_0_0_2); // @[MuxLayer.scala 22:44]
  assign _GEN_5 = _T_1058 ? $signed(io_dataIn_bits_3) : $signed(buffers_0_0_3); // @[MuxLayer.scala 22:44]
  assign _GEN_6 = _T_1058 ? $signed(io_dataIn_bits_4) : $signed(buffers_0_1_0); // @[MuxLayer.scala 22:44]
  assign _GEN_7 = _T_1058 ? $signed(io_dataIn_bits_5) : $signed(buffers_0_1_1); // @[MuxLayer.scala 22:44]
  assign _GEN_8 = _T_1058 ? $signed(io_dataIn_bits_6) : $signed(buffers_0_1_2); // @[MuxLayer.scala 22:44]
  assign _GEN_9 = _T_1058 ? $signed(io_dataIn_bits_7) : $signed(buffers_0_1_3); // @[MuxLayer.scala 22:44]
  assign _GEN_10 = _T_1058 ? $signed(io_dataIn_bits_8) : $signed(buffers_0_2_0); // @[MuxLayer.scala 22:44]
  assign _GEN_11 = _T_1058 ? $signed(io_dataIn_bits_9) : $signed(buffers_0_2_1); // @[MuxLayer.scala 22:44]
  assign _GEN_12 = _T_1058 ? $signed(io_dataIn_bits_10) : $signed(buffers_0_2_2); // @[MuxLayer.scala 22:44]
  assign _GEN_13 = _T_1058 ? $signed(io_dataIn_bits_11) : $signed(buffers_0_2_3); // @[MuxLayer.scala 22:44]
  assign _GEN_14 = _T_1058 ? $signed(io_dataIn_bits_12) : $signed(buffers_0_3_0); // @[MuxLayer.scala 22:44]
  assign _GEN_15 = _T_1058 ? $signed(io_dataIn_bits_13) : $signed(buffers_0_3_1); // @[MuxLayer.scala 22:44]
  assign _GEN_16 = _T_1058 ? $signed(io_dataIn_bits_14) : $signed(buffers_0_3_2); // @[MuxLayer.scala 22:44]
  assign _GEN_17 = _T_1058 ? $signed(io_dataIn_bits_15) : $signed(buffers_0_3_3); // @[MuxLayer.scala 22:44]
  assign _GEN_18 = _T_1058 ? $signed(io_dataIn_bits_16) : $signed(buffers_0_4_0); // @[MuxLayer.scala 22:44]
  assign _GEN_19 = _T_1058 ? $signed(io_dataIn_bits_17) : $signed(buffers_0_4_1); // @[MuxLayer.scala 22:44]
  assign _GEN_20 = _T_1058 ? $signed(io_dataIn_bits_18) : $signed(buffers_0_4_2); // @[MuxLayer.scala 22:44]
  assign _GEN_21 = _T_1058 ? $signed(io_dataIn_bits_19) : $signed(buffers_0_4_3); // @[MuxLayer.scala 22:44]
  assign _GEN_22 = _T_1058 ? $signed(io_dataIn_bits_20) : $signed(buffers_0_5_0); // @[MuxLayer.scala 22:44]
  assign _GEN_23 = _T_1058 ? $signed(io_dataIn_bits_21) : $signed(buffers_0_5_1); // @[MuxLayer.scala 22:44]
  assign _GEN_24 = _T_1058 ? $signed(io_dataIn_bits_22) : $signed(buffers_0_5_2); // @[MuxLayer.scala 22:44]
  assign _GEN_25 = _T_1058 ? $signed(io_dataIn_bits_23) : $signed(buffers_0_5_3); // @[MuxLayer.scala 22:44]
  assign _GEN_26 = _T_1058 ? $signed(io_dataIn_bits_24) : $signed(buffers_0_6_0); // @[MuxLayer.scala 22:44]
  assign _GEN_27 = _T_1058 ? $signed(io_dataIn_bits_25) : $signed(buffers_0_6_1); // @[MuxLayer.scala 22:44]
  assign _GEN_28 = _T_1058 ? $signed(io_dataIn_bits_26) : $signed(buffers_0_6_2); // @[MuxLayer.scala 22:44]
  assign _GEN_29 = _T_1058 ? $signed(io_dataIn_bits_27) : $signed(buffers_0_6_3); // @[MuxLayer.scala 22:44]
  assign _GEN_30 = _T_1058 ? $signed(io_dataIn_bits_28) : $signed(buffers_0_7_0); // @[MuxLayer.scala 22:44]
  assign _GEN_31 = _T_1058 ? $signed(io_dataIn_bits_29) : $signed(buffers_0_7_1); // @[MuxLayer.scala 22:44]
  assign _GEN_32 = _T_1058 ? $signed(io_dataIn_bits_30) : $signed(buffers_0_7_2); // @[MuxLayer.scala 22:44]
  assign _GEN_33 = _T_1058 ? $signed(io_dataIn_bits_31) : $signed(buffers_0_7_3); // @[MuxLayer.scala 22:44]
  assign _GEN_34 = _T_1058 ? $signed(io_dataIn_bits_32) : $signed(buffers_0_8_0); // @[MuxLayer.scala 22:44]
  assign _GEN_35 = _T_1058 ? $signed(io_dataIn_bits_33) : $signed(buffers_0_8_1); // @[MuxLayer.scala 22:44]
  assign _GEN_36 = _T_1058 ? $signed(io_dataIn_bits_34) : $signed(buffers_0_8_2); // @[MuxLayer.scala 22:44]
  assign _GEN_37 = _T_1058 ? $signed(io_dataIn_bits_35) : $signed(buffers_0_8_3); // @[MuxLayer.scala 22:44]
  assign _GEN_38 = _T_1058 ? $signed(io_dataIn_bits_36) : $signed(buffers_0_9_0); // @[MuxLayer.scala 22:44]
  assign _GEN_39 = _T_1058 ? $signed(io_dataIn_bits_37) : $signed(buffers_0_9_1); // @[MuxLayer.scala 22:44]
  assign _GEN_40 = _T_1058 ? $signed(io_dataIn_bits_38) : $signed(buffers_0_9_2); // @[MuxLayer.scala 22:44]
  assign _GEN_41 = _T_1058 ? $signed(io_dataIn_bits_39) : $signed(buffers_0_9_3); // @[MuxLayer.scala 22:44]
  assign _GEN_42 = _T_1058 ? $signed(io_dataIn_bits_40) : $signed(buffers_0_10_0); // @[MuxLayer.scala 22:44]
  assign _GEN_43 = _T_1058 ? $signed(io_dataIn_bits_41) : $signed(buffers_0_10_1); // @[MuxLayer.scala 22:44]
  assign _GEN_44 = _T_1058 ? $signed(io_dataIn_bits_42) : $signed(buffers_0_10_2); // @[MuxLayer.scala 22:44]
  assign _GEN_45 = _T_1058 ? $signed(io_dataIn_bits_43) : $signed(buffers_0_10_3); // @[MuxLayer.scala 22:44]
  assign _GEN_46 = _T_1058 ? $signed(io_dataIn_bits_44) : $signed(buffers_0_11_0); // @[MuxLayer.scala 22:44]
  assign _GEN_47 = _T_1058 ? $signed(io_dataIn_bits_45) : $signed(buffers_0_11_1); // @[MuxLayer.scala 22:44]
  assign _GEN_48 = _T_1058 ? $signed(io_dataIn_bits_46) : $signed(buffers_0_11_2); // @[MuxLayer.scala 22:44]
  assign _GEN_49 = _T_1058 ? $signed(io_dataIn_bits_47) : $signed(buffers_0_11_3); // @[MuxLayer.scala 22:44]
  assign _GEN_50 = _T_1058 ? $signed(io_dataIn_bits_48) : $signed(buffers_0_12_0); // @[MuxLayer.scala 22:44]
  assign _GEN_51 = _T_1058 ? $signed(io_dataIn_bits_49) : $signed(buffers_0_12_1); // @[MuxLayer.scala 22:44]
  assign _GEN_52 = _T_1058 ? $signed(io_dataIn_bits_50) : $signed(buffers_0_12_2); // @[MuxLayer.scala 22:44]
  assign _GEN_53 = _T_1058 ? $signed(io_dataIn_bits_51) : $signed(buffers_0_12_3); // @[MuxLayer.scala 22:44]
  assign _GEN_54 = _T_1058 ? $signed(io_dataIn_bits_52) : $signed(buffers_0_13_0); // @[MuxLayer.scala 22:44]
  assign _GEN_55 = _T_1058 ? $signed(io_dataIn_bits_53) : $signed(buffers_0_13_1); // @[MuxLayer.scala 22:44]
  assign _GEN_56 = _T_1058 ? $signed(io_dataIn_bits_54) : $signed(buffers_0_13_2); // @[MuxLayer.scala 22:44]
  assign _GEN_57 = _T_1058 ? $signed(io_dataIn_bits_55) : $signed(buffers_0_13_3); // @[MuxLayer.scala 22:44]
  assign _GEN_58 = _T_1058 ? $signed(io_dataIn_bits_56) : $signed(buffers_0_14_0); // @[MuxLayer.scala 22:44]
  assign _GEN_59 = _T_1058 ? $signed(io_dataIn_bits_57) : $signed(buffers_0_14_1); // @[MuxLayer.scala 22:44]
  assign _GEN_60 = _T_1058 ? $signed(io_dataIn_bits_58) : $signed(buffers_0_14_2); // @[MuxLayer.scala 22:44]
  assign _GEN_61 = _T_1058 ? $signed(io_dataIn_bits_59) : $signed(buffers_0_14_3); // @[MuxLayer.scala 22:44]
  assign _GEN_62 = _T_1058 ? $signed(io_dataIn_bits_60) : $signed(buffers_0_15_0); // @[MuxLayer.scala 22:44]
  assign _GEN_63 = _T_1058 ? $signed(io_dataIn_bits_61) : $signed(buffers_0_15_1); // @[MuxLayer.scala 22:44]
  assign _GEN_64 = _T_1058 ? $signed(io_dataIn_bits_62) : $signed(buffers_0_15_2); // @[MuxLayer.scala 22:44]
  assign _GEN_65 = _T_1058 ? $signed(io_dataIn_bits_63) : $signed(buffers_0_15_3); // @[MuxLayer.scala 22:44]
  assign _GEN_66 = _T_1058 ? $signed(io_dataIn_bits_64) : $signed(buffers_0_16_0); // @[MuxLayer.scala 22:44]
  assign _GEN_67 = _T_1058 ? $signed(io_dataIn_bits_65) : $signed(buffers_0_16_1); // @[MuxLayer.scala 22:44]
  assign _GEN_68 = _T_1058 ? $signed(io_dataIn_bits_66) : $signed(buffers_0_16_2); // @[MuxLayer.scala 22:44]
  assign _GEN_69 = _T_1058 ? $signed(io_dataIn_bits_67) : $signed(buffers_0_16_3); // @[MuxLayer.scala 22:44]
  assign _GEN_70 = _T_1058 ? $signed(io_dataIn_bits_68) : $signed(buffers_0_17_0); // @[MuxLayer.scala 22:44]
  assign _GEN_71 = _T_1058 ? $signed(io_dataIn_bits_69) : $signed(buffers_0_17_1); // @[MuxLayer.scala 22:44]
  assign _GEN_72 = _T_1058 ? $signed(io_dataIn_bits_70) : $signed(buffers_0_17_2); // @[MuxLayer.scala 22:44]
  assign _GEN_73 = _T_1058 ? $signed(io_dataIn_bits_71) : $signed(buffers_0_17_3); // @[MuxLayer.scala 22:44]
  assign _GEN_74 = _T_1058 ? $signed(io_dataIn_bits_72) : $signed(buffers_0_18_0); // @[MuxLayer.scala 22:44]
  assign _GEN_75 = _T_1058 ? $signed(io_dataIn_bits_73) : $signed(buffers_0_18_1); // @[MuxLayer.scala 22:44]
  assign _GEN_76 = _T_1058 ? $signed(io_dataIn_bits_74) : $signed(buffers_0_18_2); // @[MuxLayer.scala 22:44]
  assign _GEN_77 = _T_1058 ? $signed(io_dataIn_bits_75) : $signed(buffers_0_18_3); // @[MuxLayer.scala 22:44]
  assign _GEN_78 = _T_1058 ? $signed(io_dataIn_bits_76) : $signed(buffers_0_19_0); // @[MuxLayer.scala 22:44]
  assign _GEN_79 = _T_1058 ? $signed(io_dataIn_bits_77) : $signed(buffers_0_19_1); // @[MuxLayer.scala 22:44]
  assign _GEN_80 = _T_1058 ? $signed(io_dataIn_bits_78) : $signed(buffers_0_19_2); // @[MuxLayer.scala 22:44]
  assign _GEN_81 = _T_1058 ? $signed(io_dataIn_bits_79) : $signed(buffers_0_19_3); // @[MuxLayer.scala 22:44]
  assign _GEN_82 = _T_1058 ? $signed(io_dataIn_bits_80) : $signed(buffers_0_20_0); // @[MuxLayer.scala 22:44]
  assign _GEN_83 = _T_1058 ? $signed(io_dataIn_bits_81) : $signed(buffers_0_20_1); // @[MuxLayer.scala 22:44]
  assign _GEN_84 = _T_1058 ? $signed(io_dataIn_bits_82) : $signed(buffers_0_20_2); // @[MuxLayer.scala 22:44]
  assign _GEN_85 = _T_1058 ? $signed(io_dataIn_bits_83) : $signed(buffers_0_20_3); // @[MuxLayer.scala 22:44]
  assign _GEN_86 = _T_1058 ? $signed(io_dataIn_bits_84) : $signed(buffers_0_21_0); // @[MuxLayer.scala 22:44]
  assign _GEN_87 = _T_1058 ? $signed(io_dataIn_bits_85) : $signed(buffers_0_21_1); // @[MuxLayer.scala 22:44]
  assign _GEN_88 = _T_1058 ? $signed(io_dataIn_bits_86) : $signed(buffers_0_21_2); // @[MuxLayer.scala 22:44]
  assign _GEN_89 = _T_1058 ? $signed(io_dataIn_bits_87) : $signed(buffers_0_21_3); // @[MuxLayer.scala 22:44]
  assign _GEN_90 = _T_1058 ? $signed(io_dataIn_bits_88) : $signed(buffers_0_22_0); // @[MuxLayer.scala 22:44]
  assign _GEN_91 = _T_1058 ? $signed(io_dataIn_bits_89) : $signed(buffers_0_22_1); // @[MuxLayer.scala 22:44]
  assign _GEN_92 = _T_1058 ? $signed(io_dataIn_bits_90) : $signed(buffers_0_22_2); // @[MuxLayer.scala 22:44]
  assign _GEN_93 = _T_1058 ? $signed(io_dataIn_bits_91) : $signed(buffers_0_22_3); // @[MuxLayer.scala 22:44]
  assign _GEN_94 = _T_1058 ? $signed(io_dataIn_bits_92) : $signed(buffers_0_23_0); // @[MuxLayer.scala 22:44]
  assign _GEN_95 = _T_1058 ? $signed(io_dataIn_bits_93) : $signed(buffers_0_23_1); // @[MuxLayer.scala 22:44]
  assign _GEN_96 = _T_1058 ? $signed(io_dataIn_bits_94) : $signed(buffers_0_23_2); // @[MuxLayer.scala 22:44]
  assign _GEN_97 = _T_1058 ? $signed(io_dataIn_bits_95) : $signed(buffers_0_23_3); // @[MuxLayer.scala 22:44]
  assign _GEN_98 = _T_1058 ? $signed(io_dataIn_bits_96) : $signed(buffers_0_24_0); // @[MuxLayer.scala 22:44]
  assign _GEN_99 = _T_1058 ? $signed(io_dataIn_bits_97) : $signed(buffers_0_24_1); // @[MuxLayer.scala 22:44]
  assign _GEN_100 = _T_1058 ? $signed(io_dataIn_bits_98) : $signed(buffers_0_24_2); // @[MuxLayer.scala 22:44]
  assign _GEN_101 = _T_1058 ? $signed(io_dataIn_bits_99) : $signed(buffers_0_24_3); // @[MuxLayer.scala 22:44]
  assign _GEN_102 = _T_1058 ? $signed(io_dataIn_bits_100) : $signed(buffers_0_25_0); // @[MuxLayer.scala 22:44]
  assign _GEN_103 = _T_1058 ? $signed(io_dataIn_bits_101) : $signed(buffers_0_25_1); // @[MuxLayer.scala 22:44]
  assign _GEN_104 = _T_1058 ? $signed(io_dataIn_bits_102) : $signed(buffers_0_25_2); // @[MuxLayer.scala 22:44]
  assign _GEN_105 = _T_1058 ? $signed(io_dataIn_bits_103) : $signed(buffers_0_25_3); // @[MuxLayer.scala 22:44]
  assign _GEN_106 = _T_1058 ? $signed(io_dataIn_bits_104) : $signed(buffers_0_26_0); // @[MuxLayer.scala 22:44]
  assign _GEN_107 = _T_1058 ? $signed(io_dataIn_bits_105) : $signed(buffers_0_26_1); // @[MuxLayer.scala 22:44]
  assign _GEN_108 = _T_1058 ? $signed(io_dataIn_bits_106) : $signed(buffers_0_26_2); // @[MuxLayer.scala 22:44]
  assign _GEN_109 = _T_1058 ? $signed(io_dataIn_bits_107) : $signed(buffers_0_26_3); // @[MuxLayer.scala 22:44]
  assign _GEN_110 = _T_1058 ? $signed(io_dataIn_bits_108) : $signed(buffers_0_27_0); // @[MuxLayer.scala 22:44]
  assign _GEN_111 = _T_1058 ? $signed(io_dataIn_bits_109) : $signed(buffers_0_27_1); // @[MuxLayer.scala 22:44]
  assign _GEN_112 = _T_1058 ? $signed(io_dataIn_bits_110) : $signed(buffers_0_27_2); // @[MuxLayer.scala 22:44]
  assign _GEN_113 = _T_1058 ? $signed(io_dataIn_bits_111) : $signed(buffers_0_27_3); // @[MuxLayer.scala 22:44]
  assign _GEN_114 = _T_1058 ? $signed(io_dataIn_bits_112) : $signed(buffers_0_28_0); // @[MuxLayer.scala 22:44]
  assign _GEN_115 = _T_1058 ? $signed(io_dataIn_bits_113) : $signed(buffers_0_28_1); // @[MuxLayer.scala 22:44]
  assign _GEN_116 = _T_1058 ? $signed(io_dataIn_bits_114) : $signed(buffers_0_28_2); // @[MuxLayer.scala 22:44]
  assign _GEN_117 = _T_1058 ? $signed(io_dataIn_bits_115) : $signed(buffers_0_28_3); // @[MuxLayer.scala 22:44]
  assign _GEN_118 = _T_1058 ? $signed(io_dataIn_bits_116) : $signed(buffers_0_29_0); // @[MuxLayer.scala 22:44]
  assign _GEN_119 = _T_1058 ? $signed(io_dataIn_bits_117) : $signed(buffers_0_29_1); // @[MuxLayer.scala 22:44]
  assign _GEN_120 = _T_1058 ? $signed(io_dataIn_bits_118) : $signed(buffers_0_29_2); // @[MuxLayer.scala 22:44]
  assign _GEN_121 = _T_1058 ? $signed(io_dataIn_bits_119) : $signed(buffers_0_29_3); // @[MuxLayer.scala 22:44]
  assign _GEN_122 = _T_1058 ? $signed(io_dataIn_bits_120) : $signed(buffers_0_30_0); // @[MuxLayer.scala 22:44]
  assign _GEN_123 = _T_1058 ? $signed(io_dataIn_bits_121) : $signed(buffers_0_30_1); // @[MuxLayer.scala 22:44]
  assign _GEN_124 = _T_1058 ? $signed(io_dataIn_bits_122) : $signed(buffers_0_30_2); // @[MuxLayer.scala 22:44]
  assign _GEN_125 = _T_1058 ? $signed(io_dataIn_bits_123) : $signed(buffers_0_30_3); // @[MuxLayer.scala 22:44]
  assign _GEN_126 = _T_1058 ? $signed(io_dataIn_bits_124) : $signed(buffers_0_31_0); // @[MuxLayer.scala 22:44]
  assign _GEN_127 = _T_1058 ? $signed(io_dataIn_bits_125) : $signed(buffers_0_31_1); // @[MuxLayer.scala 22:44]
  assign _GEN_128 = _T_1058 ? $signed(io_dataIn_bits_126) : $signed(buffers_0_31_2); // @[MuxLayer.scala 22:44]
  assign _GEN_129 = _T_1058 ? $signed(io_dataIn_bits_127) : $signed(buffers_0_31_3); // @[MuxLayer.scala 22:44]
  assign _GEN_130 = _T_1058 ? $signed(io_dataIn_bits_128) : $signed(buffers_0_32_0); // @[MuxLayer.scala 22:44]
  assign _GEN_131 = _T_1058 ? $signed(io_dataIn_bits_129) : $signed(buffers_0_32_1); // @[MuxLayer.scala 22:44]
  assign _GEN_132 = _T_1058 ? $signed(io_dataIn_bits_130) : $signed(buffers_0_32_2); // @[MuxLayer.scala 22:44]
  assign _GEN_133 = _T_1058 ? $signed(io_dataIn_bits_131) : $signed(buffers_0_32_3); // @[MuxLayer.scala 22:44]
  assign _GEN_134 = _T_1058 ? $signed(io_dataIn_bits_132) : $signed(buffers_0_33_0); // @[MuxLayer.scala 22:44]
  assign _GEN_135 = _T_1058 ? $signed(io_dataIn_bits_133) : $signed(buffers_0_33_1); // @[MuxLayer.scala 22:44]
  assign _GEN_136 = _T_1058 ? $signed(io_dataIn_bits_134) : $signed(buffers_0_33_2); // @[MuxLayer.scala 22:44]
  assign _GEN_137 = _T_1058 ? $signed(io_dataIn_bits_135) : $signed(buffers_0_33_3); // @[MuxLayer.scala 22:44]
  assign _GEN_138 = _T_1058 ? $signed(io_dataIn_bits_136) : $signed(buffers_0_34_0); // @[MuxLayer.scala 22:44]
  assign _GEN_139 = _T_1058 ? $signed(io_dataIn_bits_137) : $signed(buffers_0_34_1); // @[MuxLayer.scala 22:44]
  assign _GEN_140 = _T_1058 ? $signed(io_dataIn_bits_138) : $signed(buffers_0_34_2); // @[MuxLayer.scala 22:44]
  assign _GEN_141 = _T_1058 ? $signed(io_dataIn_bits_139) : $signed(buffers_0_34_3); // @[MuxLayer.scala 22:44]
  assign _GEN_142 = _T_1058 ? $signed(io_dataIn_bits_140) : $signed(buffers_0_35_0); // @[MuxLayer.scala 22:44]
  assign _GEN_143 = _T_1058 ? $signed(io_dataIn_bits_141) : $signed(buffers_0_35_1); // @[MuxLayer.scala 22:44]
  assign _GEN_144 = _T_1058 ? $signed(io_dataIn_bits_142) : $signed(buffers_0_35_2); // @[MuxLayer.scala 22:44]
  assign _GEN_145 = _T_1058 ? $signed(io_dataIn_bits_143) : $signed(buffers_0_35_3); // @[MuxLayer.scala 22:44]
  assign _GEN_146 = _T_1058 ? $signed(io_dataIn_bits_144) : $signed(buffers_0_36_0); // @[MuxLayer.scala 22:44]
  assign _GEN_147 = _T_1058 ? $signed(io_dataIn_bits_145) : $signed(buffers_0_36_1); // @[MuxLayer.scala 22:44]
  assign _GEN_148 = _T_1058 ? $signed(io_dataIn_bits_146) : $signed(buffers_0_36_2); // @[MuxLayer.scala 22:44]
  assign _GEN_149 = _T_1058 ? $signed(io_dataIn_bits_147) : $signed(buffers_0_36_3); // @[MuxLayer.scala 22:44]
  assign _GEN_150 = _T_1058 ? $signed(io_dataIn_bits_148) : $signed(buffers_0_37_0); // @[MuxLayer.scala 22:44]
  assign _GEN_151 = _T_1058 ? $signed(io_dataIn_bits_149) : $signed(buffers_0_37_1); // @[MuxLayer.scala 22:44]
  assign _GEN_152 = _T_1058 ? $signed(io_dataIn_bits_150) : $signed(buffers_0_37_2); // @[MuxLayer.scala 22:44]
  assign _GEN_153 = _T_1058 ? $signed(io_dataIn_bits_151) : $signed(buffers_0_37_3); // @[MuxLayer.scala 22:44]
  assign _GEN_154 = _T_1058 ? $signed(io_dataIn_bits_152) : $signed(buffers_0_38_0); // @[MuxLayer.scala 22:44]
  assign _GEN_155 = _T_1058 ? $signed(io_dataIn_bits_153) : $signed(buffers_0_38_1); // @[MuxLayer.scala 22:44]
  assign _GEN_156 = _T_1058 ? $signed(io_dataIn_bits_154) : $signed(buffers_0_38_2); // @[MuxLayer.scala 22:44]
  assign _GEN_157 = _T_1058 ? $signed(io_dataIn_bits_155) : $signed(buffers_0_38_3); // @[MuxLayer.scala 22:44]
  assign _GEN_158 = _T_1058 ? $signed(io_dataIn_bits_156) : $signed(buffers_0_39_0); // @[MuxLayer.scala 22:44]
  assign _GEN_159 = _T_1058 ? $signed(io_dataIn_bits_157) : $signed(buffers_0_39_1); // @[MuxLayer.scala 22:44]
  assign _GEN_160 = _T_1058 ? $signed(io_dataIn_bits_158) : $signed(buffers_0_39_2); // @[MuxLayer.scala 22:44]
  assign _GEN_161 = _T_1058 ? $signed(io_dataIn_bits_159) : $signed(buffers_0_39_3); // @[MuxLayer.scala 22:44]
  assign _GEN_162 = _T_1058 ? $signed(io_dataIn_bits_160) : $signed(buffers_0_40_0); // @[MuxLayer.scala 22:44]
  assign _GEN_163 = _T_1058 ? $signed(io_dataIn_bits_161) : $signed(buffers_0_40_1); // @[MuxLayer.scala 22:44]
  assign _GEN_164 = _T_1058 ? $signed(io_dataIn_bits_162) : $signed(buffers_0_40_2); // @[MuxLayer.scala 22:44]
  assign _GEN_165 = _T_1058 ? $signed(io_dataIn_bits_163) : $signed(buffers_0_40_3); // @[MuxLayer.scala 22:44]
  assign _GEN_166 = _T_1058 ? $signed(io_dataIn_bits_164) : $signed(buffers_0_41_0); // @[MuxLayer.scala 22:44]
  assign _GEN_167 = _T_1058 ? $signed(io_dataIn_bits_165) : $signed(buffers_0_41_1); // @[MuxLayer.scala 22:44]
  assign _GEN_168 = _T_1058 ? $signed(io_dataIn_bits_166) : $signed(buffers_0_41_2); // @[MuxLayer.scala 22:44]
  assign _GEN_169 = _T_1058 ? $signed(io_dataIn_bits_167) : $signed(buffers_0_41_3); // @[MuxLayer.scala 22:44]
  assign _GEN_170 = _T_1058 ? $signed(io_dataIn_bits_168) : $signed(buffers_0_42_0); // @[MuxLayer.scala 22:44]
  assign _GEN_171 = _T_1058 ? $signed(io_dataIn_bits_169) : $signed(buffers_0_42_1); // @[MuxLayer.scala 22:44]
  assign _GEN_172 = _T_1058 ? $signed(io_dataIn_bits_170) : $signed(buffers_0_42_2); // @[MuxLayer.scala 22:44]
  assign _GEN_173 = _T_1058 ? $signed(io_dataIn_bits_171) : $signed(buffers_0_42_3); // @[MuxLayer.scala 22:44]
  assign _GEN_174 = _T_1058 ? $signed(io_dataIn_bits_172) : $signed(buffers_0_43_0); // @[MuxLayer.scala 22:44]
  assign _GEN_175 = _T_1058 ? $signed(io_dataIn_bits_173) : $signed(buffers_0_43_1); // @[MuxLayer.scala 22:44]
  assign _GEN_176 = _T_1058 ? $signed(io_dataIn_bits_174) : $signed(buffers_0_43_2); // @[MuxLayer.scala 22:44]
  assign _GEN_177 = _T_1058 ? $signed(io_dataIn_bits_175) : $signed(buffers_0_43_3); // @[MuxLayer.scala 22:44]
  assign _GEN_178 = _T_1058 ? $signed(io_dataIn_bits_176) : $signed(buffers_0_44_0); // @[MuxLayer.scala 22:44]
  assign _GEN_179 = _T_1058 ? $signed(io_dataIn_bits_177) : $signed(buffers_0_44_1); // @[MuxLayer.scala 22:44]
  assign _GEN_180 = _T_1058 ? $signed(io_dataIn_bits_178) : $signed(buffers_0_44_2); // @[MuxLayer.scala 22:44]
  assign _GEN_181 = _T_1058 ? $signed(io_dataIn_bits_179) : $signed(buffers_0_44_3); // @[MuxLayer.scala 22:44]
  assign _GEN_182 = _T_1058 ? $signed(io_dataIn_bits_180) : $signed(buffers_0_45_0); // @[MuxLayer.scala 22:44]
  assign _GEN_183 = _T_1058 ? $signed(io_dataIn_bits_181) : $signed(buffers_0_45_1); // @[MuxLayer.scala 22:44]
  assign _GEN_184 = _T_1058 ? $signed(io_dataIn_bits_182) : $signed(buffers_0_45_2); // @[MuxLayer.scala 22:44]
  assign _GEN_185 = _T_1058 ? $signed(io_dataIn_bits_183) : $signed(buffers_0_45_3); // @[MuxLayer.scala 22:44]
  assign _GEN_186 = _T_1058 ? $signed(io_dataIn_bits_184) : $signed(buffers_0_46_0); // @[MuxLayer.scala 22:44]
  assign _GEN_187 = _T_1058 ? $signed(io_dataIn_bits_185) : $signed(buffers_0_46_1); // @[MuxLayer.scala 22:44]
  assign _GEN_188 = _T_1058 ? $signed(io_dataIn_bits_186) : $signed(buffers_0_46_2); // @[MuxLayer.scala 22:44]
  assign _GEN_189 = _T_1058 ? $signed(io_dataIn_bits_187) : $signed(buffers_0_46_3); // @[MuxLayer.scala 22:44]
  assign _GEN_190 = _T_1058 ? $signed(io_dataIn_bits_188) : $signed(buffers_0_47_0); // @[MuxLayer.scala 22:44]
  assign _GEN_191 = _T_1058 ? $signed(io_dataIn_bits_189) : $signed(buffers_0_47_1); // @[MuxLayer.scala 22:44]
  assign _GEN_192 = _T_1058 ? $signed(io_dataIn_bits_190) : $signed(buffers_0_47_2); // @[MuxLayer.scala 22:44]
  assign _GEN_193 = _T_1058 ? $signed(io_dataIn_bits_191) : $signed(buffers_0_47_3); // @[MuxLayer.scala 22:44]
  assign _GEN_194 = _T_1058 ? $signed(io_dataIn_bits_192) : $signed(buffers_0_48_0); // @[MuxLayer.scala 22:44]
  assign _GEN_195 = _T_1058 ? $signed(io_dataIn_bits_193) : $signed(buffers_0_48_1); // @[MuxLayer.scala 22:44]
  assign _GEN_196 = _T_1058 ? $signed(io_dataIn_bits_194) : $signed(buffers_0_48_2); // @[MuxLayer.scala 22:44]
  assign _GEN_197 = _T_1058 ? $signed(io_dataIn_bits_195) : $signed(buffers_0_48_3); // @[MuxLayer.scala 22:44]
  assign _GEN_198 = _T_1058 ? $signed(io_dataIn_bits_196) : $signed(buffers_0_49_0); // @[MuxLayer.scala 22:44]
  assign _GEN_199 = _T_1058 ? $signed(io_dataIn_bits_197) : $signed(buffers_0_49_1); // @[MuxLayer.scala 22:44]
  assign _GEN_200 = _T_1058 ? $signed(io_dataIn_bits_198) : $signed(buffers_0_49_2); // @[MuxLayer.scala 22:44]
  assign _GEN_201 = _T_1058 ? $signed(io_dataIn_bits_199) : $signed(buffers_0_49_3); // @[MuxLayer.scala 22:44]
  assign _GEN_202 = _T_1058 ? $signed(io_dataIn_bits_200) : $signed(buffers_0_50_0); // @[MuxLayer.scala 22:44]
  assign _GEN_203 = _T_1058 ? $signed(io_dataIn_bits_201) : $signed(buffers_0_50_1); // @[MuxLayer.scala 22:44]
  assign _GEN_204 = _T_1058 ? $signed(io_dataIn_bits_202) : $signed(buffers_0_50_2); // @[MuxLayer.scala 22:44]
  assign _GEN_205 = _T_1058 ? $signed(io_dataIn_bits_203) : $signed(buffers_0_50_3); // @[MuxLayer.scala 22:44]
  assign _GEN_206 = _T_1058 ? $signed(io_dataIn_bits_204) : $signed(buffers_0_51_0); // @[MuxLayer.scala 22:44]
  assign _GEN_207 = _T_1058 ? $signed(io_dataIn_bits_205) : $signed(buffers_0_51_1); // @[MuxLayer.scala 22:44]
  assign _GEN_208 = _T_1058 ? $signed(io_dataIn_bits_206) : $signed(buffers_0_51_2); // @[MuxLayer.scala 22:44]
  assign _GEN_209 = _T_1058 ? $signed(io_dataIn_bits_207) : $signed(buffers_0_51_3); // @[MuxLayer.scala 22:44]
  assign _GEN_210 = _T_1058 ? $signed(io_dataIn_bits_208) : $signed(buffers_0_52_0); // @[MuxLayer.scala 22:44]
  assign _GEN_211 = _T_1058 ? $signed(io_dataIn_bits_209) : $signed(buffers_0_52_1); // @[MuxLayer.scala 22:44]
  assign _GEN_212 = _T_1058 ? $signed(io_dataIn_bits_210) : $signed(buffers_0_52_2); // @[MuxLayer.scala 22:44]
  assign _GEN_213 = _T_1058 ? $signed(io_dataIn_bits_211) : $signed(buffers_0_52_3); // @[MuxLayer.scala 22:44]
  assign _GEN_214 = _T_1058 ? $signed(io_dataIn_bits_212) : $signed(buffers_0_53_0); // @[MuxLayer.scala 22:44]
  assign _GEN_215 = _T_1058 ? $signed(io_dataIn_bits_213) : $signed(buffers_0_53_1); // @[MuxLayer.scala 22:44]
  assign _GEN_216 = _T_1058 ? $signed(io_dataIn_bits_214) : $signed(buffers_0_53_2); // @[MuxLayer.scala 22:44]
  assign _GEN_217 = _T_1058 ? $signed(io_dataIn_bits_215) : $signed(buffers_0_53_3); // @[MuxLayer.scala 22:44]
  assign _GEN_218 = _T_1058 ? $signed(io_dataIn_bits_216) : $signed(buffers_0_54_0); // @[MuxLayer.scala 22:44]
  assign _GEN_219 = _T_1058 ? $signed(io_dataIn_bits_217) : $signed(buffers_0_54_1); // @[MuxLayer.scala 22:44]
  assign _GEN_220 = _T_1058 ? $signed(io_dataIn_bits_218) : $signed(buffers_0_54_2); // @[MuxLayer.scala 22:44]
  assign _GEN_221 = _T_1058 ? $signed(io_dataIn_bits_219) : $signed(buffers_0_54_3); // @[MuxLayer.scala 22:44]
  assign _GEN_222 = _T_1058 ? $signed(io_dataIn_bits_220) : $signed(buffers_0_55_0); // @[MuxLayer.scala 22:44]
  assign _GEN_223 = _T_1058 ? $signed(io_dataIn_bits_221) : $signed(buffers_0_55_1); // @[MuxLayer.scala 22:44]
  assign _GEN_224 = _T_1058 ? $signed(io_dataIn_bits_222) : $signed(buffers_0_55_2); // @[MuxLayer.scala 22:44]
  assign _GEN_225 = _T_1058 ? $signed(io_dataIn_bits_223) : $signed(buffers_0_55_3); // @[MuxLayer.scala 22:44]
  assign _GEN_226 = _T_1058 ? $signed(io_dataIn_bits_224) : $signed(buffers_0_56_0); // @[MuxLayer.scala 22:44]
  assign _GEN_227 = _T_1058 ? $signed(io_dataIn_bits_225) : $signed(buffers_0_56_1); // @[MuxLayer.scala 22:44]
  assign _GEN_228 = _T_1058 ? $signed(io_dataIn_bits_226) : $signed(buffers_0_56_2); // @[MuxLayer.scala 22:44]
  assign _GEN_229 = _T_1058 ? $signed(io_dataIn_bits_227) : $signed(buffers_0_56_3); // @[MuxLayer.scala 22:44]
  assign _GEN_230 = _T_1058 ? $signed(io_dataIn_bits_228) : $signed(buffers_0_57_0); // @[MuxLayer.scala 22:44]
  assign _GEN_231 = _T_1058 ? $signed(io_dataIn_bits_229) : $signed(buffers_0_57_1); // @[MuxLayer.scala 22:44]
  assign _GEN_232 = _T_1058 ? $signed(io_dataIn_bits_230) : $signed(buffers_0_57_2); // @[MuxLayer.scala 22:44]
  assign _GEN_233 = _T_1058 ? $signed(io_dataIn_bits_231) : $signed(buffers_0_57_3); // @[MuxLayer.scala 22:44]
  assign _GEN_234 = _T_1058 ? $signed(io_dataIn_bits_232) : $signed(buffers_0_58_0); // @[MuxLayer.scala 22:44]
  assign _GEN_235 = _T_1058 ? $signed(io_dataIn_bits_233) : $signed(buffers_0_58_1); // @[MuxLayer.scala 22:44]
  assign _GEN_236 = _T_1058 ? $signed(io_dataIn_bits_234) : $signed(buffers_0_58_2); // @[MuxLayer.scala 22:44]
  assign _GEN_237 = _T_1058 ? $signed(io_dataIn_bits_235) : $signed(buffers_0_58_3); // @[MuxLayer.scala 22:44]
  assign _GEN_238 = _T_1058 ? $signed(io_dataIn_bits_236) : $signed(buffers_0_59_0); // @[MuxLayer.scala 22:44]
  assign _GEN_239 = _T_1058 ? $signed(io_dataIn_bits_237) : $signed(buffers_0_59_1); // @[MuxLayer.scala 22:44]
  assign _GEN_240 = _T_1058 ? $signed(io_dataIn_bits_238) : $signed(buffers_0_59_2); // @[MuxLayer.scala 22:44]
  assign _GEN_241 = _T_1058 ? $signed(io_dataIn_bits_239) : $signed(buffers_0_59_3); // @[MuxLayer.scala 22:44]
  assign _GEN_242 = _T_1058 ? $signed(io_dataIn_bits_240) : $signed(buffers_0_60_0); // @[MuxLayer.scala 22:44]
  assign _GEN_243 = _T_1058 ? $signed(io_dataIn_bits_241) : $signed(buffers_0_60_1); // @[MuxLayer.scala 22:44]
  assign _GEN_244 = _T_1058 ? $signed(io_dataIn_bits_242) : $signed(buffers_0_60_2); // @[MuxLayer.scala 22:44]
  assign _GEN_245 = _T_1058 ? $signed(io_dataIn_bits_243) : $signed(buffers_0_60_3); // @[MuxLayer.scala 22:44]
  assign _GEN_246 = _T_1058 ? $signed(io_dataIn_bits_244) : $signed(buffers_0_61_0); // @[MuxLayer.scala 22:44]
  assign _GEN_247 = _T_1058 ? $signed(io_dataIn_bits_245) : $signed(buffers_0_61_1); // @[MuxLayer.scala 22:44]
  assign _GEN_248 = _T_1058 ? $signed(io_dataIn_bits_246) : $signed(buffers_0_61_2); // @[MuxLayer.scala 22:44]
  assign _GEN_249 = _T_1058 ? $signed(io_dataIn_bits_247) : $signed(buffers_0_61_3); // @[MuxLayer.scala 22:44]
  assign _GEN_250 = _T_1058 ? $signed(io_dataIn_bits_248) : $signed(buffers_0_62_0); // @[MuxLayer.scala 22:44]
  assign _GEN_251 = _T_1058 ? $signed(io_dataIn_bits_249) : $signed(buffers_0_62_1); // @[MuxLayer.scala 22:44]
  assign _GEN_252 = _T_1058 ? $signed(io_dataIn_bits_250) : $signed(buffers_0_62_2); // @[MuxLayer.scala 22:44]
  assign _GEN_253 = _T_1058 ? $signed(io_dataIn_bits_251) : $signed(buffers_0_62_3); // @[MuxLayer.scala 22:44]
  assign _GEN_254 = _T_1058 ? $signed(io_dataIn_bits_252) : $signed(buffers_0_63_0); // @[MuxLayer.scala 22:44]
  assign _GEN_255 = _T_1058 ? $signed(io_dataIn_bits_253) : $signed(buffers_0_63_1); // @[MuxLayer.scala 22:44]
  assign _GEN_256 = _T_1058 ? $signed(io_dataIn_bits_254) : $signed(buffers_0_63_2); // @[MuxLayer.scala 22:44]
  assign _GEN_257 = _T_1058 ? $signed(io_dataIn_bits_255) : $signed(buffers_0_63_3); // @[MuxLayer.scala 22:44]
  assign _T_1061 = cntr == 6'h3f; // @[MuxLayer.scala 29:15]
  assign _GEN_258 = _T_1061 ? 1'h1 : rdyReg; // @[MuxLayer.scala 29:36]
  assign _T_1063 = io_dataIn_valid & rdyReg; // @[MuxLayer.scala 32:26]
  assign _GEN_259 = _T_1063 ? 1'h0 : _GEN_258; // @[MuxLayer.scala 32:38]
  assign _T_1065 = cntr[1:0]; // @[MuxLayer.scala 45:19]
  assign _T_1068 = cntr[3:2]; // @[MuxLayer.scala 45:19]
  assign _T_1073 = cntr[5:4]; // @[MuxLayer.scala 45:19]
  assign _T_1090 = cntrs_0 == 2'h1; // @[MuxLayer.scala 55:25]
  assign _GEN_266 = _T_1090 ? $signed(buffers_0_1_0) : $signed(buffers_0_0_0); // @[MuxLayer.scala 55:35]
  assign _GEN_267 = _T_1090 ? $signed(buffers_0_1_1) : $signed(buffers_0_0_1); // @[MuxLayer.scala 55:35]
  assign _GEN_268 = _T_1090 ? $signed(buffers_0_1_2) : $signed(buffers_0_0_2); // @[MuxLayer.scala 55:35]
  assign _GEN_269 = _T_1090 ? $signed(buffers_0_1_3) : $signed(buffers_0_0_3); // @[MuxLayer.scala 55:35]
  assign _T_1092 = cntrs_0 == 2'h2; // @[MuxLayer.scala 55:25]
  assign _GEN_270 = _T_1092 ? $signed(buffers_0_2_0) : $signed(_GEN_266); // @[MuxLayer.scala 55:35]
  assign _GEN_271 = _T_1092 ? $signed(buffers_0_2_1) : $signed(_GEN_267); // @[MuxLayer.scala 55:35]
  assign _GEN_272 = _T_1092 ? $signed(buffers_0_2_2) : $signed(_GEN_268); // @[MuxLayer.scala 55:35]
  assign _GEN_273 = _T_1092 ? $signed(buffers_0_2_3) : $signed(_GEN_269); // @[MuxLayer.scala 55:35]
  assign _T_1094 = cntrs_0 == 2'h3; // @[MuxLayer.scala 55:25]
  assign _GEN_274 = _T_1094 ? $signed(buffers_0_3_0) : $signed(_GEN_270); // @[MuxLayer.scala 55:35]
  assign _GEN_275 = _T_1094 ? $signed(buffers_0_3_1) : $signed(_GEN_271); // @[MuxLayer.scala 55:35]
  assign _GEN_276 = _T_1094 ? $signed(buffers_0_3_2) : $signed(_GEN_272); // @[MuxLayer.scala 55:35]
  assign _GEN_277 = _T_1094 ? $signed(buffers_0_3_3) : $signed(_GEN_273); // @[MuxLayer.scala 55:35]
  assign _GEN_278 = _T_1090 ? $signed(buffers_0_5_0) : $signed(buffers_0_4_0); // @[MuxLayer.scala 55:35]
  assign _GEN_279 = _T_1090 ? $signed(buffers_0_5_1) : $signed(buffers_0_4_1); // @[MuxLayer.scala 55:35]
  assign _GEN_280 = _T_1090 ? $signed(buffers_0_5_2) : $signed(buffers_0_4_2); // @[MuxLayer.scala 55:35]
  assign _GEN_281 = _T_1090 ? $signed(buffers_0_5_3) : $signed(buffers_0_4_3); // @[MuxLayer.scala 55:35]
  assign _GEN_282 = _T_1092 ? $signed(buffers_0_6_0) : $signed(_GEN_278); // @[MuxLayer.scala 55:35]
  assign _GEN_283 = _T_1092 ? $signed(buffers_0_6_1) : $signed(_GEN_279); // @[MuxLayer.scala 55:35]
  assign _GEN_284 = _T_1092 ? $signed(buffers_0_6_2) : $signed(_GEN_280); // @[MuxLayer.scala 55:35]
  assign _GEN_285 = _T_1092 ? $signed(buffers_0_6_3) : $signed(_GEN_281); // @[MuxLayer.scala 55:35]
  assign _GEN_286 = _T_1094 ? $signed(buffers_0_7_0) : $signed(_GEN_282); // @[MuxLayer.scala 55:35]
  assign _GEN_287 = _T_1094 ? $signed(buffers_0_7_1) : $signed(_GEN_283); // @[MuxLayer.scala 55:35]
  assign _GEN_288 = _T_1094 ? $signed(buffers_0_7_2) : $signed(_GEN_284); // @[MuxLayer.scala 55:35]
  assign _GEN_289 = _T_1094 ? $signed(buffers_0_7_3) : $signed(_GEN_285); // @[MuxLayer.scala 55:35]
  assign _GEN_290 = _T_1090 ? $signed(buffers_0_9_0) : $signed(buffers_0_8_0); // @[MuxLayer.scala 55:35]
  assign _GEN_291 = _T_1090 ? $signed(buffers_0_9_1) : $signed(buffers_0_8_1); // @[MuxLayer.scala 55:35]
  assign _GEN_292 = _T_1090 ? $signed(buffers_0_9_2) : $signed(buffers_0_8_2); // @[MuxLayer.scala 55:35]
  assign _GEN_293 = _T_1090 ? $signed(buffers_0_9_3) : $signed(buffers_0_8_3); // @[MuxLayer.scala 55:35]
  assign _GEN_294 = _T_1092 ? $signed(buffers_0_10_0) : $signed(_GEN_290); // @[MuxLayer.scala 55:35]
  assign _GEN_295 = _T_1092 ? $signed(buffers_0_10_1) : $signed(_GEN_291); // @[MuxLayer.scala 55:35]
  assign _GEN_296 = _T_1092 ? $signed(buffers_0_10_2) : $signed(_GEN_292); // @[MuxLayer.scala 55:35]
  assign _GEN_297 = _T_1092 ? $signed(buffers_0_10_3) : $signed(_GEN_293); // @[MuxLayer.scala 55:35]
  assign _GEN_298 = _T_1094 ? $signed(buffers_0_11_0) : $signed(_GEN_294); // @[MuxLayer.scala 55:35]
  assign _GEN_299 = _T_1094 ? $signed(buffers_0_11_1) : $signed(_GEN_295); // @[MuxLayer.scala 55:35]
  assign _GEN_300 = _T_1094 ? $signed(buffers_0_11_2) : $signed(_GEN_296); // @[MuxLayer.scala 55:35]
  assign _GEN_301 = _T_1094 ? $signed(buffers_0_11_3) : $signed(_GEN_297); // @[MuxLayer.scala 55:35]
  assign _GEN_302 = _T_1090 ? $signed(buffers_0_13_0) : $signed(buffers_0_12_0); // @[MuxLayer.scala 55:35]
  assign _GEN_303 = _T_1090 ? $signed(buffers_0_13_1) : $signed(buffers_0_12_1); // @[MuxLayer.scala 55:35]
  assign _GEN_304 = _T_1090 ? $signed(buffers_0_13_2) : $signed(buffers_0_12_2); // @[MuxLayer.scala 55:35]
  assign _GEN_305 = _T_1090 ? $signed(buffers_0_13_3) : $signed(buffers_0_12_3); // @[MuxLayer.scala 55:35]
  assign _GEN_306 = _T_1092 ? $signed(buffers_0_14_0) : $signed(_GEN_302); // @[MuxLayer.scala 55:35]
  assign _GEN_307 = _T_1092 ? $signed(buffers_0_14_1) : $signed(_GEN_303); // @[MuxLayer.scala 55:35]
  assign _GEN_308 = _T_1092 ? $signed(buffers_0_14_2) : $signed(_GEN_304); // @[MuxLayer.scala 55:35]
  assign _GEN_309 = _T_1092 ? $signed(buffers_0_14_3) : $signed(_GEN_305); // @[MuxLayer.scala 55:35]
  assign _GEN_310 = _T_1094 ? $signed(buffers_0_15_0) : $signed(_GEN_306); // @[MuxLayer.scala 55:35]
  assign _GEN_311 = _T_1094 ? $signed(buffers_0_15_1) : $signed(_GEN_307); // @[MuxLayer.scala 55:35]
  assign _GEN_312 = _T_1094 ? $signed(buffers_0_15_2) : $signed(_GEN_308); // @[MuxLayer.scala 55:35]
  assign _GEN_313 = _T_1094 ? $signed(buffers_0_15_3) : $signed(_GEN_309); // @[MuxLayer.scala 55:35]
  assign _GEN_314 = _T_1090 ? $signed(buffers_0_17_0) : $signed(buffers_0_16_0); // @[MuxLayer.scala 55:35]
  assign _GEN_315 = _T_1090 ? $signed(buffers_0_17_1) : $signed(buffers_0_16_1); // @[MuxLayer.scala 55:35]
  assign _GEN_316 = _T_1090 ? $signed(buffers_0_17_2) : $signed(buffers_0_16_2); // @[MuxLayer.scala 55:35]
  assign _GEN_317 = _T_1090 ? $signed(buffers_0_17_3) : $signed(buffers_0_16_3); // @[MuxLayer.scala 55:35]
  assign _GEN_318 = _T_1092 ? $signed(buffers_0_18_0) : $signed(_GEN_314); // @[MuxLayer.scala 55:35]
  assign _GEN_319 = _T_1092 ? $signed(buffers_0_18_1) : $signed(_GEN_315); // @[MuxLayer.scala 55:35]
  assign _GEN_320 = _T_1092 ? $signed(buffers_0_18_2) : $signed(_GEN_316); // @[MuxLayer.scala 55:35]
  assign _GEN_321 = _T_1092 ? $signed(buffers_0_18_3) : $signed(_GEN_317); // @[MuxLayer.scala 55:35]
  assign _GEN_322 = _T_1094 ? $signed(buffers_0_19_0) : $signed(_GEN_318); // @[MuxLayer.scala 55:35]
  assign _GEN_323 = _T_1094 ? $signed(buffers_0_19_1) : $signed(_GEN_319); // @[MuxLayer.scala 55:35]
  assign _GEN_324 = _T_1094 ? $signed(buffers_0_19_2) : $signed(_GEN_320); // @[MuxLayer.scala 55:35]
  assign _GEN_325 = _T_1094 ? $signed(buffers_0_19_3) : $signed(_GEN_321); // @[MuxLayer.scala 55:35]
  assign _GEN_326 = _T_1090 ? $signed(buffers_0_21_0) : $signed(buffers_0_20_0); // @[MuxLayer.scala 55:35]
  assign _GEN_327 = _T_1090 ? $signed(buffers_0_21_1) : $signed(buffers_0_20_1); // @[MuxLayer.scala 55:35]
  assign _GEN_328 = _T_1090 ? $signed(buffers_0_21_2) : $signed(buffers_0_20_2); // @[MuxLayer.scala 55:35]
  assign _GEN_329 = _T_1090 ? $signed(buffers_0_21_3) : $signed(buffers_0_20_3); // @[MuxLayer.scala 55:35]
  assign _GEN_330 = _T_1092 ? $signed(buffers_0_22_0) : $signed(_GEN_326); // @[MuxLayer.scala 55:35]
  assign _GEN_331 = _T_1092 ? $signed(buffers_0_22_1) : $signed(_GEN_327); // @[MuxLayer.scala 55:35]
  assign _GEN_332 = _T_1092 ? $signed(buffers_0_22_2) : $signed(_GEN_328); // @[MuxLayer.scala 55:35]
  assign _GEN_333 = _T_1092 ? $signed(buffers_0_22_3) : $signed(_GEN_329); // @[MuxLayer.scala 55:35]
  assign _GEN_334 = _T_1094 ? $signed(buffers_0_23_0) : $signed(_GEN_330); // @[MuxLayer.scala 55:35]
  assign _GEN_335 = _T_1094 ? $signed(buffers_0_23_1) : $signed(_GEN_331); // @[MuxLayer.scala 55:35]
  assign _GEN_336 = _T_1094 ? $signed(buffers_0_23_2) : $signed(_GEN_332); // @[MuxLayer.scala 55:35]
  assign _GEN_337 = _T_1094 ? $signed(buffers_0_23_3) : $signed(_GEN_333); // @[MuxLayer.scala 55:35]
  assign _GEN_338 = _T_1090 ? $signed(buffers_0_25_0) : $signed(buffers_0_24_0); // @[MuxLayer.scala 55:35]
  assign _GEN_339 = _T_1090 ? $signed(buffers_0_25_1) : $signed(buffers_0_24_1); // @[MuxLayer.scala 55:35]
  assign _GEN_340 = _T_1090 ? $signed(buffers_0_25_2) : $signed(buffers_0_24_2); // @[MuxLayer.scala 55:35]
  assign _GEN_341 = _T_1090 ? $signed(buffers_0_25_3) : $signed(buffers_0_24_3); // @[MuxLayer.scala 55:35]
  assign _GEN_342 = _T_1092 ? $signed(buffers_0_26_0) : $signed(_GEN_338); // @[MuxLayer.scala 55:35]
  assign _GEN_343 = _T_1092 ? $signed(buffers_0_26_1) : $signed(_GEN_339); // @[MuxLayer.scala 55:35]
  assign _GEN_344 = _T_1092 ? $signed(buffers_0_26_2) : $signed(_GEN_340); // @[MuxLayer.scala 55:35]
  assign _GEN_345 = _T_1092 ? $signed(buffers_0_26_3) : $signed(_GEN_341); // @[MuxLayer.scala 55:35]
  assign _GEN_346 = _T_1094 ? $signed(buffers_0_27_0) : $signed(_GEN_342); // @[MuxLayer.scala 55:35]
  assign _GEN_347 = _T_1094 ? $signed(buffers_0_27_1) : $signed(_GEN_343); // @[MuxLayer.scala 55:35]
  assign _GEN_348 = _T_1094 ? $signed(buffers_0_27_2) : $signed(_GEN_344); // @[MuxLayer.scala 55:35]
  assign _GEN_349 = _T_1094 ? $signed(buffers_0_27_3) : $signed(_GEN_345); // @[MuxLayer.scala 55:35]
  assign _GEN_350 = _T_1090 ? $signed(buffers_0_29_0) : $signed(buffers_0_28_0); // @[MuxLayer.scala 55:35]
  assign _GEN_351 = _T_1090 ? $signed(buffers_0_29_1) : $signed(buffers_0_28_1); // @[MuxLayer.scala 55:35]
  assign _GEN_352 = _T_1090 ? $signed(buffers_0_29_2) : $signed(buffers_0_28_2); // @[MuxLayer.scala 55:35]
  assign _GEN_353 = _T_1090 ? $signed(buffers_0_29_3) : $signed(buffers_0_28_3); // @[MuxLayer.scala 55:35]
  assign _GEN_354 = _T_1092 ? $signed(buffers_0_30_0) : $signed(_GEN_350); // @[MuxLayer.scala 55:35]
  assign _GEN_355 = _T_1092 ? $signed(buffers_0_30_1) : $signed(_GEN_351); // @[MuxLayer.scala 55:35]
  assign _GEN_356 = _T_1092 ? $signed(buffers_0_30_2) : $signed(_GEN_352); // @[MuxLayer.scala 55:35]
  assign _GEN_357 = _T_1092 ? $signed(buffers_0_30_3) : $signed(_GEN_353); // @[MuxLayer.scala 55:35]
  assign _GEN_358 = _T_1094 ? $signed(buffers_0_31_0) : $signed(_GEN_354); // @[MuxLayer.scala 55:35]
  assign _GEN_359 = _T_1094 ? $signed(buffers_0_31_1) : $signed(_GEN_355); // @[MuxLayer.scala 55:35]
  assign _GEN_360 = _T_1094 ? $signed(buffers_0_31_2) : $signed(_GEN_356); // @[MuxLayer.scala 55:35]
  assign _GEN_361 = _T_1094 ? $signed(buffers_0_31_3) : $signed(_GEN_357); // @[MuxLayer.scala 55:35]
  assign _GEN_362 = _T_1090 ? $signed(buffers_0_33_0) : $signed(buffers_0_32_0); // @[MuxLayer.scala 55:35]
  assign _GEN_363 = _T_1090 ? $signed(buffers_0_33_1) : $signed(buffers_0_32_1); // @[MuxLayer.scala 55:35]
  assign _GEN_364 = _T_1090 ? $signed(buffers_0_33_2) : $signed(buffers_0_32_2); // @[MuxLayer.scala 55:35]
  assign _GEN_365 = _T_1090 ? $signed(buffers_0_33_3) : $signed(buffers_0_32_3); // @[MuxLayer.scala 55:35]
  assign _GEN_366 = _T_1092 ? $signed(buffers_0_34_0) : $signed(_GEN_362); // @[MuxLayer.scala 55:35]
  assign _GEN_367 = _T_1092 ? $signed(buffers_0_34_1) : $signed(_GEN_363); // @[MuxLayer.scala 55:35]
  assign _GEN_368 = _T_1092 ? $signed(buffers_0_34_2) : $signed(_GEN_364); // @[MuxLayer.scala 55:35]
  assign _GEN_369 = _T_1092 ? $signed(buffers_0_34_3) : $signed(_GEN_365); // @[MuxLayer.scala 55:35]
  assign _GEN_370 = _T_1094 ? $signed(buffers_0_35_0) : $signed(_GEN_366); // @[MuxLayer.scala 55:35]
  assign _GEN_371 = _T_1094 ? $signed(buffers_0_35_1) : $signed(_GEN_367); // @[MuxLayer.scala 55:35]
  assign _GEN_372 = _T_1094 ? $signed(buffers_0_35_2) : $signed(_GEN_368); // @[MuxLayer.scala 55:35]
  assign _GEN_373 = _T_1094 ? $signed(buffers_0_35_3) : $signed(_GEN_369); // @[MuxLayer.scala 55:35]
  assign _GEN_374 = _T_1090 ? $signed(buffers_0_37_0) : $signed(buffers_0_36_0); // @[MuxLayer.scala 55:35]
  assign _GEN_375 = _T_1090 ? $signed(buffers_0_37_1) : $signed(buffers_0_36_1); // @[MuxLayer.scala 55:35]
  assign _GEN_376 = _T_1090 ? $signed(buffers_0_37_2) : $signed(buffers_0_36_2); // @[MuxLayer.scala 55:35]
  assign _GEN_377 = _T_1090 ? $signed(buffers_0_37_3) : $signed(buffers_0_36_3); // @[MuxLayer.scala 55:35]
  assign _GEN_378 = _T_1092 ? $signed(buffers_0_38_0) : $signed(_GEN_374); // @[MuxLayer.scala 55:35]
  assign _GEN_379 = _T_1092 ? $signed(buffers_0_38_1) : $signed(_GEN_375); // @[MuxLayer.scala 55:35]
  assign _GEN_380 = _T_1092 ? $signed(buffers_0_38_2) : $signed(_GEN_376); // @[MuxLayer.scala 55:35]
  assign _GEN_381 = _T_1092 ? $signed(buffers_0_38_3) : $signed(_GEN_377); // @[MuxLayer.scala 55:35]
  assign _GEN_382 = _T_1094 ? $signed(buffers_0_39_0) : $signed(_GEN_378); // @[MuxLayer.scala 55:35]
  assign _GEN_383 = _T_1094 ? $signed(buffers_0_39_1) : $signed(_GEN_379); // @[MuxLayer.scala 55:35]
  assign _GEN_384 = _T_1094 ? $signed(buffers_0_39_2) : $signed(_GEN_380); // @[MuxLayer.scala 55:35]
  assign _GEN_385 = _T_1094 ? $signed(buffers_0_39_3) : $signed(_GEN_381); // @[MuxLayer.scala 55:35]
  assign _GEN_386 = _T_1090 ? $signed(buffers_0_41_0) : $signed(buffers_0_40_0); // @[MuxLayer.scala 55:35]
  assign _GEN_387 = _T_1090 ? $signed(buffers_0_41_1) : $signed(buffers_0_40_1); // @[MuxLayer.scala 55:35]
  assign _GEN_388 = _T_1090 ? $signed(buffers_0_41_2) : $signed(buffers_0_40_2); // @[MuxLayer.scala 55:35]
  assign _GEN_389 = _T_1090 ? $signed(buffers_0_41_3) : $signed(buffers_0_40_3); // @[MuxLayer.scala 55:35]
  assign _GEN_390 = _T_1092 ? $signed(buffers_0_42_0) : $signed(_GEN_386); // @[MuxLayer.scala 55:35]
  assign _GEN_391 = _T_1092 ? $signed(buffers_0_42_1) : $signed(_GEN_387); // @[MuxLayer.scala 55:35]
  assign _GEN_392 = _T_1092 ? $signed(buffers_0_42_2) : $signed(_GEN_388); // @[MuxLayer.scala 55:35]
  assign _GEN_393 = _T_1092 ? $signed(buffers_0_42_3) : $signed(_GEN_389); // @[MuxLayer.scala 55:35]
  assign _GEN_394 = _T_1094 ? $signed(buffers_0_43_0) : $signed(_GEN_390); // @[MuxLayer.scala 55:35]
  assign _GEN_395 = _T_1094 ? $signed(buffers_0_43_1) : $signed(_GEN_391); // @[MuxLayer.scala 55:35]
  assign _GEN_396 = _T_1094 ? $signed(buffers_0_43_2) : $signed(_GEN_392); // @[MuxLayer.scala 55:35]
  assign _GEN_397 = _T_1094 ? $signed(buffers_0_43_3) : $signed(_GEN_393); // @[MuxLayer.scala 55:35]
  assign _GEN_398 = _T_1090 ? $signed(buffers_0_45_0) : $signed(buffers_0_44_0); // @[MuxLayer.scala 55:35]
  assign _GEN_399 = _T_1090 ? $signed(buffers_0_45_1) : $signed(buffers_0_44_1); // @[MuxLayer.scala 55:35]
  assign _GEN_400 = _T_1090 ? $signed(buffers_0_45_2) : $signed(buffers_0_44_2); // @[MuxLayer.scala 55:35]
  assign _GEN_401 = _T_1090 ? $signed(buffers_0_45_3) : $signed(buffers_0_44_3); // @[MuxLayer.scala 55:35]
  assign _GEN_402 = _T_1092 ? $signed(buffers_0_46_0) : $signed(_GEN_398); // @[MuxLayer.scala 55:35]
  assign _GEN_403 = _T_1092 ? $signed(buffers_0_46_1) : $signed(_GEN_399); // @[MuxLayer.scala 55:35]
  assign _GEN_404 = _T_1092 ? $signed(buffers_0_46_2) : $signed(_GEN_400); // @[MuxLayer.scala 55:35]
  assign _GEN_405 = _T_1092 ? $signed(buffers_0_46_3) : $signed(_GEN_401); // @[MuxLayer.scala 55:35]
  assign _GEN_406 = _T_1094 ? $signed(buffers_0_47_0) : $signed(_GEN_402); // @[MuxLayer.scala 55:35]
  assign _GEN_407 = _T_1094 ? $signed(buffers_0_47_1) : $signed(_GEN_403); // @[MuxLayer.scala 55:35]
  assign _GEN_408 = _T_1094 ? $signed(buffers_0_47_2) : $signed(_GEN_404); // @[MuxLayer.scala 55:35]
  assign _GEN_409 = _T_1094 ? $signed(buffers_0_47_3) : $signed(_GEN_405); // @[MuxLayer.scala 55:35]
  assign _GEN_410 = _T_1090 ? $signed(buffers_0_49_0) : $signed(buffers_0_48_0); // @[MuxLayer.scala 55:35]
  assign _GEN_411 = _T_1090 ? $signed(buffers_0_49_1) : $signed(buffers_0_48_1); // @[MuxLayer.scala 55:35]
  assign _GEN_412 = _T_1090 ? $signed(buffers_0_49_2) : $signed(buffers_0_48_2); // @[MuxLayer.scala 55:35]
  assign _GEN_413 = _T_1090 ? $signed(buffers_0_49_3) : $signed(buffers_0_48_3); // @[MuxLayer.scala 55:35]
  assign _GEN_414 = _T_1092 ? $signed(buffers_0_50_0) : $signed(_GEN_410); // @[MuxLayer.scala 55:35]
  assign _GEN_415 = _T_1092 ? $signed(buffers_0_50_1) : $signed(_GEN_411); // @[MuxLayer.scala 55:35]
  assign _GEN_416 = _T_1092 ? $signed(buffers_0_50_2) : $signed(_GEN_412); // @[MuxLayer.scala 55:35]
  assign _GEN_417 = _T_1092 ? $signed(buffers_0_50_3) : $signed(_GEN_413); // @[MuxLayer.scala 55:35]
  assign _GEN_418 = _T_1094 ? $signed(buffers_0_51_0) : $signed(_GEN_414); // @[MuxLayer.scala 55:35]
  assign _GEN_419 = _T_1094 ? $signed(buffers_0_51_1) : $signed(_GEN_415); // @[MuxLayer.scala 55:35]
  assign _GEN_420 = _T_1094 ? $signed(buffers_0_51_2) : $signed(_GEN_416); // @[MuxLayer.scala 55:35]
  assign _GEN_421 = _T_1094 ? $signed(buffers_0_51_3) : $signed(_GEN_417); // @[MuxLayer.scala 55:35]
  assign _GEN_422 = _T_1090 ? $signed(buffers_0_53_0) : $signed(buffers_0_52_0); // @[MuxLayer.scala 55:35]
  assign _GEN_423 = _T_1090 ? $signed(buffers_0_53_1) : $signed(buffers_0_52_1); // @[MuxLayer.scala 55:35]
  assign _GEN_424 = _T_1090 ? $signed(buffers_0_53_2) : $signed(buffers_0_52_2); // @[MuxLayer.scala 55:35]
  assign _GEN_425 = _T_1090 ? $signed(buffers_0_53_3) : $signed(buffers_0_52_3); // @[MuxLayer.scala 55:35]
  assign _GEN_426 = _T_1092 ? $signed(buffers_0_54_0) : $signed(_GEN_422); // @[MuxLayer.scala 55:35]
  assign _GEN_427 = _T_1092 ? $signed(buffers_0_54_1) : $signed(_GEN_423); // @[MuxLayer.scala 55:35]
  assign _GEN_428 = _T_1092 ? $signed(buffers_0_54_2) : $signed(_GEN_424); // @[MuxLayer.scala 55:35]
  assign _GEN_429 = _T_1092 ? $signed(buffers_0_54_3) : $signed(_GEN_425); // @[MuxLayer.scala 55:35]
  assign _GEN_430 = _T_1094 ? $signed(buffers_0_55_0) : $signed(_GEN_426); // @[MuxLayer.scala 55:35]
  assign _GEN_431 = _T_1094 ? $signed(buffers_0_55_1) : $signed(_GEN_427); // @[MuxLayer.scala 55:35]
  assign _GEN_432 = _T_1094 ? $signed(buffers_0_55_2) : $signed(_GEN_428); // @[MuxLayer.scala 55:35]
  assign _GEN_433 = _T_1094 ? $signed(buffers_0_55_3) : $signed(_GEN_429); // @[MuxLayer.scala 55:35]
  assign _GEN_434 = _T_1090 ? $signed(buffers_0_57_0) : $signed(buffers_0_56_0); // @[MuxLayer.scala 55:35]
  assign _GEN_435 = _T_1090 ? $signed(buffers_0_57_1) : $signed(buffers_0_56_1); // @[MuxLayer.scala 55:35]
  assign _GEN_436 = _T_1090 ? $signed(buffers_0_57_2) : $signed(buffers_0_56_2); // @[MuxLayer.scala 55:35]
  assign _GEN_437 = _T_1090 ? $signed(buffers_0_57_3) : $signed(buffers_0_56_3); // @[MuxLayer.scala 55:35]
  assign _GEN_438 = _T_1092 ? $signed(buffers_0_58_0) : $signed(_GEN_434); // @[MuxLayer.scala 55:35]
  assign _GEN_439 = _T_1092 ? $signed(buffers_0_58_1) : $signed(_GEN_435); // @[MuxLayer.scala 55:35]
  assign _GEN_440 = _T_1092 ? $signed(buffers_0_58_2) : $signed(_GEN_436); // @[MuxLayer.scala 55:35]
  assign _GEN_441 = _T_1092 ? $signed(buffers_0_58_3) : $signed(_GEN_437); // @[MuxLayer.scala 55:35]
  assign _GEN_442 = _T_1094 ? $signed(buffers_0_59_0) : $signed(_GEN_438); // @[MuxLayer.scala 55:35]
  assign _GEN_443 = _T_1094 ? $signed(buffers_0_59_1) : $signed(_GEN_439); // @[MuxLayer.scala 55:35]
  assign _GEN_444 = _T_1094 ? $signed(buffers_0_59_2) : $signed(_GEN_440); // @[MuxLayer.scala 55:35]
  assign _GEN_445 = _T_1094 ? $signed(buffers_0_59_3) : $signed(_GEN_441); // @[MuxLayer.scala 55:35]
  assign _GEN_446 = _T_1090 ? $signed(buffers_0_61_0) : $signed(buffers_0_60_0); // @[MuxLayer.scala 55:35]
  assign _GEN_447 = _T_1090 ? $signed(buffers_0_61_1) : $signed(buffers_0_60_1); // @[MuxLayer.scala 55:35]
  assign _GEN_448 = _T_1090 ? $signed(buffers_0_61_2) : $signed(buffers_0_60_2); // @[MuxLayer.scala 55:35]
  assign _GEN_449 = _T_1090 ? $signed(buffers_0_61_3) : $signed(buffers_0_60_3); // @[MuxLayer.scala 55:35]
  assign _GEN_450 = _T_1092 ? $signed(buffers_0_62_0) : $signed(_GEN_446); // @[MuxLayer.scala 55:35]
  assign _GEN_451 = _T_1092 ? $signed(buffers_0_62_1) : $signed(_GEN_447); // @[MuxLayer.scala 55:35]
  assign _GEN_452 = _T_1092 ? $signed(buffers_0_62_2) : $signed(_GEN_448); // @[MuxLayer.scala 55:35]
  assign _GEN_453 = _T_1092 ? $signed(buffers_0_62_3) : $signed(_GEN_449); // @[MuxLayer.scala 55:35]
  assign _GEN_454 = _T_1094 ? $signed(buffers_0_63_0) : $signed(_GEN_450); // @[MuxLayer.scala 55:35]
  assign _GEN_455 = _T_1094 ? $signed(buffers_0_63_1) : $signed(_GEN_451); // @[MuxLayer.scala 55:35]
  assign _GEN_456 = _T_1094 ? $signed(buffers_0_63_2) : $signed(_GEN_452); // @[MuxLayer.scala 55:35]
  assign _GEN_457 = _T_1094 ? $signed(buffers_0_63_3) : $signed(_GEN_453); // @[MuxLayer.scala 55:35]
  assign _T_1778 = cntrs_1 == 2'h1; // @[MuxLayer.scala 55:25]
  assign _GEN_458 = _T_1778 ? $signed(buffers_1_1_0) : $signed(buffers_1_0_0); // @[MuxLayer.scala 55:35]
  assign _GEN_459 = _T_1778 ? $signed(buffers_1_1_1) : $signed(buffers_1_0_1); // @[MuxLayer.scala 55:35]
  assign _GEN_460 = _T_1778 ? $signed(buffers_1_1_2) : $signed(buffers_1_0_2); // @[MuxLayer.scala 55:35]
  assign _GEN_461 = _T_1778 ? $signed(buffers_1_1_3) : $signed(buffers_1_0_3); // @[MuxLayer.scala 55:35]
  assign _T_1780 = cntrs_1 == 2'h2; // @[MuxLayer.scala 55:25]
  assign _GEN_462 = _T_1780 ? $signed(buffers_1_2_0) : $signed(_GEN_458); // @[MuxLayer.scala 55:35]
  assign _GEN_463 = _T_1780 ? $signed(buffers_1_2_1) : $signed(_GEN_459); // @[MuxLayer.scala 55:35]
  assign _GEN_464 = _T_1780 ? $signed(buffers_1_2_2) : $signed(_GEN_460); // @[MuxLayer.scala 55:35]
  assign _GEN_465 = _T_1780 ? $signed(buffers_1_2_3) : $signed(_GEN_461); // @[MuxLayer.scala 55:35]
  assign _T_1782 = cntrs_1 == 2'h3; // @[MuxLayer.scala 55:25]
  assign _GEN_466 = _T_1782 ? $signed(buffers_1_3_0) : $signed(_GEN_462); // @[MuxLayer.scala 55:35]
  assign _GEN_467 = _T_1782 ? $signed(buffers_1_3_1) : $signed(_GEN_463); // @[MuxLayer.scala 55:35]
  assign _GEN_468 = _T_1782 ? $signed(buffers_1_3_2) : $signed(_GEN_464); // @[MuxLayer.scala 55:35]
  assign _GEN_469 = _T_1782 ? $signed(buffers_1_3_3) : $signed(_GEN_465); // @[MuxLayer.scala 55:35]
  assign _GEN_470 = _T_1778 ? $signed(buffers_1_5_0) : $signed(buffers_1_4_0); // @[MuxLayer.scala 55:35]
  assign _GEN_471 = _T_1778 ? $signed(buffers_1_5_1) : $signed(buffers_1_4_1); // @[MuxLayer.scala 55:35]
  assign _GEN_472 = _T_1778 ? $signed(buffers_1_5_2) : $signed(buffers_1_4_2); // @[MuxLayer.scala 55:35]
  assign _GEN_473 = _T_1778 ? $signed(buffers_1_5_3) : $signed(buffers_1_4_3); // @[MuxLayer.scala 55:35]
  assign _GEN_474 = _T_1780 ? $signed(buffers_1_6_0) : $signed(_GEN_470); // @[MuxLayer.scala 55:35]
  assign _GEN_475 = _T_1780 ? $signed(buffers_1_6_1) : $signed(_GEN_471); // @[MuxLayer.scala 55:35]
  assign _GEN_476 = _T_1780 ? $signed(buffers_1_6_2) : $signed(_GEN_472); // @[MuxLayer.scala 55:35]
  assign _GEN_477 = _T_1780 ? $signed(buffers_1_6_3) : $signed(_GEN_473); // @[MuxLayer.scala 55:35]
  assign _GEN_478 = _T_1782 ? $signed(buffers_1_7_0) : $signed(_GEN_474); // @[MuxLayer.scala 55:35]
  assign _GEN_479 = _T_1782 ? $signed(buffers_1_7_1) : $signed(_GEN_475); // @[MuxLayer.scala 55:35]
  assign _GEN_480 = _T_1782 ? $signed(buffers_1_7_2) : $signed(_GEN_476); // @[MuxLayer.scala 55:35]
  assign _GEN_481 = _T_1782 ? $signed(buffers_1_7_3) : $signed(_GEN_477); // @[MuxLayer.scala 55:35]
  assign _GEN_482 = _T_1778 ? $signed(buffers_1_9_0) : $signed(buffers_1_8_0); // @[MuxLayer.scala 55:35]
  assign _GEN_483 = _T_1778 ? $signed(buffers_1_9_1) : $signed(buffers_1_8_1); // @[MuxLayer.scala 55:35]
  assign _GEN_484 = _T_1778 ? $signed(buffers_1_9_2) : $signed(buffers_1_8_2); // @[MuxLayer.scala 55:35]
  assign _GEN_485 = _T_1778 ? $signed(buffers_1_9_3) : $signed(buffers_1_8_3); // @[MuxLayer.scala 55:35]
  assign _GEN_486 = _T_1780 ? $signed(buffers_1_10_0) : $signed(_GEN_482); // @[MuxLayer.scala 55:35]
  assign _GEN_487 = _T_1780 ? $signed(buffers_1_10_1) : $signed(_GEN_483); // @[MuxLayer.scala 55:35]
  assign _GEN_488 = _T_1780 ? $signed(buffers_1_10_2) : $signed(_GEN_484); // @[MuxLayer.scala 55:35]
  assign _GEN_489 = _T_1780 ? $signed(buffers_1_10_3) : $signed(_GEN_485); // @[MuxLayer.scala 55:35]
  assign _GEN_490 = _T_1782 ? $signed(buffers_1_11_0) : $signed(_GEN_486); // @[MuxLayer.scala 55:35]
  assign _GEN_491 = _T_1782 ? $signed(buffers_1_11_1) : $signed(_GEN_487); // @[MuxLayer.scala 55:35]
  assign _GEN_492 = _T_1782 ? $signed(buffers_1_11_2) : $signed(_GEN_488); // @[MuxLayer.scala 55:35]
  assign _GEN_493 = _T_1782 ? $signed(buffers_1_11_3) : $signed(_GEN_489); // @[MuxLayer.scala 55:35]
  assign _GEN_494 = _T_1778 ? $signed(buffers_1_13_0) : $signed(buffers_1_12_0); // @[MuxLayer.scala 55:35]
  assign _GEN_495 = _T_1778 ? $signed(buffers_1_13_1) : $signed(buffers_1_12_1); // @[MuxLayer.scala 55:35]
  assign _GEN_496 = _T_1778 ? $signed(buffers_1_13_2) : $signed(buffers_1_12_2); // @[MuxLayer.scala 55:35]
  assign _GEN_497 = _T_1778 ? $signed(buffers_1_13_3) : $signed(buffers_1_12_3); // @[MuxLayer.scala 55:35]
  assign _GEN_498 = _T_1780 ? $signed(buffers_1_14_0) : $signed(_GEN_494); // @[MuxLayer.scala 55:35]
  assign _GEN_499 = _T_1780 ? $signed(buffers_1_14_1) : $signed(_GEN_495); // @[MuxLayer.scala 55:35]
  assign _GEN_500 = _T_1780 ? $signed(buffers_1_14_2) : $signed(_GEN_496); // @[MuxLayer.scala 55:35]
  assign _GEN_501 = _T_1780 ? $signed(buffers_1_14_3) : $signed(_GEN_497); // @[MuxLayer.scala 55:35]
  assign _GEN_502 = _T_1782 ? $signed(buffers_1_15_0) : $signed(_GEN_498); // @[MuxLayer.scala 55:35]
  assign _GEN_503 = _T_1782 ? $signed(buffers_1_15_1) : $signed(_GEN_499); // @[MuxLayer.scala 55:35]
  assign _GEN_504 = _T_1782 ? $signed(buffers_1_15_2) : $signed(_GEN_500); // @[MuxLayer.scala 55:35]
  assign _GEN_505 = _T_1782 ? $signed(buffers_1_15_3) : $signed(_GEN_501); // @[MuxLayer.scala 55:35]
  assign _T_1950 = cntrs_2 == 2'h1; // @[MuxLayer.scala 55:25]
  assign _GEN_506 = _T_1950 ? $signed(buffers_2_1_0) : $signed(buffers_2_0_0); // @[MuxLayer.scala 55:35]
  assign _GEN_507 = _T_1950 ? $signed(buffers_2_1_1) : $signed(buffers_2_0_1); // @[MuxLayer.scala 55:35]
  assign _GEN_508 = _T_1950 ? $signed(buffers_2_1_2) : $signed(buffers_2_0_2); // @[MuxLayer.scala 55:35]
  assign _GEN_509 = _T_1950 ? $signed(buffers_2_1_3) : $signed(buffers_2_0_3); // @[MuxLayer.scala 55:35]
  assign _T_1952 = cntrs_2 == 2'h2; // @[MuxLayer.scala 55:25]
  assign _GEN_510 = _T_1952 ? $signed(buffers_2_2_0) : $signed(_GEN_506); // @[MuxLayer.scala 55:35]
  assign _GEN_511 = _T_1952 ? $signed(buffers_2_2_1) : $signed(_GEN_507); // @[MuxLayer.scala 55:35]
  assign _GEN_512 = _T_1952 ? $signed(buffers_2_2_2) : $signed(_GEN_508); // @[MuxLayer.scala 55:35]
  assign _GEN_513 = _T_1952 ? $signed(buffers_2_2_3) : $signed(_GEN_509); // @[MuxLayer.scala 55:35]
  assign _T_1954 = cntrs_2 == 2'h3; // @[MuxLayer.scala 55:25]
  assign _GEN_514 = _T_1954 ? $signed(buffers_2_3_0) : $signed(_GEN_510); // @[MuxLayer.scala 55:35]
  assign _GEN_515 = _T_1954 ? $signed(buffers_2_3_1) : $signed(_GEN_511); // @[MuxLayer.scala 55:35]
  assign _GEN_516 = _T_1954 ? $signed(buffers_2_3_2) : $signed(_GEN_512); // @[MuxLayer.scala 55:35]
  assign _GEN_517 = _T_1954 ? $signed(buffers_2_3_3) : $signed(_GEN_513); // @[MuxLayer.scala 55:35]
  assign _T_1994 = vld | lastVld; // @[MuxLayer.scala 68:27]
  assign io_dataIn_ready = rdyReg;
  assign io_dataOut_valid = _T_1994;
  assign io_dataOut_bits_0 = buffers_3_0_0;
  assign io_dataOut_bits_1 = buffers_3_0_1;
  assign io_dataOut_bits_2 = buffers_3_0_2;
  assign io_dataOut_bits_3 = buffers_3_0_3;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  rdyReg = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  cntr = _RAND_1[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  buffers_0_0_0 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  buffers_0_0_1 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  buffers_0_0_2 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  buffers_0_0_3 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  buffers_0_1_0 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  buffers_0_1_1 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  buffers_0_1_2 = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  buffers_0_1_3 = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  buffers_0_2_0 = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  buffers_0_2_1 = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  buffers_0_2_2 = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  buffers_0_2_3 = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  buffers_0_3_0 = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  buffers_0_3_1 = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  buffers_0_3_2 = _RAND_16[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  buffers_0_3_3 = _RAND_17[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  buffers_0_4_0 = _RAND_18[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  buffers_0_4_1 = _RAND_19[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  buffers_0_4_2 = _RAND_20[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  buffers_0_4_3 = _RAND_21[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  buffers_0_5_0 = _RAND_22[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  buffers_0_5_1 = _RAND_23[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  buffers_0_5_2 = _RAND_24[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  buffers_0_5_3 = _RAND_25[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  buffers_0_6_0 = _RAND_26[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  buffers_0_6_1 = _RAND_27[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  buffers_0_6_2 = _RAND_28[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  buffers_0_6_3 = _RAND_29[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  buffers_0_7_0 = _RAND_30[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  buffers_0_7_1 = _RAND_31[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  buffers_0_7_2 = _RAND_32[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{$random}};
  buffers_0_7_3 = _RAND_33[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{$random}};
  buffers_0_8_0 = _RAND_34[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{$random}};
  buffers_0_8_1 = _RAND_35[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{$random}};
  buffers_0_8_2 = _RAND_36[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{$random}};
  buffers_0_8_3 = _RAND_37[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{$random}};
  buffers_0_9_0 = _RAND_38[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{$random}};
  buffers_0_9_1 = _RAND_39[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{$random}};
  buffers_0_9_2 = _RAND_40[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{$random}};
  buffers_0_9_3 = _RAND_41[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{$random}};
  buffers_0_10_0 = _RAND_42[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{$random}};
  buffers_0_10_1 = _RAND_43[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{$random}};
  buffers_0_10_2 = _RAND_44[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{$random}};
  buffers_0_10_3 = _RAND_45[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{$random}};
  buffers_0_11_0 = _RAND_46[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{$random}};
  buffers_0_11_1 = _RAND_47[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{$random}};
  buffers_0_11_2 = _RAND_48[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{$random}};
  buffers_0_11_3 = _RAND_49[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{$random}};
  buffers_0_12_0 = _RAND_50[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{$random}};
  buffers_0_12_1 = _RAND_51[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{$random}};
  buffers_0_12_2 = _RAND_52[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{$random}};
  buffers_0_12_3 = _RAND_53[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{$random}};
  buffers_0_13_0 = _RAND_54[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{$random}};
  buffers_0_13_1 = _RAND_55[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{$random}};
  buffers_0_13_2 = _RAND_56[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{$random}};
  buffers_0_13_3 = _RAND_57[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{$random}};
  buffers_0_14_0 = _RAND_58[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{$random}};
  buffers_0_14_1 = _RAND_59[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{$random}};
  buffers_0_14_2 = _RAND_60[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{$random}};
  buffers_0_14_3 = _RAND_61[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{$random}};
  buffers_0_15_0 = _RAND_62[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{$random}};
  buffers_0_15_1 = _RAND_63[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{$random}};
  buffers_0_15_2 = _RAND_64[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{$random}};
  buffers_0_15_3 = _RAND_65[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{$random}};
  buffers_0_16_0 = _RAND_66[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{$random}};
  buffers_0_16_1 = _RAND_67[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{$random}};
  buffers_0_16_2 = _RAND_68[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{$random}};
  buffers_0_16_3 = _RAND_69[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{$random}};
  buffers_0_17_0 = _RAND_70[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{$random}};
  buffers_0_17_1 = _RAND_71[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{$random}};
  buffers_0_17_2 = _RAND_72[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{$random}};
  buffers_0_17_3 = _RAND_73[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{$random}};
  buffers_0_18_0 = _RAND_74[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{$random}};
  buffers_0_18_1 = _RAND_75[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{$random}};
  buffers_0_18_2 = _RAND_76[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{$random}};
  buffers_0_18_3 = _RAND_77[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{$random}};
  buffers_0_19_0 = _RAND_78[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{$random}};
  buffers_0_19_1 = _RAND_79[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{$random}};
  buffers_0_19_2 = _RAND_80[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{$random}};
  buffers_0_19_3 = _RAND_81[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{$random}};
  buffers_0_20_0 = _RAND_82[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{$random}};
  buffers_0_20_1 = _RAND_83[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{$random}};
  buffers_0_20_2 = _RAND_84[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{$random}};
  buffers_0_20_3 = _RAND_85[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{$random}};
  buffers_0_21_0 = _RAND_86[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{$random}};
  buffers_0_21_1 = _RAND_87[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{$random}};
  buffers_0_21_2 = _RAND_88[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{$random}};
  buffers_0_21_3 = _RAND_89[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{$random}};
  buffers_0_22_0 = _RAND_90[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{$random}};
  buffers_0_22_1 = _RAND_91[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{$random}};
  buffers_0_22_2 = _RAND_92[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{$random}};
  buffers_0_22_3 = _RAND_93[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{$random}};
  buffers_0_23_0 = _RAND_94[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{$random}};
  buffers_0_23_1 = _RAND_95[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{$random}};
  buffers_0_23_2 = _RAND_96[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{$random}};
  buffers_0_23_3 = _RAND_97[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{$random}};
  buffers_0_24_0 = _RAND_98[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{$random}};
  buffers_0_24_1 = _RAND_99[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{$random}};
  buffers_0_24_2 = _RAND_100[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{$random}};
  buffers_0_24_3 = _RAND_101[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{$random}};
  buffers_0_25_0 = _RAND_102[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{$random}};
  buffers_0_25_1 = _RAND_103[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{$random}};
  buffers_0_25_2 = _RAND_104[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{$random}};
  buffers_0_25_3 = _RAND_105[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{$random}};
  buffers_0_26_0 = _RAND_106[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{$random}};
  buffers_0_26_1 = _RAND_107[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{$random}};
  buffers_0_26_2 = _RAND_108[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{$random}};
  buffers_0_26_3 = _RAND_109[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{$random}};
  buffers_0_27_0 = _RAND_110[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{$random}};
  buffers_0_27_1 = _RAND_111[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{$random}};
  buffers_0_27_2 = _RAND_112[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{$random}};
  buffers_0_27_3 = _RAND_113[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{$random}};
  buffers_0_28_0 = _RAND_114[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{$random}};
  buffers_0_28_1 = _RAND_115[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{$random}};
  buffers_0_28_2 = _RAND_116[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{$random}};
  buffers_0_28_3 = _RAND_117[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{$random}};
  buffers_0_29_0 = _RAND_118[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{$random}};
  buffers_0_29_1 = _RAND_119[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{$random}};
  buffers_0_29_2 = _RAND_120[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{$random}};
  buffers_0_29_3 = _RAND_121[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{$random}};
  buffers_0_30_0 = _RAND_122[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{$random}};
  buffers_0_30_1 = _RAND_123[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{$random}};
  buffers_0_30_2 = _RAND_124[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{$random}};
  buffers_0_30_3 = _RAND_125[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{$random}};
  buffers_0_31_0 = _RAND_126[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{$random}};
  buffers_0_31_1 = _RAND_127[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{$random}};
  buffers_0_31_2 = _RAND_128[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{$random}};
  buffers_0_31_3 = _RAND_129[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{$random}};
  buffers_0_32_0 = _RAND_130[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{$random}};
  buffers_0_32_1 = _RAND_131[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{$random}};
  buffers_0_32_2 = _RAND_132[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{$random}};
  buffers_0_32_3 = _RAND_133[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{$random}};
  buffers_0_33_0 = _RAND_134[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{$random}};
  buffers_0_33_1 = _RAND_135[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{$random}};
  buffers_0_33_2 = _RAND_136[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{$random}};
  buffers_0_33_3 = _RAND_137[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{$random}};
  buffers_0_34_0 = _RAND_138[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{$random}};
  buffers_0_34_1 = _RAND_139[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{$random}};
  buffers_0_34_2 = _RAND_140[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{$random}};
  buffers_0_34_3 = _RAND_141[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{$random}};
  buffers_0_35_0 = _RAND_142[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{$random}};
  buffers_0_35_1 = _RAND_143[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{$random}};
  buffers_0_35_2 = _RAND_144[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{$random}};
  buffers_0_35_3 = _RAND_145[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{$random}};
  buffers_0_36_0 = _RAND_146[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{$random}};
  buffers_0_36_1 = _RAND_147[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{$random}};
  buffers_0_36_2 = _RAND_148[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{$random}};
  buffers_0_36_3 = _RAND_149[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{$random}};
  buffers_0_37_0 = _RAND_150[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{$random}};
  buffers_0_37_1 = _RAND_151[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{$random}};
  buffers_0_37_2 = _RAND_152[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{$random}};
  buffers_0_37_3 = _RAND_153[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{$random}};
  buffers_0_38_0 = _RAND_154[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{$random}};
  buffers_0_38_1 = _RAND_155[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{$random}};
  buffers_0_38_2 = _RAND_156[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{$random}};
  buffers_0_38_3 = _RAND_157[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{$random}};
  buffers_0_39_0 = _RAND_158[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{$random}};
  buffers_0_39_1 = _RAND_159[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{$random}};
  buffers_0_39_2 = _RAND_160[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{$random}};
  buffers_0_39_3 = _RAND_161[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{$random}};
  buffers_0_40_0 = _RAND_162[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{$random}};
  buffers_0_40_1 = _RAND_163[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{$random}};
  buffers_0_40_2 = _RAND_164[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{$random}};
  buffers_0_40_3 = _RAND_165[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{$random}};
  buffers_0_41_0 = _RAND_166[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{$random}};
  buffers_0_41_1 = _RAND_167[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{$random}};
  buffers_0_41_2 = _RAND_168[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{$random}};
  buffers_0_41_3 = _RAND_169[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{$random}};
  buffers_0_42_0 = _RAND_170[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{$random}};
  buffers_0_42_1 = _RAND_171[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{$random}};
  buffers_0_42_2 = _RAND_172[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{$random}};
  buffers_0_42_3 = _RAND_173[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{$random}};
  buffers_0_43_0 = _RAND_174[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{$random}};
  buffers_0_43_1 = _RAND_175[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{$random}};
  buffers_0_43_2 = _RAND_176[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{$random}};
  buffers_0_43_3 = _RAND_177[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{$random}};
  buffers_0_44_0 = _RAND_178[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{$random}};
  buffers_0_44_1 = _RAND_179[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{$random}};
  buffers_0_44_2 = _RAND_180[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{$random}};
  buffers_0_44_3 = _RAND_181[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{$random}};
  buffers_0_45_0 = _RAND_182[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{$random}};
  buffers_0_45_1 = _RAND_183[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{$random}};
  buffers_0_45_2 = _RAND_184[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{$random}};
  buffers_0_45_3 = _RAND_185[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{$random}};
  buffers_0_46_0 = _RAND_186[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{$random}};
  buffers_0_46_1 = _RAND_187[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{$random}};
  buffers_0_46_2 = _RAND_188[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{$random}};
  buffers_0_46_3 = _RAND_189[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{$random}};
  buffers_0_47_0 = _RAND_190[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{$random}};
  buffers_0_47_1 = _RAND_191[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{$random}};
  buffers_0_47_2 = _RAND_192[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{$random}};
  buffers_0_47_3 = _RAND_193[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{$random}};
  buffers_0_48_0 = _RAND_194[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{$random}};
  buffers_0_48_1 = _RAND_195[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{$random}};
  buffers_0_48_2 = _RAND_196[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{$random}};
  buffers_0_48_3 = _RAND_197[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{$random}};
  buffers_0_49_0 = _RAND_198[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{$random}};
  buffers_0_49_1 = _RAND_199[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{$random}};
  buffers_0_49_2 = _RAND_200[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{$random}};
  buffers_0_49_3 = _RAND_201[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{$random}};
  buffers_0_50_0 = _RAND_202[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{$random}};
  buffers_0_50_1 = _RAND_203[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{$random}};
  buffers_0_50_2 = _RAND_204[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{$random}};
  buffers_0_50_3 = _RAND_205[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{$random}};
  buffers_0_51_0 = _RAND_206[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{$random}};
  buffers_0_51_1 = _RAND_207[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{$random}};
  buffers_0_51_2 = _RAND_208[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{$random}};
  buffers_0_51_3 = _RAND_209[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{$random}};
  buffers_0_52_0 = _RAND_210[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{$random}};
  buffers_0_52_1 = _RAND_211[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{$random}};
  buffers_0_52_2 = _RAND_212[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{$random}};
  buffers_0_52_3 = _RAND_213[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{$random}};
  buffers_0_53_0 = _RAND_214[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{$random}};
  buffers_0_53_1 = _RAND_215[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{$random}};
  buffers_0_53_2 = _RAND_216[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{$random}};
  buffers_0_53_3 = _RAND_217[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{$random}};
  buffers_0_54_0 = _RAND_218[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{$random}};
  buffers_0_54_1 = _RAND_219[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{$random}};
  buffers_0_54_2 = _RAND_220[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{$random}};
  buffers_0_54_3 = _RAND_221[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{$random}};
  buffers_0_55_0 = _RAND_222[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{$random}};
  buffers_0_55_1 = _RAND_223[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{$random}};
  buffers_0_55_2 = _RAND_224[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{$random}};
  buffers_0_55_3 = _RAND_225[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{$random}};
  buffers_0_56_0 = _RAND_226[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{$random}};
  buffers_0_56_1 = _RAND_227[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{$random}};
  buffers_0_56_2 = _RAND_228[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{$random}};
  buffers_0_56_3 = _RAND_229[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{$random}};
  buffers_0_57_0 = _RAND_230[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{$random}};
  buffers_0_57_1 = _RAND_231[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{$random}};
  buffers_0_57_2 = _RAND_232[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{$random}};
  buffers_0_57_3 = _RAND_233[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{$random}};
  buffers_0_58_0 = _RAND_234[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{$random}};
  buffers_0_58_1 = _RAND_235[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{$random}};
  buffers_0_58_2 = _RAND_236[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{$random}};
  buffers_0_58_3 = _RAND_237[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{$random}};
  buffers_0_59_0 = _RAND_238[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{$random}};
  buffers_0_59_1 = _RAND_239[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{$random}};
  buffers_0_59_2 = _RAND_240[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{$random}};
  buffers_0_59_3 = _RAND_241[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{$random}};
  buffers_0_60_0 = _RAND_242[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{$random}};
  buffers_0_60_1 = _RAND_243[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{$random}};
  buffers_0_60_2 = _RAND_244[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{$random}};
  buffers_0_60_3 = _RAND_245[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{$random}};
  buffers_0_61_0 = _RAND_246[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{$random}};
  buffers_0_61_1 = _RAND_247[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{$random}};
  buffers_0_61_2 = _RAND_248[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{$random}};
  buffers_0_61_3 = _RAND_249[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{$random}};
  buffers_0_62_0 = _RAND_250[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{$random}};
  buffers_0_62_1 = _RAND_251[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{$random}};
  buffers_0_62_2 = _RAND_252[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{$random}};
  buffers_0_62_3 = _RAND_253[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{$random}};
  buffers_0_63_0 = _RAND_254[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{$random}};
  buffers_0_63_1 = _RAND_255[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{$random}};
  buffers_0_63_2 = _RAND_256[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{$random}};
  buffers_0_63_3 = _RAND_257[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{$random}};
  cntrs_0 = _RAND_258[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{$random}};
  _T_1071 = _RAND_259[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{$random}};
  cntrs_1 = _RAND_260[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{$random}};
  _T_1076 = _RAND_261[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{$random}};
  _T_1078 = _RAND_262[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{$random}};
  cntrs_2 = _RAND_263[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{$random}};
  buffers_1_0_0 = _RAND_264[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{$random}};
  buffers_1_0_1 = _RAND_265[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{$random}};
  buffers_1_0_2 = _RAND_266[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{$random}};
  buffers_1_0_3 = _RAND_267[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{$random}};
  buffers_1_1_0 = _RAND_268[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{$random}};
  buffers_1_1_1 = _RAND_269[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{$random}};
  buffers_1_1_2 = _RAND_270[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{$random}};
  buffers_1_1_3 = _RAND_271[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{$random}};
  buffers_1_2_0 = _RAND_272[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{$random}};
  buffers_1_2_1 = _RAND_273[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{$random}};
  buffers_1_2_2 = _RAND_274[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{$random}};
  buffers_1_2_3 = _RAND_275[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{$random}};
  buffers_1_3_0 = _RAND_276[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{$random}};
  buffers_1_3_1 = _RAND_277[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{$random}};
  buffers_1_3_2 = _RAND_278[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{$random}};
  buffers_1_3_3 = _RAND_279[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{$random}};
  buffers_1_4_0 = _RAND_280[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{$random}};
  buffers_1_4_1 = _RAND_281[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{$random}};
  buffers_1_4_2 = _RAND_282[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{$random}};
  buffers_1_4_3 = _RAND_283[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{$random}};
  buffers_1_5_0 = _RAND_284[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{$random}};
  buffers_1_5_1 = _RAND_285[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{$random}};
  buffers_1_5_2 = _RAND_286[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{$random}};
  buffers_1_5_3 = _RAND_287[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{$random}};
  buffers_1_6_0 = _RAND_288[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{$random}};
  buffers_1_6_1 = _RAND_289[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{$random}};
  buffers_1_6_2 = _RAND_290[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{$random}};
  buffers_1_6_3 = _RAND_291[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{$random}};
  buffers_1_7_0 = _RAND_292[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{$random}};
  buffers_1_7_1 = _RAND_293[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{$random}};
  buffers_1_7_2 = _RAND_294[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{$random}};
  buffers_1_7_3 = _RAND_295[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{$random}};
  buffers_1_8_0 = _RAND_296[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{$random}};
  buffers_1_8_1 = _RAND_297[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{$random}};
  buffers_1_8_2 = _RAND_298[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{$random}};
  buffers_1_8_3 = _RAND_299[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{$random}};
  buffers_1_9_0 = _RAND_300[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{$random}};
  buffers_1_9_1 = _RAND_301[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{$random}};
  buffers_1_9_2 = _RAND_302[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{$random}};
  buffers_1_9_3 = _RAND_303[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{$random}};
  buffers_1_10_0 = _RAND_304[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{$random}};
  buffers_1_10_1 = _RAND_305[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{$random}};
  buffers_1_10_2 = _RAND_306[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{$random}};
  buffers_1_10_3 = _RAND_307[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{$random}};
  buffers_1_11_0 = _RAND_308[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{$random}};
  buffers_1_11_1 = _RAND_309[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{$random}};
  buffers_1_11_2 = _RAND_310[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{$random}};
  buffers_1_11_3 = _RAND_311[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{$random}};
  buffers_1_12_0 = _RAND_312[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{$random}};
  buffers_1_12_1 = _RAND_313[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{$random}};
  buffers_1_12_2 = _RAND_314[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{$random}};
  buffers_1_12_3 = _RAND_315[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{$random}};
  buffers_1_13_0 = _RAND_316[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{$random}};
  buffers_1_13_1 = _RAND_317[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{$random}};
  buffers_1_13_2 = _RAND_318[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{$random}};
  buffers_1_13_3 = _RAND_319[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{$random}};
  buffers_1_14_0 = _RAND_320[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{$random}};
  buffers_1_14_1 = _RAND_321[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{$random}};
  buffers_1_14_2 = _RAND_322[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{$random}};
  buffers_1_14_3 = _RAND_323[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{$random}};
  buffers_1_15_0 = _RAND_324[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{$random}};
  buffers_1_15_1 = _RAND_325[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{$random}};
  buffers_1_15_2 = _RAND_326[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{$random}};
  buffers_1_15_3 = _RAND_327[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{$random}};
  buffers_2_0_0 = _RAND_328[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{$random}};
  buffers_2_0_1 = _RAND_329[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{$random}};
  buffers_2_0_2 = _RAND_330[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{$random}};
  buffers_2_0_3 = _RAND_331[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{$random}};
  buffers_2_1_0 = _RAND_332[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{$random}};
  buffers_2_1_1 = _RAND_333[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{$random}};
  buffers_2_1_2 = _RAND_334[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{$random}};
  buffers_2_1_3 = _RAND_335[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{$random}};
  buffers_2_2_0 = _RAND_336[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{$random}};
  buffers_2_2_1 = _RAND_337[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{$random}};
  buffers_2_2_2 = _RAND_338[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{$random}};
  buffers_2_2_3 = _RAND_339[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{$random}};
  buffers_2_3_0 = _RAND_340[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{$random}};
  buffers_2_3_1 = _RAND_341[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{$random}};
  buffers_2_3_2 = _RAND_342[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{$random}};
  buffers_2_3_3 = _RAND_343[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{$random}};
  buffers_3_0_0 = _RAND_344[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{$random}};
  buffers_3_0_1 = _RAND_345[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{$random}};
  buffers_3_0_2 = _RAND_346[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{$random}};
  buffers_3_0_3 = _RAND_347[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{$random}};
  _T_1988 = _RAND_348[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{$random}};
  _T_1990 = _RAND_349[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{$random}};
  vld = _RAND_350[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{$random}};
  lastVld = _RAND_351[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      rdyReg <= 1'h1;
    end else begin
      if (_T_1063) begin
        rdyReg <= 1'h0;
      end else begin
        if (_T_1061) begin
          rdyReg <= 1'h1;
        end
      end
    end
    if (reset) begin
      cntr <= 6'h0;
    end else begin
      if (_T_1058) begin
        cntr <= 6'h1;
      end else begin
        if (_T_1052) begin
          cntr <= _T_1055;
        end
      end
    end
    if (_T_1058) begin
      buffers_0_0_0 <= io_dataIn_bits_0;
    end
    if (_T_1058) begin
      buffers_0_0_1 <= io_dataIn_bits_1;
    end
    if (_T_1058) begin
      buffers_0_0_2 <= io_dataIn_bits_2;
    end
    if (_T_1058) begin
      buffers_0_0_3 <= io_dataIn_bits_3;
    end
    if (_T_1058) begin
      buffers_0_1_0 <= io_dataIn_bits_4;
    end
    if (_T_1058) begin
      buffers_0_1_1 <= io_dataIn_bits_5;
    end
    if (_T_1058) begin
      buffers_0_1_2 <= io_dataIn_bits_6;
    end
    if (_T_1058) begin
      buffers_0_1_3 <= io_dataIn_bits_7;
    end
    if (_T_1058) begin
      buffers_0_2_0 <= io_dataIn_bits_8;
    end
    if (_T_1058) begin
      buffers_0_2_1 <= io_dataIn_bits_9;
    end
    if (_T_1058) begin
      buffers_0_2_2 <= io_dataIn_bits_10;
    end
    if (_T_1058) begin
      buffers_0_2_3 <= io_dataIn_bits_11;
    end
    if (_T_1058) begin
      buffers_0_3_0 <= io_dataIn_bits_12;
    end
    if (_T_1058) begin
      buffers_0_3_1 <= io_dataIn_bits_13;
    end
    if (_T_1058) begin
      buffers_0_3_2 <= io_dataIn_bits_14;
    end
    if (_T_1058) begin
      buffers_0_3_3 <= io_dataIn_bits_15;
    end
    if (_T_1058) begin
      buffers_0_4_0 <= io_dataIn_bits_16;
    end
    if (_T_1058) begin
      buffers_0_4_1 <= io_dataIn_bits_17;
    end
    if (_T_1058) begin
      buffers_0_4_2 <= io_dataIn_bits_18;
    end
    if (_T_1058) begin
      buffers_0_4_3 <= io_dataIn_bits_19;
    end
    if (_T_1058) begin
      buffers_0_5_0 <= io_dataIn_bits_20;
    end
    if (_T_1058) begin
      buffers_0_5_1 <= io_dataIn_bits_21;
    end
    if (_T_1058) begin
      buffers_0_5_2 <= io_dataIn_bits_22;
    end
    if (_T_1058) begin
      buffers_0_5_3 <= io_dataIn_bits_23;
    end
    if (_T_1058) begin
      buffers_0_6_0 <= io_dataIn_bits_24;
    end
    if (_T_1058) begin
      buffers_0_6_1 <= io_dataIn_bits_25;
    end
    if (_T_1058) begin
      buffers_0_6_2 <= io_dataIn_bits_26;
    end
    if (_T_1058) begin
      buffers_0_6_3 <= io_dataIn_bits_27;
    end
    if (_T_1058) begin
      buffers_0_7_0 <= io_dataIn_bits_28;
    end
    if (_T_1058) begin
      buffers_0_7_1 <= io_dataIn_bits_29;
    end
    if (_T_1058) begin
      buffers_0_7_2 <= io_dataIn_bits_30;
    end
    if (_T_1058) begin
      buffers_0_7_3 <= io_dataIn_bits_31;
    end
    if (_T_1058) begin
      buffers_0_8_0 <= io_dataIn_bits_32;
    end
    if (_T_1058) begin
      buffers_0_8_1 <= io_dataIn_bits_33;
    end
    if (_T_1058) begin
      buffers_0_8_2 <= io_dataIn_bits_34;
    end
    if (_T_1058) begin
      buffers_0_8_3 <= io_dataIn_bits_35;
    end
    if (_T_1058) begin
      buffers_0_9_0 <= io_dataIn_bits_36;
    end
    if (_T_1058) begin
      buffers_0_9_1 <= io_dataIn_bits_37;
    end
    if (_T_1058) begin
      buffers_0_9_2 <= io_dataIn_bits_38;
    end
    if (_T_1058) begin
      buffers_0_9_3 <= io_dataIn_bits_39;
    end
    if (_T_1058) begin
      buffers_0_10_0 <= io_dataIn_bits_40;
    end
    if (_T_1058) begin
      buffers_0_10_1 <= io_dataIn_bits_41;
    end
    if (_T_1058) begin
      buffers_0_10_2 <= io_dataIn_bits_42;
    end
    if (_T_1058) begin
      buffers_0_10_3 <= io_dataIn_bits_43;
    end
    if (_T_1058) begin
      buffers_0_11_0 <= io_dataIn_bits_44;
    end
    if (_T_1058) begin
      buffers_0_11_1 <= io_dataIn_bits_45;
    end
    if (_T_1058) begin
      buffers_0_11_2 <= io_dataIn_bits_46;
    end
    if (_T_1058) begin
      buffers_0_11_3 <= io_dataIn_bits_47;
    end
    if (_T_1058) begin
      buffers_0_12_0 <= io_dataIn_bits_48;
    end
    if (_T_1058) begin
      buffers_0_12_1 <= io_dataIn_bits_49;
    end
    if (_T_1058) begin
      buffers_0_12_2 <= io_dataIn_bits_50;
    end
    if (_T_1058) begin
      buffers_0_12_3 <= io_dataIn_bits_51;
    end
    if (_T_1058) begin
      buffers_0_13_0 <= io_dataIn_bits_52;
    end
    if (_T_1058) begin
      buffers_0_13_1 <= io_dataIn_bits_53;
    end
    if (_T_1058) begin
      buffers_0_13_2 <= io_dataIn_bits_54;
    end
    if (_T_1058) begin
      buffers_0_13_3 <= io_dataIn_bits_55;
    end
    if (_T_1058) begin
      buffers_0_14_0 <= io_dataIn_bits_56;
    end
    if (_T_1058) begin
      buffers_0_14_1 <= io_dataIn_bits_57;
    end
    if (_T_1058) begin
      buffers_0_14_2 <= io_dataIn_bits_58;
    end
    if (_T_1058) begin
      buffers_0_14_3 <= io_dataIn_bits_59;
    end
    if (_T_1058) begin
      buffers_0_15_0 <= io_dataIn_bits_60;
    end
    if (_T_1058) begin
      buffers_0_15_1 <= io_dataIn_bits_61;
    end
    if (_T_1058) begin
      buffers_0_15_2 <= io_dataIn_bits_62;
    end
    if (_T_1058) begin
      buffers_0_15_3 <= io_dataIn_bits_63;
    end
    if (_T_1058) begin
      buffers_0_16_0 <= io_dataIn_bits_64;
    end
    if (_T_1058) begin
      buffers_0_16_1 <= io_dataIn_bits_65;
    end
    if (_T_1058) begin
      buffers_0_16_2 <= io_dataIn_bits_66;
    end
    if (_T_1058) begin
      buffers_0_16_3 <= io_dataIn_bits_67;
    end
    if (_T_1058) begin
      buffers_0_17_0 <= io_dataIn_bits_68;
    end
    if (_T_1058) begin
      buffers_0_17_1 <= io_dataIn_bits_69;
    end
    if (_T_1058) begin
      buffers_0_17_2 <= io_dataIn_bits_70;
    end
    if (_T_1058) begin
      buffers_0_17_3 <= io_dataIn_bits_71;
    end
    if (_T_1058) begin
      buffers_0_18_0 <= io_dataIn_bits_72;
    end
    if (_T_1058) begin
      buffers_0_18_1 <= io_dataIn_bits_73;
    end
    if (_T_1058) begin
      buffers_0_18_2 <= io_dataIn_bits_74;
    end
    if (_T_1058) begin
      buffers_0_18_3 <= io_dataIn_bits_75;
    end
    if (_T_1058) begin
      buffers_0_19_0 <= io_dataIn_bits_76;
    end
    if (_T_1058) begin
      buffers_0_19_1 <= io_dataIn_bits_77;
    end
    if (_T_1058) begin
      buffers_0_19_2 <= io_dataIn_bits_78;
    end
    if (_T_1058) begin
      buffers_0_19_3 <= io_dataIn_bits_79;
    end
    if (_T_1058) begin
      buffers_0_20_0 <= io_dataIn_bits_80;
    end
    if (_T_1058) begin
      buffers_0_20_1 <= io_dataIn_bits_81;
    end
    if (_T_1058) begin
      buffers_0_20_2 <= io_dataIn_bits_82;
    end
    if (_T_1058) begin
      buffers_0_20_3 <= io_dataIn_bits_83;
    end
    if (_T_1058) begin
      buffers_0_21_0 <= io_dataIn_bits_84;
    end
    if (_T_1058) begin
      buffers_0_21_1 <= io_dataIn_bits_85;
    end
    if (_T_1058) begin
      buffers_0_21_2 <= io_dataIn_bits_86;
    end
    if (_T_1058) begin
      buffers_0_21_3 <= io_dataIn_bits_87;
    end
    if (_T_1058) begin
      buffers_0_22_0 <= io_dataIn_bits_88;
    end
    if (_T_1058) begin
      buffers_0_22_1 <= io_dataIn_bits_89;
    end
    if (_T_1058) begin
      buffers_0_22_2 <= io_dataIn_bits_90;
    end
    if (_T_1058) begin
      buffers_0_22_3 <= io_dataIn_bits_91;
    end
    if (_T_1058) begin
      buffers_0_23_0 <= io_dataIn_bits_92;
    end
    if (_T_1058) begin
      buffers_0_23_1 <= io_dataIn_bits_93;
    end
    if (_T_1058) begin
      buffers_0_23_2 <= io_dataIn_bits_94;
    end
    if (_T_1058) begin
      buffers_0_23_3 <= io_dataIn_bits_95;
    end
    if (_T_1058) begin
      buffers_0_24_0 <= io_dataIn_bits_96;
    end
    if (_T_1058) begin
      buffers_0_24_1 <= io_dataIn_bits_97;
    end
    if (_T_1058) begin
      buffers_0_24_2 <= io_dataIn_bits_98;
    end
    if (_T_1058) begin
      buffers_0_24_3 <= io_dataIn_bits_99;
    end
    if (_T_1058) begin
      buffers_0_25_0 <= io_dataIn_bits_100;
    end
    if (_T_1058) begin
      buffers_0_25_1 <= io_dataIn_bits_101;
    end
    if (_T_1058) begin
      buffers_0_25_2 <= io_dataIn_bits_102;
    end
    if (_T_1058) begin
      buffers_0_25_3 <= io_dataIn_bits_103;
    end
    if (_T_1058) begin
      buffers_0_26_0 <= io_dataIn_bits_104;
    end
    if (_T_1058) begin
      buffers_0_26_1 <= io_dataIn_bits_105;
    end
    if (_T_1058) begin
      buffers_0_26_2 <= io_dataIn_bits_106;
    end
    if (_T_1058) begin
      buffers_0_26_3 <= io_dataIn_bits_107;
    end
    if (_T_1058) begin
      buffers_0_27_0 <= io_dataIn_bits_108;
    end
    if (_T_1058) begin
      buffers_0_27_1 <= io_dataIn_bits_109;
    end
    if (_T_1058) begin
      buffers_0_27_2 <= io_dataIn_bits_110;
    end
    if (_T_1058) begin
      buffers_0_27_3 <= io_dataIn_bits_111;
    end
    if (_T_1058) begin
      buffers_0_28_0 <= io_dataIn_bits_112;
    end
    if (_T_1058) begin
      buffers_0_28_1 <= io_dataIn_bits_113;
    end
    if (_T_1058) begin
      buffers_0_28_2 <= io_dataIn_bits_114;
    end
    if (_T_1058) begin
      buffers_0_28_3 <= io_dataIn_bits_115;
    end
    if (_T_1058) begin
      buffers_0_29_0 <= io_dataIn_bits_116;
    end
    if (_T_1058) begin
      buffers_0_29_1 <= io_dataIn_bits_117;
    end
    if (_T_1058) begin
      buffers_0_29_2 <= io_dataIn_bits_118;
    end
    if (_T_1058) begin
      buffers_0_29_3 <= io_dataIn_bits_119;
    end
    if (_T_1058) begin
      buffers_0_30_0 <= io_dataIn_bits_120;
    end
    if (_T_1058) begin
      buffers_0_30_1 <= io_dataIn_bits_121;
    end
    if (_T_1058) begin
      buffers_0_30_2 <= io_dataIn_bits_122;
    end
    if (_T_1058) begin
      buffers_0_30_3 <= io_dataIn_bits_123;
    end
    if (_T_1058) begin
      buffers_0_31_0 <= io_dataIn_bits_124;
    end
    if (_T_1058) begin
      buffers_0_31_1 <= io_dataIn_bits_125;
    end
    if (_T_1058) begin
      buffers_0_31_2 <= io_dataIn_bits_126;
    end
    if (_T_1058) begin
      buffers_0_31_3 <= io_dataIn_bits_127;
    end
    if (_T_1058) begin
      buffers_0_32_0 <= io_dataIn_bits_128;
    end
    if (_T_1058) begin
      buffers_0_32_1 <= io_dataIn_bits_129;
    end
    if (_T_1058) begin
      buffers_0_32_2 <= io_dataIn_bits_130;
    end
    if (_T_1058) begin
      buffers_0_32_3 <= io_dataIn_bits_131;
    end
    if (_T_1058) begin
      buffers_0_33_0 <= io_dataIn_bits_132;
    end
    if (_T_1058) begin
      buffers_0_33_1 <= io_dataIn_bits_133;
    end
    if (_T_1058) begin
      buffers_0_33_2 <= io_dataIn_bits_134;
    end
    if (_T_1058) begin
      buffers_0_33_3 <= io_dataIn_bits_135;
    end
    if (_T_1058) begin
      buffers_0_34_0 <= io_dataIn_bits_136;
    end
    if (_T_1058) begin
      buffers_0_34_1 <= io_dataIn_bits_137;
    end
    if (_T_1058) begin
      buffers_0_34_2 <= io_dataIn_bits_138;
    end
    if (_T_1058) begin
      buffers_0_34_3 <= io_dataIn_bits_139;
    end
    if (_T_1058) begin
      buffers_0_35_0 <= io_dataIn_bits_140;
    end
    if (_T_1058) begin
      buffers_0_35_1 <= io_dataIn_bits_141;
    end
    if (_T_1058) begin
      buffers_0_35_2 <= io_dataIn_bits_142;
    end
    if (_T_1058) begin
      buffers_0_35_3 <= io_dataIn_bits_143;
    end
    if (_T_1058) begin
      buffers_0_36_0 <= io_dataIn_bits_144;
    end
    if (_T_1058) begin
      buffers_0_36_1 <= io_dataIn_bits_145;
    end
    if (_T_1058) begin
      buffers_0_36_2 <= io_dataIn_bits_146;
    end
    if (_T_1058) begin
      buffers_0_36_3 <= io_dataIn_bits_147;
    end
    if (_T_1058) begin
      buffers_0_37_0 <= io_dataIn_bits_148;
    end
    if (_T_1058) begin
      buffers_0_37_1 <= io_dataIn_bits_149;
    end
    if (_T_1058) begin
      buffers_0_37_2 <= io_dataIn_bits_150;
    end
    if (_T_1058) begin
      buffers_0_37_3 <= io_dataIn_bits_151;
    end
    if (_T_1058) begin
      buffers_0_38_0 <= io_dataIn_bits_152;
    end
    if (_T_1058) begin
      buffers_0_38_1 <= io_dataIn_bits_153;
    end
    if (_T_1058) begin
      buffers_0_38_2 <= io_dataIn_bits_154;
    end
    if (_T_1058) begin
      buffers_0_38_3 <= io_dataIn_bits_155;
    end
    if (_T_1058) begin
      buffers_0_39_0 <= io_dataIn_bits_156;
    end
    if (_T_1058) begin
      buffers_0_39_1 <= io_dataIn_bits_157;
    end
    if (_T_1058) begin
      buffers_0_39_2 <= io_dataIn_bits_158;
    end
    if (_T_1058) begin
      buffers_0_39_3 <= io_dataIn_bits_159;
    end
    if (_T_1058) begin
      buffers_0_40_0 <= io_dataIn_bits_160;
    end
    if (_T_1058) begin
      buffers_0_40_1 <= io_dataIn_bits_161;
    end
    if (_T_1058) begin
      buffers_0_40_2 <= io_dataIn_bits_162;
    end
    if (_T_1058) begin
      buffers_0_40_3 <= io_dataIn_bits_163;
    end
    if (_T_1058) begin
      buffers_0_41_0 <= io_dataIn_bits_164;
    end
    if (_T_1058) begin
      buffers_0_41_1 <= io_dataIn_bits_165;
    end
    if (_T_1058) begin
      buffers_0_41_2 <= io_dataIn_bits_166;
    end
    if (_T_1058) begin
      buffers_0_41_3 <= io_dataIn_bits_167;
    end
    if (_T_1058) begin
      buffers_0_42_0 <= io_dataIn_bits_168;
    end
    if (_T_1058) begin
      buffers_0_42_1 <= io_dataIn_bits_169;
    end
    if (_T_1058) begin
      buffers_0_42_2 <= io_dataIn_bits_170;
    end
    if (_T_1058) begin
      buffers_0_42_3 <= io_dataIn_bits_171;
    end
    if (_T_1058) begin
      buffers_0_43_0 <= io_dataIn_bits_172;
    end
    if (_T_1058) begin
      buffers_0_43_1 <= io_dataIn_bits_173;
    end
    if (_T_1058) begin
      buffers_0_43_2 <= io_dataIn_bits_174;
    end
    if (_T_1058) begin
      buffers_0_43_3 <= io_dataIn_bits_175;
    end
    if (_T_1058) begin
      buffers_0_44_0 <= io_dataIn_bits_176;
    end
    if (_T_1058) begin
      buffers_0_44_1 <= io_dataIn_bits_177;
    end
    if (_T_1058) begin
      buffers_0_44_2 <= io_dataIn_bits_178;
    end
    if (_T_1058) begin
      buffers_0_44_3 <= io_dataIn_bits_179;
    end
    if (_T_1058) begin
      buffers_0_45_0 <= io_dataIn_bits_180;
    end
    if (_T_1058) begin
      buffers_0_45_1 <= io_dataIn_bits_181;
    end
    if (_T_1058) begin
      buffers_0_45_2 <= io_dataIn_bits_182;
    end
    if (_T_1058) begin
      buffers_0_45_3 <= io_dataIn_bits_183;
    end
    if (_T_1058) begin
      buffers_0_46_0 <= io_dataIn_bits_184;
    end
    if (_T_1058) begin
      buffers_0_46_1 <= io_dataIn_bits_185;
    end
    if (_T_1058) begin
      buffers_0_46_2 <= io_dataIn_bits_186;
    end
    if (_T_1058) begin
      buffers_0_46_3 <= io_dataIn_bits_187;
    end
    if (_T_1058) begin
      buffers_0_47_0 <= io_dataIn_bits_188;
    end
    if (_T_1058) begin
      buffers_0_47_1 <= io_dataIn_bits_189;
    end
    if (_T_1058) begin
      buffers_0_47_2 <= io_dataIn_bits_190;
    end
    if (_T_1058) begin
      buffers_0_47_3 <= io_dataIn_bits_191;
    end
    if (_T_1058) begin
      buffers_0_48_0 <= io_dataIn_bits_192;
    end
    if (_T_1058) begin
      buffers_0_48_1 <= io_dataIn_bits_193;
    end
    if (_T_1058) begin
      buffers_0_48_2 <= io_dataIn_bits_194;
    end
    if (_T_1058) begin
      buffers_0_48_3 <= io_dataIn_bits_195;
    end
    if (_T_1058) begin
      buffers_0_49_0 <= io_dataIn_bits_196;
    end
    if (_T_1058) begin
      buffers_0_49_1 <= io_dataIn_bits_197;
    end
    if (_T_1058) begin
      buffers_0_49_2 <= io_dataIn_bits_198;
    end
    if (_T_1058) begin
      buffers_0_49_3 <= io_dataIn_bits_199;
    end
    if (_T_1058) begin
      buffers_0_50_0 <= io_dataIn_bits_200;
    end
    if (_T_1058) begin
      buffers_0_50_1 <= io_dataIn_bits_201;
    end
    if (_T_1058) begin
      buffers_0_50_2 <= io_dataIn_bits_202;
    end
    if (_T_1058) begin
      buffers_0_50_3 <= io_dataIn_bits_203;
    end
    if (_T_1058) begin
      buffers_0_51_0 <= io_dataIn_bits_204;
    end
    if (_T_1058) begin
      buffers_0_51_1 <= io_dataIn_bits_205;
    end
    if (_T_1058) begin
      buffers_0_51_2 <= io_dataIn_bits_206;
    end
    if (_T_1058) begin
      buffers_0_51_3 <= io_dataIn_bits_207;
    end
    if (_T_1058) begin
      buffers_0_52_0 <= io_dataIn_bits_208;
    end
    if (_T_1058) begin
      buffers_0_52_1 <= io_dataIn_bits_209;
    end
    if (_T_1058) begin
      buffers_0_52_2 <= io_dataIn_bits_210;
    end
    if (_T_1058) begin
      buffers_0_52_3 <= io_dataIn_bits_211;
    end
    if (_T_1058) begin
      buffers_0_53_0 <= io_dataIn_bits_212;
    end
    if (_T_1058) begin
      buffers_0_53_1 <= io_dataIn_bits_213;
    end
    if (_T_1058) begin
      buffers_0_53_2 <= io_dataIn_bits_214;
    end
    if (_T_1058) begin
      buffers_0_53_3 <= io_dataIn_bits_215;
    end
    if (_T_1058) begin
      buffers_0_54_0 <= io_dataIn_bits_216;
    end
    if (_T_1058) begin
      buffers_0_54_1 <= io_dataIn_bits_217;
    end
    if (_T_1058) begin
      buffers_0_54_2 <= io_dataIn_bits_218;
    end
    if (_T_1058) begin
      buffers_0_54_3 <= io_dataIn_bits_219;
    end
    if (_T_1058) begin
      buffers_0_55_0 <= io_dataIn_bits_220;
    end
    if (_T_1058) begin
      buffers_0_55_1 <= io_dataIn_bits_221;
    end
    if (_T_1058) begin
      buffers_0_55_2 <= io_dataIn_bits_222;
    end
    if (_T_1058) begin
      buffers_0_55_3 <= io_dataIn_bits_223;
    end
    if (_T_1058) begin
      buffers_0_56_0 <= io_dataIn_bits_224;
    end
    if (_T_1058) begin
      buffers_0_56_1 <= io_dataIn_bits_225;
    end
    if (_T_1058) begin
      buffers_0_56_2 <= io_dataIn_bits_226;
    end
    if (_T_1058) begin
      buffers_0_56_3 <= io_dataIn_bits_227;
    end
    if (_T_1058) begin
      buffers_0_57_0 <= io_dataIn_bits_228;
    end
    if (_T_1058) begin
      buffers_0_57_1 <= io_dataIn_bits_229;
    end
    if (_T_1058) begin
      buffers_0_57_2 <= io_dataIn_bits_230;
    end
    if (_T_1058) begin
      buffers_0_57_3 <= io_dataIn_bits_231;
    end
    if (_T_1058) begin
      buffers_0_58_0 <= io_dataIn_bits_232;
    end
    if (_T_1058) begin
      buffers_0_58_1 <= io_dataIn_bits_233;
    end
    if (_T_1058) begin
      buffers_0_58_2 <= io_dataIn_bits_234;
    end
    if (_T_1058) begin
      buffers_0_58_3 <= io_dataIn_bits_235;
    end
    if (_T_1058) begin
      buffers_0_59_0 <= io_dataIn_bits_236;
    end
    if (_T_1058) begin
      buffers_0_59_1 <= io_dataIn_bits_237;
    end
    if (_T_1058) begin
      buffers_0_59_2 <= io_dataIn_bits_238;
    end
    if (_T_1058) begin
      buffers_0_59_3 <= io_dataIn_bits_239;
    end
    if (_T_1058) begin
      buffers_0_60_0 <= io_dataIn_bits_240;
    end
    if (_T_1058) begin
      buffers_0_60_1 <= io_dataIn_bits_241;
    end
    if (_T_1058) begin
      buffers_0_60_2 <= io_dataIn_bits_242;
    end
    if (_T_1058) begin
      buffers_0_60_3 <= io_dataIn_bits_243;
    end
    if (_T_1058) begin
      buffers_0_61_0 <= io_dataIn_bits_244;
    end
    if (_T_1058) begin
      buffers_0_61_1 <= io_dataIn_bits_245;
    end
    if (_T_1058) begin
      buffers_0_61_2 <= io_dataIn_bits_246;
    end
    if (_T_1058) begin
      buffers_0_61_3 <= io_dataIn_bits_247;
    end
    if (_T_1058) begin
      buffers_0_62_0 <= io_dataIn_bits_248;
    end
    if (_T_1058) begin
      buffers_0_62_1 <= io_dataIn_bits_249;
    end
    if (_T_1058) begin
      buffers_0_62_2 <= io_dataIn_bits_250;
    end
    if (_T_1058) begin
      buffers_0_62_3 <= io_dataIn_bits_251;
    end
    if (_T_1058) begin
      buffers_0_63_0 <= io_dataIn_bits_252;
    end
    if (_T_1058) begin
      buffers_0_63_1 <= io_dataIn_bits_253;
    end
    if (_T_1058) begin
      buffers_0_63_2 <= io_dataIn_bits_254;
    end
    if (_T_1058) begin
      buffers_0_63_3 <= io_dataIn_bits_255;
    end
    cntrs_0 <= _T_1065;
    _T_1071 <= _T_1068;
    cntrs_1 <= _T_1071;
    _T_1076 <= _T_1073;
    _T_1078 <= _T_1076;
    cntrs_2 <= _T_1078;
    if (_T_1094) begin
      buffers_1_0_0 <= buffers_0_3_0;
    end else begin
      if (_T_1092) begin
        buffers_1_0_0 <= buffers_0_2_0;
      end else begin
        if (_T_1090) begin
          buffers_1_0_0 <= buffers_0_1_0;
        end else begin
          buffers_1_0_0 <= buffers_0_0_0;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_0_1 <= buffers_0_3_1;
    end else begin
      if (_T_1092) begin
        buffers_1_0_1 <= buffers_0_2_1;
      end else begin
        if (_T_1090) begin
          buffers_1_0_1 <= buffers_0_1_1;
        end else begin
          buffers_1_0_1 <= buffers_0_0_1;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_0_2 <= buffers_0_3_2;
    end else begin
      if (_T_1092) begin
        buffers_1_0_2 <= buffers_0_2_2;
      end else begin
        if (_T_1090) begin
          buffers_1_0_2 <= buffers_0_1_2;
        end else begin
          buffers_1_0_2 <= buffers_0_0_2;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_0_3 <= buffers_0_3_3;
    end else begin
      if (_T_1092) begin
        buffers_1_0_3 <= buffers_0_2_3;
      end else begin
        if (_T_1090) begin
          buffers_1_0_3 <= buffers_0_1_3;
        end else begin
          buffers_1_0_3 <= buffers_0_0_3;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_1_0 <= buffers_0_7_0;
    end else begin
      if (_T_1092) begin
        buffers_1_1_0 <= buffers_0_6_0;
      end else begin
        if (_T_1090) begin
          buffers_1_1_0 <= buffers_0_5_0;
        end else begin
          buffers_1_1_0 <= buffers_0_4_0;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_1_1 <= buffers_0_7_1;
    end else begin
      if (_T_1092) begin
        buffers_1_1_1 <= buffers_0_6_1;
      end else begin
        if (_T_1090) begin
          buffers_1_1_1 <= buffers_0_5_1;
        end else begin
          buffers_1_1_1 <= buffers_0_4_1;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_1_2 <= buffers_0_7_2;
    end else begin
      if (_T_1092) begin
        buffers_1_1_2 <= buffers_0_6_2;
      end else begin
        if (_T_1090) begin
          buffers_1_1_2 <= buffers_0_5_2;
        end else begin
          buffers_1_1_2 <= buffers_0_4_2;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_1_3 <= buffers_0_7_3;
    end else begin
      if (_T_1092) begin
        buffers_1_1_3 <= buffers_0_6_3;
      end else begin
        if (_T_1090) begin
          buffers_1_1_3 <= buffers_0_5_3;
        end else begin
          buffers_1_1_3 <= buffers_0_4_3;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_2_0 <= buffers_0_11_0;
    end else begin
      if (_T_1092) begin
        buffers_1_2_0 <= buffers_0_10_0;
      end else begin
        if (_T_1090) begin
          buffers_1_2_0 <= buffers_0_9_0;
        end else begin
          buffers_1_2_0 <= buffers_0_8_0;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_2_1 <= buffers_0_11_1;
    end else begin
      if (_T_1092) begin
        buffers_1_2_1 <= buffers_0_10_1;
      end else begin
        if (_T_1090) begin
          buffers_1_2_1 <= buffers_0_9_1;
        end else begin
          buffers_1_2_1 <= buffers_0_8_1;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_2_2 <= buffers_0_11_2;
    end else begin
      if (_T_1092) begin
        buffers_1_2_2 <= buffers_0_10_2;
      end else begin
        if (_T_1090) begin
          buffers_1_2_2 <= buffers_0_9_2;
        end else begin
          buffers_1_2_2 <= buffers_0_8_2;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_2_3 <= buffers_0_11_3;
    end else begin
      if (_T_1092) begin
        buffers_1_2_3 <= buffers_0_10_3;
      end else begin
        if (_T_1090) begin
          buffers_1_2_3 <= buffers_0_9_3;
        end else begin
          buffers_1_2_3 <= buffers_0_8_3;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_3_0 <= buffers_0_15_0;
    end else begin
      if (_T_1092) begin
        buffers_1_3_0 <= buffers_0_14_0;
      end else begin
        if (_T_1090) begin
          buffers_1_3_0 <= buffers_0_13_0;
        end else begin
          buffers_1_3_0 <= buffers_0_12_0;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_3_1 <= buffers_0_15_1;
    end else begin
      if (_T_1092) begin
        buffers_1_3_1 <= buffers_0_14_1;
      end else begin
        if (_T_1090) begin
          buffers_1_3_1 <= buffers_0_13_1;
        end else begin
          buffers_1_3_1 <= buffers_0_12_1;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_3_2 <= buffers_0_15_2;
    end else begin
      if (_T_1092) begin
        buffers_1_3_2 <= buffers_0_14_2;
      end else begin
        if (_T_1090) begin
          buffers_1_3_2 <= buffers_0_13_2;
        end else begin
          buffers_1_3_2 <= buffers_0_12_2;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_3_3 <= buffers_0_15_3;
    end else begin
      if (_T_1092) begin
        buffers_1_3_3 <= buffers_0_14_3;
      end else begin
        if (_T_1090) begin
          buffers_1_3_3 <= buffers_0_13_3;
        end else begin
          buffers_1_3_3 <= buffers_0_12_3;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_4_0 <= buffers_0_19_0;
    end else begin
      if (_T_1092) begin
        buffers_1_4_0 <= buffers_0_18_0;
      end else begin
        if (_T_1090) begin
          buffers_1_4_0 <= buffers_0_17_0;
        end else begin
          buffers_1_4_0 <= buffers_0_16_0;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_4_1 <= buffers_0_19_1;
    end else begin
      if (_T_1092) begin
        buffers_1_4_1 <= buffers_0_18_1;
      end else begin
        if (_T_1090) begin
          buffers_1_4_1 <= buffers_0_17_1;
        end else begin
          buffers_1_4_1 <= buffers_0_16_1;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_4_2 <= buffers_0_19_2;
    end else begin
      if (_T_1092) begin
        buffers_1_4_2 <= buffers_0_18_2;
      end else begin
        if (_T_1090) begin
          buffers_1_4_2 <= buffers_0_17_2;
        end else begin
          buffers_1_4_2 <= buffers_0_16_2;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_4_3 <= buffers_0_19_3;
    end else begin
      if (_T_1092) begin
        buffers_1_4_3 <= buffers_0_18_3;
      end else begin
        if (_T_1090) begin
          buffers_1_4_3 <= buffers_0_17_3;
        end else begin
          buffers_1_4_3 <= buffers_0_16_3;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_5_0 <= buffers_0_23_0;
    end else begin
      if (_T_1092) begin
        buffers_1_5_0 <= buffers_0_22_0;
      end else begin
        if (_T_1090) begin
          buffers_1_5_0 <= buffers_0_21_0;
        end else begin
          buffers_1_5_0 <= buffers_0_20_0;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_5_1 <= buffers_0_23_1;
    end else begin
      if (_T_1092) begin
        buffers_1_5_1 <= buffers_0_22_1;
      end else begin
        if (_T_1090) begin
          buffers_1_5_1 <= buffers_0_21_1;
        end else begin
          buffers_1_5_1 <= buffers_0_20_1;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_5_2 <= buffers_0_23_2;
    end else begin
      if (_T_1092) begin
        buffers_1_5_2 <= buffers_0_22_2;
      end else begin
        if (_T_1090) begin
          buffers_1_5_2 <= buffers_0_21_2;
        end else begin
          buffers_1_5_2 <= buffers_0_20_2;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_5_3 <= buffers_0_23_3;
    end else begin
      if (_T_1092) begin
        buffers_1_5_3 <= buffers_0_22_3;
      end else begin
        if (_T_1090) begin
          buffers_1_5_3 <= buffers_0_21_3;
        end else begin
          buffers_1_5_3 <= buffers_0_20_3;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_6_0 <= buffers_0_27_0;
    end else begin
      if (_T_1092) begin
        buffers_1_6_0 <= buffers_0_26_0;
      end else begin
        if (_T_1090) begin
          buffers_1_6_0 <= buffers_0_25_0;
        end else begin
          buffers_1_6_0 <= buffers_0_24_0;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_6_1 <= buffers_0_27_1;
    end else begin
      if (_T_1092) begin
        buffers_1_6_1 <= buffers_0_26_1;
      end else begin
        if (_T_1090) begin
          buffers_1_6_1 <= buffers_0_25_1;
        end else begin
          buffers_1_6_1 <= buffers_0_24_1;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_6_2 <= buffers_0_27_2;
    end else begin
      if (_T_1092) begin
        buffers_1_6_2 <= buffers_0_26_2;
      end else begin
        if (_T_1090) begin
          buffers_1_6_2 <= buffers_0_25_2;
        end else begin
          buffers_1_6_2 <= buffers_0_24_2;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_6_3 <= buffers_0_27_3;
    end else begin
      if (_T_1092) begin
        buffers_1_6_3 <= buffers_0_26_3;
      end else begin
        if (_T_1090) begin
          buffers_1_6_3 <= buffers_0_25_3;
        end else begin
          buffers_1_6_3 <= buffers_0_24_3;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_7_0 <= buffers_0_31_0;
    end else begin
      if (_T_1092) begin
        buffers_1_7_0 <= buffers_0_30_0;
      end else begin
        if (_T_1090) begin
          buffers_1_7_0 <= buffers_0_29_0;
        end else begin
          buffers_1_7_0 <= buffers_0_28_0;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_7_1 <= buffers_0_31_1;
    end else begin
      if (_T_1092) begin
        buffers_1_7_1 <= buffers_0_30_1;
      end else begin
        if (_T_1090) begin
          buffers_1_7_1 <= buffers_0_29_1;
        end else begin
          buffers_1_7_1 <= buffers_0_28_1;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_7_2 <= buffers_0_31_2;
    end else begin
      if (_T_1092) begin
        buffers_1_7_2 <= buffers_0_30_2;
      end else begin
        if (_T_1090) begin
          buffers_1_7_2 <= buffers_0_29_2;
        end else begin
          buffers_1_7_2 <= buffers_0_28_2;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_7_3 <= buffers_0_31_3;
    end else begin
      if (_T_1092) begin
        buffers_1_7_3 <= buffers_0_30_3;
      end else begin
        if (_T_1090) begin
          buffers_1_7_3 <= buffers_0_29_3;
        end else begin
          buffers_1_7_3 <= buffers_0_28_3;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_8_0 <= buffers_0_35_0;
    end else begin
      if (_T_1092) begin
        buffers_1_8_0 <= buffers_0_34_0;
      end else begin
        if (_T_1090) begin
          buffers_1_8_0 <= buffers_0_33_0;
        end else begin
          buffers_1_8_0 <= buffers_0_32_0;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_8_1 <= buffers_0_35_1;
    end else begin
      if (_T_1092) begin
        buffers_1_8_1 <= buffers_0_34_1;
      end else begin
        if (_T_1090) begin
          buffers_1_8_1 <= buffers_0_33_1;
        end else begin
          buffers_1_8_1 <= buffers_0_32_1;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_8_2 <= buffers_0_35_2;
    end else begin
      if (_T_1092) begin
        buffers_1_8_2 <= buffers_0_34_2;
      end else begin
        if (_T_1090) begin
          buffers_1_8_2 <= buffers_0_33_2;
        end else begin
          buffers_1_8_2 <= buffers_0_32_2;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_8_3 <= buffers_0_35_3;
    end else begin
      if (_T_1092) begin
        buffers_1_8_3 <= buffers_0_34_3;
      end else begin
        if (_T_1090) begin
          buffers_1_8_3 <= buffers_0_33_3;
        end else begin
          buffers_1_8_3 <= buffers_0_32_3;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_9_0 <= buffers_0_39_0;
    end else begin
      if (_T_1092) begin
        buffers_1_9_0 <= buffers_0_38_0;
      end else begin
        if (_T_1090) begin
          buffers_1_9_0 <= buffers_0_37_0;
        end else begin
          buffers_1_9_0 <= buffers_0_36_0;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_9_1 <= buffers_0_39_1;
    end else begin
      if (_T_1092) begin
        buffers_1_9_1 <= buffers_0_38_1;
      end else begin
        if (_T_1090) begin
          buffers_1_9_1 <= buffers_0_37_1;
        end else begin
          buffers_1_9_1 <= buffers_0_36_1;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_9_2 <= buffers_0_39_2;
    end else begin
      if (_T_1092) begin
        buffers_1_9_2 <= buffers_0_38_2;
      end else begin
        if (_T_1090) begin
          buffers_1_9_2 <= buffers_0_37_2;
        end else begin
          buffers_1_9_2 <= buffers_0_36_2;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_9_3 <= buffers_0_39_3;
    end else begin
      if (_T_1092) begin
        buffers_1_9_3 <= buffers_0_38_3;
      end else begin
        if (_T_1090) begin
          buffers_1_9_3 <= buffers_0_37_3;
        end else begin
          buffers_1_9_3 <= buffers_0_36_3;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_10_0 <= buffers_0_43_0;
    end else begin
      if (_T_1092) begin
        buffers_1_10_0 <= buffers_0_42_0;
      end else begin
        if (_T_1090) begin
          buffers_1_10_0 <= buffers_0_41_0;
        end else begin
          buffers_1_10_0 <= buffers_0_40_0;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_10_1 <= buffers_0_43_1;
    end else begin
      if (_T_1092) begin
        buffers_1_10_1 <= buffers_0_42_1;
      end else begin
        if (_T_1090) begin
          buffers_1_10_1 <= buffers_0_41_1;
        end else begin
          buffers_1_10_1 <= buffers_0_40_1;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_10_2 <= buffers_0_43_2;
    end else begin
      if (_T_1092) begin
        buffers_1_10_2 <= buffers_0_42_2;
      end else begin
        if (_T_1090) begin
          buffers_1_10_2 <= buffers_0_41_2;
        end else begin
          buffers_1_10_2 <= buffers_0_40_2;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_10_3 <= buffers_0_43_3;
    end else begin
      if (_T_1092) begin
        buffers_1_10_3 <= buffers_0_42_3;
      end else begin
        if (_T_1090) begin
          buffers_1_10_3 <= buffers_0_41_3;
        end else begin
          buffers_1_10_3 <= buffers_0_40_3;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_11_0 <= buffers_0_47_0;
    end else begin
      if (_T_1092) begin
        buffers_1_11_0 <= buffers_0_46_0;
      end else begin
        if (_T_1090) begin
          buffers_1_11_0 <= buffers_0_45_0;
        end else begin
          buffers_1_11_0 <= buffers_0_44_0;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_11_1 <= buffers_0_47_1;
    end else begin
      if (_T_1092) begin
        buffers_1_11_1 <= buffers_0_46_1;
      end else begin
        if (_T_1090) begin
          buffers_1_11_1 <= buffers_0_45_1;
        end else begin
          buffers_1_11_1 <= buffers_0_44_1;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_11_2 <= buffers_0_47_2;
    end else begin
      if (_T_1092) begin
        buffers_1_11_2 <= buffers_0_46_2;
      end else begin
        if (_T_1090) begin
          buffers_1_11_2 <= buffers_0_45_2;
        end else begin
          buffers_1_11_2 <= buffers_0_44_2;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_11_3 <= buffers_0_47_3;
    end else begin
      if (_T_1092) begin
        buffers_1_11_3 <= buffers_0_46_3;
      end else begin
        if (_T_1090) begin
          buffers_1_11_3 <= buffers_0_45_3;
        end else begin
          buffers_1_11_3 <= buffers_0_44_3;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_12_0 <= buffers_0_51_0;
    end else begin
      if (_T_1092) begin
        buffers_1_12_0 <= buffers_0_50_0;
      end else begin
        if (_T_1090) begin
          buffers_1_12_0 <= buffers_0_49_0;
        end else begin
          buffers_1_12_0 <= buffers_0_48_0;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_12_1 <= buffers_0_51_1;
    end else begin
      if (_T_1092) begin
        buffers_1_12_1 <= buffers_0_50_1;
      end else begin
        if (_T_1090) begin
          buffers_1_12_1 <= buffers_0_49_1;
        end else begin
          buffers_1_12_1 <= buffers_0_48_1;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_12_2 <= buffers_0_51_2;
    end else begin
      if (_T_1092) begin
        buffers_1_12_2 <= buffers_0_50_2;
      end else begin
        if (_T_1090) begin
          buffers_1_12_2 <= buffers_0_49_2;
        end else begin
          buffers_1_12_2 <= buffers_0_48_2;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_12_3 <= buffers_0_51_3;
    end else begin
      if (_T_1092) begin
        buffers_1_12_3 <= buffers_0_50_3;
      end else begin
        if (_T_1090) begin
          buffers_1_12_3 <= buffers_0_49_3;
        end else begin
          buffers_1_12_3 <= buffers_0_48_3;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_13_0 <= buffers_0_55_0;
    end else begin
      if (_T_1092) begin
        buffers_1_13_0 <= buffers_0_54_0;
      end else begin
        if (_T_1090) begin
          buffers_1_13_0 <= buffers_0_53_0;
        end else begin
          buffers_1_13_0 <= buffers_0_52_0;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_13_1 <= buffers_0_55_1;
    end else begin
      if (_T_1092) begin
        buffers_1_13_1 <= buffers_0_54_1;
      end else begin
        if (_T_1090) begin
          buffers_1_13_1 <= buffers_0_53_1;
        end else begin
          buffers_1_13_1 <= buffers_0_52_1;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_13_2 <= buffers_0_55_2;
    end else begin
      if (_T_1092) begin
        buffers_1_13_2 <= buffers_0_54_2;
      end else begin
        if (_T_1090) begin
          buffers_1_13_2 <= buffers_0_53_2;
        end else begin
          buffers_1_13_2 <= buffers_0_52_2;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_13_3 <= buffers_0_55_3;
    end else begin
      if (_T_1092) begin
        buffers_1_13_3 <= buffers_0_54_3;
      end else begin
        if (_T_1090) begin
          buffers_1_13_3 <= buffers_0_53_3;
        end else begin
          buffers_1_13_3 <= buffers_0_52_3;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_14_0 <= buffers_0_59_0;
    end else begin
      if (_T_1092) begin
        buffers_1_14_0 <= buffers_0_58_0;
      end else begin
        if (_T_1090) begin
          buffers_1_14_0 <= buffers_0_57_0;
        end else begin
          buffers_1_14_0 <= buffers_0_56_0;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_14_1 <= buffers_0_59_1;
    end else begin
      if (_T_1092) begin
        buffers_1_14_1 <= buffers_0_58_1;
      end else begin
        if (_T_1090) begin
          buffers_1_14_1 <= buffers_0_57_1;
        end else begin
          buffers_1_14_1 <= buffers_0_56_1;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_14_2 <= buffers_0_59_2;
    end else begin
      if (_T_1092) begin
        buffers_1_14_2 <= buffers_0_58_2;
      end else begin
        if (_T_1090) begin
          buffers_1_14_2 <= buffers_0_57_2;
        end else begin
          buffers_1_14_2 <= buffers_0_56_2;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_14_3 <= buffers_0_59_3;
    end else begin
      if (_T_1092) begin
        buffers_1_14_3 <= buffers_0_58_3;
      end else begin
        if (_T_1090) begin
          buffers_1_14_3 <= buffers_0_57_3;
        end else begin
          buffers_1_14_3 <= buffers_0_56_3;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_15_0 <= buffers_0_63_0;
    end else begin
      if (_T_1092) begin
        buffers_1_15_0 <= buffers_0_62_0;
      end else begin
        if (_T_1090) begin
          buffers_1_15_0 <= buffers_0_61_0;
        end else begin
          buffers_1_15_0 <= buffers_0_60_0;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_15_1 <= buffers_0_63_1;
    end else begin
      if (_T_1092) begin
        buffers_1_15_1 <= buffers_0_62_1;
      end else begin
        if (_T_1090) begin
          buffers_1_15_1 <= buffers_0_61_1;
        end else begin
          buffers_1_15_1 <= buffers_0_60_1;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_15_2 <= buffers_0_63_2;
    end else begin
      if (_T_1092) begin
        buffers_1_15_2 <= buffers_0_62_2;
      end else begin
        if (_T_1090) begin
          buffers_1_15_2 <= buffers_0_61_2;
        end else begin
          buffers_1_15_2 <= buffers_0_60_2;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_15_3 <= buffers_0_63_3;
    end else begin
      if (_T_1092) begin
        buffers_1_15_3 <= buffers_0_62_3;
      end else begin
        if (_T_1090) begin
          buffers_1_15_3 <= buffers_0_61_3;
        end else begin
          buffers_1_15_3 <= buffers_0_60_3;
        end
      end
    end
    if (_T_1782) begin
      buffers_2_0_0 <= buffers_1_3_0;
    end else begin
      if (_T_1780) begin
        buffers_2_0_0 <= buffers_1_2_0;
      end else begin
        if (_T_1778) begin
          buffers_2_0_0 <= buffers_1_1_0;
        end else begin
          buffers_2_0_0 <= buffers_1_0_0;
        end
      end
    end
    if (_T_1782) begin
      buffers_2_0_1 <= buffers_1_3_1;
    end else begin
      if (_T_1780) begin
        buffers_2_0_1 <= buffers_1_2_1;
      end else begin
        if (_T_1778) begin
          buffers_2_0_1 <= buffers_1_1_1;
        end else begin
          buffers_2_0_1 <= buffers_1_0_1;
        end
      end
    end
    if (_T_1782) begin
      buffers_2_0_2 <= buffers_1_3_2;
    end else begin
      if (_T_1780) begin
        buffers_2_0_2 <= buffers_1_2_2;
      end else begin
        if (_T_1778) begin
          buffers_2_0_2 <= buffers_1_1_2;
        end else begin
          buffers_2_0_2 <= buffers_1_0_2;
        end
      end
    end
    if (_T_1782) begin
      buffers_2_0_3 <= buffers_1_3_3;
    end else begin
      if (_T_1780) begin
        buffers_2_0_3 <= buffers_1_2_3;
      end else begin
        if (_T_1778) begin
          buffers_2_0_3 <= buffers_1_1_3;
        end else begin
          buffers_2_0_3 <= buffers_1_0_3;
        end
      end
    end
    if (_T_1782) begin
      buffers_2_1_0 <= buffers_1_7_0;
    end else begin
      if (_T_1780) begin
        buffers_2_1_0 <= buffers_1_6_0;
      end else begin
        if (_T_1778) begin
          buffers_2_1_0 <= buffers_1_5_0;
        end else begin
          buffers_2_1_0 <= buffers_1_4_0;
        end
      end
    end
    if (_T_1782) begin
      buffers_2_1_1 <= buffers_1_7_1;
    end else begin
      if (_T_1780) begin
        buffers_2_1_1 <= buffers_1_6_1;
      end else begin
        if (_T_1778) begin
          buffers_2_1_1 <= buffers_1_5_1;
        end else begin
          buffers_2_1_1 <= buffers_1_4_1;
        end
      end
    end
    if (_T_1782) begin
      buffers_2_1_2 <= buffers_1_7_2;
    end else begin
      if (_T_1780) begin
        buffers_2_1_2 <= buffers_1_6_2;
      end else begin
        if (_T_1778) begin
          buffers_2_1_2 <= buffers_1_5_2;
        end else begin
          buffers_2_1_2 <= buffers_1_4_2;
        end
      end
    end
    if (_T_1782) begin
      buffers_2_1_3 <= buffers_1_7_3;
    end else begin
      if (_T_1780) begin
        buffers_2_1_3 <= buffers_1_6_3;
      end else begin
        if (_T_1778) begin
          buffers_2_1_3 <= buffers_1_5_3;
        end else begin
          buffers_2_1_3 <= buffers_1_4_3;
        end
      end
    end
    if (_T_1782) begin
      buffers_2_2_0 <= buffers_1_11_0;
    end else begin
      if (_T_1780) begin
        buffers_2_2_0 <= buffers_1_10_0;
      end else begin
        if (_T_1778) begin
          buffers_2_2_0 <= buffers_1_9_0;
        end else begin
          buffers_2_2_0 <= buffers_1_8_0;
        end
      end
    end
    if (_T_1782) begin
      buffers_2_2_1 <= buffers_1_11_1;
    end else begin
      if (_T_1780) begin
        buffers_2_2_1 <= buffers_1_10_1;
      end else begin
        if (_T_1778) begin
          buffers_2_2_1 <= buffers_1_9_1;
        end else begin
          buffers_2_2_1 <= buffers_1_8_1;
        end
      end
    end
    if (_T_1782) begin
      buffers_2_2_2 <= buffers_1_11_2;
    end else begin
      if (_T_1780) begin
        buffers_2_2_2 <= buffers_1_10_2;
      end else begin
        if (_T_1778) begin
          buffers_2_2_2 <= buffers_1_9_2;
        end else begin
          buffers_2_2_2 <= buffers_1_8_2;
        end
      end
    end
    if (_T_1782) begin
      buffers_2_2_3 <= buffers_1_11_3;
    end else begin
      if (_T_1780) begin
        buffers_2_2_3 <= buffers_1_10_3;
      end else begin
        if (_T_1778) begin
          buffers_2_2_3 <= buffers_1_9_3;
        end else begin
          buffers_2_2_3 <= buffers_1_8_3;
        end
      end
    end
    if (_T_1782) begin
      buffers_2_3_0 <= buffers_1_15_0;
    end else begin
      if (_T_1780) begin
        buffers_2_3_0 <= buffers_1_14_0;
      end else begin
        if (_T_1778) begin
          buffers_2_3_0 <= buffers_1_13_0;
        end else begin
          buffers_2_3_0 <= buffers_1_12_0;
        end
      end
    end
    if (_T_1782) begin
      buffers_2_3_1 <= buffers_1_15_1;
    end else begin
      if (_T_1780) begin
        buffers_2_3_1 <= buffers_1_14_1;
      end else begin
        if (_T_1778) begin
          buffers_2_3_1 <= buffers_1_13_1;
        end else begin
          buffers_2_3_1 <= buffers_1_12_1;
        end
      end
    end
    if (_T_1782) begin
      buffers_2_3_2 <= buffers_1_15_2;
    end else begin
      if (_T_1780) begin
        buffers_2_3_2 <= buffers_1_14_2;
      end else begin
        if (_T_1778) begin
          buffers_2_3_2 <= buffers_1_13_2;
        end else begin
          buffers_2_3_2 <= buffers_1_12_2;
        end
      end
    end
    if (_T_1782) begin
      buffers_2_3_3 <= buffers_1_15_3;
    end else begin
      if (_T_1780) begin
        buffers_2_3_3 <= buffers_1_14_3;
      end else begin
        if (_T_1778) begin
          buffers_2_3_3 <= buffers_1_13_3;
        end else begin
          buffers_2_3_3 <= buffers_1_12_3;
        end
      end
    end
    if (_T_1954) begin
      buffers_3_0_0 <= buffers_2_3_0;
    end else begin
      if (_T_1952) begin
        buffers_3_0_0 <= buffers_2_2_0;
      end else begin
        if (_T_1950) begin
          buffers_3_0_0 <= buffers_2_1_0;
        end else begin
          buffers_3_0_0 <= buffers_2_0_0;
        end
      end
    end
    if (_T_1954) begin
      buffers_3_0_1 <= buffers_2_3_1;
    end else begin
      if (_T_1952) begin
        buffers_3_0_1 <= buffers_2_2_1;
      end else begin
        if (_T_1950) begin
          buffers_3_0_1 <= buffers_2_1_1;
        end else begin
          buffers_3_0_1 <= buffers_2_0_1;
        end
      end
    end
    if (_T_1954) begin
      buffers_3_0_2 <= buffers_2_3_2;
    end else begin
      if (_T_1952) begin
        buffers_3_0_2 <= buffers_2_2_2;
      end else begin
        if (_T_1950) begin
          buffers_3_0_2 <= buffers_2_1_2;
        end else begin
          buffers_3_0_2 <= buffers_2_0_2;
        end
      end
    end
    if (_T_1954) begin
      buffers_3_0_3 <= buffers_2_3_3;
    end else begin
      if (_T_1952) begin
        buffers_3_0_3 <= buffers_2_2_3;
      end else begin
        if (_T_1950) begin
          buffers_3_0_3 <= buffers_2_1_3;
        end else begin
          buffers_3_0_3 <= buffers_2_0_3;
        end
      end
    end
    if (reset) begin
      _T_1988 <= 1'h0;
    end else begin
      _T_1988 <= _T_1052;
    end
    if (reset) begin
      _T_1990 <= 1'h0;
    end else begin
      _T_1990 <= _T_1988;
    end
    if (reset) begin
      vld <= 1'h0;
    end else begin
      vld <= _T_1990;
    end
    if (reset) begin
      lastVld <= 1'h0;
    end else begin
      lastVld <= vld;
    end
  end
endmodule
module AWSVggWrapper(
  input         clock,
  input         reset,
  output        io_dataIn_ready,
  input         io_dataIn_valid,
  input  [15:0] io_dataIn_bits_0,
  input  [15:0] io_dataIn_bits_1,
  input  [15:0] io_dataIn_bits_2,
  input         io_dataOut_ready,
  output        io_dataOut_valid,
  output [15:0] io_dataOut_bits_0,
  output [15:0] io_dataOut_bits_1,
  output [15:0] io_dataOut_bits_2,
  output [15:0] io_dataOut_bits_3
);
  wire  vgg_clock; // @[AWSVggWrapper.scala 46:27]
  wire  vgg_reset; // @[AWSVggWrapper.scala 46:27]
  wire  vgg_io_dataIn_ready; // @[AWSVggWrapper.scala 46:27]
  wire  vgg_io_dataIn_valid; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataIn_bits_0; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataIn_bits_1; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataIn_bits_2; // @[AWSVggWrapper.scala 46:27]
  wire  vgg_io_dataOut_ready; // @[AWSVggWrapper.scala 46:27]
  wire  vgg_io_dataOut_valid; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_0; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_1; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_2; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_3; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_4; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_5; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_6; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_7; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_8; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_9; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_10; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_11; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_12; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_13; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_14; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_15; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_16; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_17; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_18; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_19; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_20; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_21; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_22; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_23; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_24; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_25; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_26; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_27; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_28; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_29; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_30; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_31; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_32; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_33; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_34; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_35; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_36; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_37; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_38; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_39; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_40; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_41; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_42; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_43; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_44; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_45; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_46; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_47; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_48; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_49; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_50; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_51; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_52; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_53; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_54; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_55; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_56; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_57; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_58; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_59; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_60; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_61; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_62; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_63; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_64; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_65; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_66; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_67; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_68; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_69; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_70; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_71; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_72; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_73; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_74; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_75; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_76; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_77; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_78; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_79; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_80; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_81; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_82; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_83; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_84; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_85; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_86; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_87; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_88; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_89; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_90; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_91; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_92; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_93; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_94; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_95; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_96; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_97; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_98; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_99; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_100; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_101; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_102; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_103; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_104; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_105; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_106; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_107; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_108; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_109; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_110; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_111; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_112; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_113; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_114; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_115; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_116; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_117; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_118; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_119; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_120; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_121; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_122; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_123; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_124; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_125; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_126; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_127; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_128; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_129; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_130; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_131; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_132; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_133; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_134; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_135; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_136; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_137; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_138; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_139; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_140; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_141; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_142; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_143; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_144; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_145; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_146; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_147; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_148; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_149; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_150; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_151; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_152; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_153; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_154; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_155; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_156; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_157; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_158; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_159; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_160; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_161; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_162; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_163; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_164; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_165; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_166; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_167; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_168; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_169; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_170; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_171; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_172; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_173; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_174; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_175; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_176; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_177; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_178; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_179; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_180; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_181; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_182; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_183; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_184; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_185; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_186; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_187; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_188; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_189; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_190; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_191; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_192; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_193; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_194; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_195; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_196; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_197; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_198; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_199; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_200; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_201; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_202; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_203; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_204; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_205; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_206; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_207; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_208; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_209; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_210; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_211; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_212; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_213; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_214; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_215; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_216; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_217; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_218; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_219; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_220; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_221; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_222; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_223; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_224; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_225; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_226; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_227; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_228; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_229; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_230; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_231; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_232; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_233; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_234; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_235; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_236; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_237; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_238; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_239; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_240; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_241; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_242; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_243; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_244; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_245; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_246; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_247; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_248; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_249; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_250; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_251; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_252; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_253; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_254; // @[AWSVggWrapper.scala 46:27]
  wire [15:0] vgg_io_dataOut_bits_255; // @[AWSVggWrapper.scala 46:27]
  wire  queueIOOut_clock; // @[Decoupled.scala 289:19]
  wire  queueIOOut_reset; // @[Decoupled.scala 289:19]
  wire  queueIOOut_io_enq_ready; // @[Decoupled.scala 289:19]
  wire  queueIOOut_io_enq_valid; // @[Decoupled.scala 289:19]
  wire [4095:0] queueIOOut_io_enq_bits; // @[Decoupled.scala 289:19]
  wire  queueIOOut_io_deq_ready; // @[Decoupled.scala 289:19]
  wire  queueIOOut_io_deq_valid; // @[Decoupled.scala 289:19]
  wire [4095:0] queueIOOut_io_deq_bits; // @[Decoupled.scala 289:19]
  wire  muxLyr_clock; // @[AWSVggWrapper.scala 65:22]
  wire  muxLyr_reset; // @[AWSVggWrapper.scala 65:22]
  wire  muxLyr_io_dataIn_ready; // @[AWSVggWrapper.scala 65:22]
  wire  muxLyr_io_dataIn_valid; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_0; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_1; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_2; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_3; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_4; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_5; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_6; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_7; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_8; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_9; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_10; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_11; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_12; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_13; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_14; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_15; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_16; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_17; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_18; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_19; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_20; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_21; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_22; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_23; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_24; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_25; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_26; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_27; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_28; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_29; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_30; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_31; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_32; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_33; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_34; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_35; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_36; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_37; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_38; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_39; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_40; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_41; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_42; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_43; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_44; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_45; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_46; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_47; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_48; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_49; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_50; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_51; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_52; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_53; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_54; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_55; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_56; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_57; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_58; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_59; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_60; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_61; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_62; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_63; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_64; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_65; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_66; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_67; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_68; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_69; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_70; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_71; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_72; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_73; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_74; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_75; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_76; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_77; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_78; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_79; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_80; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_81; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_82; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_83; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_84; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_85; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_86; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_87; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_88; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_89; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_90; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_91; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_92; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_93; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_94; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_95; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_96; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_97; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_98; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_99; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_100; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_101; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_102; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_103; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_104; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_105; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_106; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_107; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_108; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_109; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_110; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_111; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_112; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_113; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_114; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_115; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_116; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_117; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_118; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_119; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_120; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_121; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_122; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_123; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_124; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_125; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_126; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_127; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_128; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_129; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_130; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_131; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_132; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_133; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_134; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_135; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_136; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_137; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_138; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_139; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_140; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_141; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_142; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_143; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_144; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_145; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_146; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_147; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_148; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_149; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_150; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_151; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_152; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_153; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_154; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_155; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_156; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_157; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_158; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_159; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_160; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_161; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_162; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_163; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_164; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_165; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_166; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_167; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_168; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_169; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_170; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_171; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_172; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_173; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_174; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_175; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_176; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_177; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_178; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_179; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_180; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_181; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_182; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_183; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_184; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_185; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_186; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_187; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_188; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_189; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_190; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_191; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_192; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_193; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_194; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_195; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_196; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_197; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_198; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_199; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_200; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_201; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_202; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_203; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_204; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_205; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_206; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_207; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_208; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_209; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_210; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_211; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_212; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_213; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_214; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_215; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_216; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_217; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_218; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_219; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_220; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_221; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_222; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_223; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_224; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_225; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_226; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_227; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_228; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_229; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_230; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_231; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_232; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_233; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_234; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_235; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_236; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_237; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_238; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_239; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_240; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_241; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_242; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_243; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_244; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_245; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_246; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_247; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_248; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_249; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_250; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_251; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_252; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_253; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_254; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataIn_bits_255; // @[AWSVggWrapper.scala 65:22]
  wire  muxLyr_io_dataOut_valid; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataOut_bits_0; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataOut_bits_1; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataOut_bits_2; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] muxLyr_io_dataOut_bits_3; // @[AWSVggWrapper.scala 65:22]
  wire [15:0] _T_29; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_30; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_31; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_32; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_33; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_34; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_35; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_36; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_37; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_38; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_39; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_40; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_41; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_42; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_43; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_44; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_45; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_46; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_47; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_48; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_49; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_50; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_51; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_52; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_53; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_54; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_55; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_56; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_57; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_58; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_59; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_60; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_61; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_62; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_63; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_64; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_65; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_66; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_67; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_68; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_69; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_70; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_71; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_72; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_73; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_74; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_75; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_76; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_77; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_78; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_79; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_80; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_81; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_82; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_83; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_84; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_85; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_86; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_87; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_88; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_89; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_90; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_91; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_92; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_93; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_94; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_95; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_96; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_97; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_98; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_99; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_100; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_101; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_102; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_103; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_104; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_105; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_106; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_107; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_108; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_109; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_110; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_111; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_112; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_113; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_114; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_115; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_116; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_117; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_118; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_119; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_120; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_121; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_122; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_123; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_124; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_125; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_126; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_127; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_128; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_129; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_130; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_131; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_132; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_133; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_134; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_135; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_136; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_137; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_138; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_139; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_140; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_141; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_142; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_143; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_144; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_145; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_146; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_147; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_148; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_149; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_150; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_151; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_152; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_153; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_154; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_155; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_156; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_157; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_158; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_159; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_160; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_161; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_162; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_163; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_164; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_165; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_166; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_167; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_168; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_169; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_170; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_171; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_172; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_173; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_174; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_175; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_176; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_177; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_178; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_179; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_180; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_181; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_182; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_183; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_184; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_185; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_186; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_187; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_188; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_189; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_190; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_191; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_192; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_193; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_194; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_195; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_196; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_197; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_198; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_199; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_200; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_201; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_202; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_203; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_204; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_205; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_206; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_207; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_208; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_209; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_210; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_211; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_212; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_213; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_214; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_215; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_216; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_217; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_218; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_219; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_220; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_221; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_222; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_223; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_224; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_225; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_226; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_227; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_228; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_229; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_230; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_231; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_232; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_233; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_234; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_235; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_236; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_237; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_238; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_239; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_240; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_241; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_242; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_243; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_244; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_245; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_246; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_247; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_248; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_249; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_250; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_251; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_252; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_253; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_254; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_255; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_256; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_257; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_258; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_259; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_260; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_261; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_262; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_263; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_264; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_265; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_266; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_267; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_268; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_269; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_270; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_271; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_272; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_273; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_274; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_275; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_276; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_277; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_278; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_279; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_280; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_281; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_282; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_283; // @[AWSVggWrapper.scala 52:79]
  wire [15:0] _T_284; // @[AWSVggWrapper.scala 52:79]
  wire [31:0] _T_285; // @[AWSVggWrapper.scala 52:94]
  wire [47:0] _T_286; // @[AWSVggWrapper.scala 52:94]
  wire [63:0] _T_287; // @[AWSVggWrapper.scala 52:94]
  wire [79:0] _T_288; // @[AWSVggWrapper.scala 52:94]
  wire [95:0] _T_289; // @[AWSVggWrapper.scala 52:94]
  wire [111:0] _T_290; // @[AWSVggWrapper.scala 52:94]
  wire [127:0] _T_291; // @[AWSVggWrapper.scala 52:94]
  wire [143:0] _T_292; // @[AWSVggWrapper.scala 52:94]
  wire [159:0] _T_293; // @[AWSVggWrapper.scala 52:94]
  wire [175:0] _T_294; // @[AWSVggWrapper.scala 52:94]
  wire [191:0] _T_295; // @[AWSVggWrapper.scala 52:94]
  wire [207:0] _T_296; // @[AWSVggWrapper.scala 52:94]
  wire [223:0] _T_297; // @[AWSVggWrapper.scala 52:94]
  wire [239:0] _T_298; // @[AWSVggWrapper.scala 52:94]
  wire [255:0] _T_299; // @[AWSVggWrapper.scala 52:94]
  wire [271:0] _T_300; // @[AWSVggWrapper.scala 52:94]
  wire [287:0] _T_301; // @[AWSVggWrapper.scala 52:94]
  wire [303:0] _T_302; // @[AWSVggWrapper.scala 52:94]
  wire [319:0] _T_303; // @[AWSVggWrapper.scala 52:94]
  wire [335:0] _T_304; // @[AWSVggWrapper.scala 52:94]
  wire [351:0] _T_305; // @[AWSVggWrapper.scala 52:94]
  wire [367:0] _T_306; // @[AWSVggWrapper.scala 52:94]
  wire [383:0] _T_307; // @[AWSVggWrapper.scala 52:94]
  wire [399:0] _T_308; // @[AWSVggWrapper.scala 52:94]
  wire [415:0] _T_309; // @[AWSVggWrapper.scala 52:94]
  wire [431:0] _T_310; // @[AWSVggWrapper.scala 52:94]
  wire [447:0] _T_311; // @[AWSVggWrapper.scala 52:94]
  wire [463:0] _T_312; // @[AWSVggWrapper.scala 52:94]
  wire [479:0] _T_313; // @[AWSVggWrapper.scala 52:94]
  wire [495:0] _T_314; // @[AWSVggWrapper.scala 52:94]
  wire [511:0] _T_315; // @[AWSVggWrapper.scala 52:94]
  wire [527:0] _T_316; // @[AWSVggWrapper.scala 52:94]
  wire [543:0] _T_317; // @[AWSVggWrapper.scala 52:94]
  wire [559:0] _T_318; // @[AWSVggWrapper.scala 52:94]
  wire [575:0] _T_319; // @[AWSVggWrapper.scala 52:94]
  wire [591:0] _T_320; // @[AWSVggWrapper.scala 52:94]
  wire [607:0] _T_321; // @[AWSVggWrapper.scala 52:94]
  wire [623:0] _T_322; // @[AWSVggWrapper.scala 52:94]
  wire [639:0] _T_323; // @[AWSVggWrapper.scala 52:94]
  wire [655:0] _T_324; // @[AWSVggWrapper.scala 52:94]
  wire [671:0] _T_325; // @[AWSVggWrapper.scala 52:94]
  wire [687:0] _T_326; // @[AWSVggWrapper.scala 52:94]
  wire [703:0] _T_327; // @[AWSVggWrapper.scala 52:94]
  wire [719:0] _T_328; // @[AWSVggWrapper.scala 52:94]
  wire [735:0] _T_329; // @[AWSVggWrapper.scala 52:94]
  wire [751:0] _T_330; // @[AWSVggWrapper.scala 52:94]
  wire [767:0] _T_331; // @[AWSVggWrapper.scala 52:94]
  wire [783:0] _T_332; // @[AWSVggWrapper.scala 52:94]
  wire [799:0] _T_333; // @[AWSVggWrapper.scala 52:94]
  wire [815:0] _T_334; // @[AWSVggWrapper.scala 52:94]
  wire [831:0] _T_335; // @[AWSVggWrapper.scala 52:94]
  wire [847:0] _T_336; // @[AWSVggWrapper.scala 52:94]
  wire [863:0] _T_337; // @[AWSVggWrapper.scala 52:94]
  wire [879:0] _T_338; // @[AWSVggWrapper.scala 52:94]
  wire [895:0] _T_339; // @[AWSVggWrapper.scala 52:94]
  wire [911:0] _T_340; // @[AWSVggWrapper.scala 52:94]
  wire [927:0] _T_341; // @[AWSVggWrapper.scala 52:94]
  wire [943:0] _T_342; // @[AWSVggWrapper.scala 52:94]
  wire [959:0] _T_343; // @[AWSVggWrapper.scala 52:94]
  wire [975:0] _T_344; // @[AWSVggWrapper.scala 52:94]
  wire [991:0] _T_345; // @[AWSVggWrapper.scala 52:94]
  wire [1007:0] _T_346; // @[AWSVggWrapper.scala 52:94]
  wire [1023:0] _T_347; // @[AWSVggWrapper.scala 52:94]
  wire [1039:0] _T_348; // @[AWSVggWrapper.scala 52:94]
  wire [1055:0] _T_349; // @[AWSVggWrapper.scala 52:94]
  wire [1071:0] _T_350; // @[AWSVggWrapper.scala 52:94]
  wire [1087:0] _T_351; // @[AWSVggWrapper.scala 52:94]
  wire [1103:0] _T_352; // @[AWSVggWrapper.scala 52:94]
  wire [1119:0] _T_353; // @[AWSVggWrapper.scala 52:94]
  wire [1135:0] _T_354; // @[AWSVggWrapper.scala 52:94]
  wire [1151:0] _T_355; // @[AWSVggWrapper.scala 52:94]
  wire [1167:0] _T_356; // @[AWSVggWrapper.scala 52:94]
  wire [1183:0] _T_357; // @[AWSVggWrapper.scala 52:94]
  wire [1199:0] _T_358; // @[AWSVggWrapper.scala 52:94]
  wire [1215:0] _T_359; // @[AWSVggWrapper.scala 52:94]
  wire [1231:0] _T_360; // @[AWSVggWrapper.scala 52:94]
  wire [1247:0] _T_361; // @[AWSVggWrapper.scala 52:94]
  wire [1263:0] _T_362; // @[AWSVggWrapper.scala 52:94]
  wire [1279:0] _T_363; // @[AWSVggWrapper.scala 52:94]
  wire [1295:0] _T_364; // @[AWSVggWrapper.scala 52:94]
  wire [1311:0] _T_365; // @[AWSVggWrapper.scala 52:94]
  wire [1327:0] _T_366; // @[AWSVggWrapper.scala 52:94]
  wire [1343:0] _T_367; // @[AWSVggWrapper.scala 52:94]
  wire [1359:0] _T_368; // @[AWSVggWrapper.scala 52:94]
  wire [1375:0] _T_369; // @[AWSVggWrapper.scala 52:94]
  wire [1391:0] _T_370; // @[AWSVggWrapper.scala 52:94]
  wire [1407:0] _T_371; // @[AWSVggWrapper.scala 52:94]
  wire [1423:0] _T_372; // @[AWSVggWrapper.scala 52:94]
  wire [1439:0] _T_373; // @[AWSVggWrapper.scala 52:94]
  wire [1455:0] _T_374; // @[AWSVggWrapper.scala 52:94]
  wire [1471:0] _T_375; // @[AWSVggWrapper.scala 52:94]
  wire [1487:0] _T_376; // @[AWSVggWrapper.scala 52:94]
  wire [1503:0] _T_377; // @[AWSVggWrapper.scala 52:94]
  wire [1519:0] _T_378; // @[AWSVggWrapper.scala 52:94]
  wire [1535:0] _T_379; // @[AWSVggWrapper.scala 52:94]
  wire [1551:0] _T_380; // @[AWSVggWrapper.scala 52:94]
  wire [1567:0] _T_381; // @[AWSVggWrapper.scala 52:94]
  wire [1583:0] _T_382; // @[AWSVggWrapper.scala 52:94]
  wire [1599:0] _T_383; // @[AWSVggWrapper.scala 52:94]
  wire [1615:0] _T_384; // @[AWSVggWrapper.scala 52:94]
  wire [1631:0] _T_385; // @[AWSVggWrapper.scala 52:94]
  wire [1647:0] _T_386; // @[AWSVggWrapper.scala 52:94]
  wire [1663:0] _T_387; // @[AWSVggWrapper.scala 52:94]
  wire [1679:0] _T_388; // @[AWSVggWrapper.scala 52:94]
  wire [1695:0] _T_389; // @[AWSVggWrapper.scala 52:94]
  wire [1711:0] _T_390; // @[AWSVggWrapper.scala 52:94]
  wire [1727:0] _T_391; // @[AWSVggWrapper.scala 52:94]
  wire [1743:0] _T_392; // @[AWSVggWrapper.scala 52:94]
  wire [1759:0] _T_393; // @[AWSVggWrapper.scala 52:94]
  wire [1775:0] _T_394; // @[AWSVggWrapper.scala 52:94]
  wire [1791:0] _T_395; // @[AWSVggWrapper.scala 52:94]
  wire [1807:0] _T_396; // @[AWSVggWrapper.scala 52:94]
  wire [1823:0] _T_397; // @[AWSVggWrapper.scala 52:94]
  wire [1839:0] _T_398; // @[AWSVggWrapper.scala 52:94]
  wire [1855:0] _T_399; // @[AWSVggWrapper.scala 52:94]
  wire [1871:0] _T_400; // @[AWSVggWrapper.scala 52:94]
  wire [1887:0] _T_401; // @[AWSVggWrapper.scala 52:94]
  wire [1903:0] _T_402; // @[AWSVggWrapper.scala 52:94]
  wire [1919:0] _T_403; // @[AWSVggWrapper.scala 52:94]
  wire [1935:0] _T_404; // @[AWSVggWrapper.scala 52:94]
  wire [1951:0] _T_405; // @[AWSVggWrapper.scala 52:94]
  wire [1967:0] _T_406; // @[AWSVggWrapper.scala 52:94]
  wire [1983:0] _T_407; // @[AWSVggWrapper.scala 52:94]
  wire [1999:0] _T_408; // @[AWSVggWrapper.scala 52:94]
  wire [2015:0] _T_409; // @[AWSVggWrapper.scala 52:94]
  wire [2031:0] _T_410; // @[AWSVggWrapper.scala 52:94]
  wire [2047:0] _T_411; // @[AWSVggWrapper.scala 52:94]
  wire [2063:0] _T_412; // @[AWSVggWrapper.scala 52:94]
  wire [2079:0] _T_413; // @[AWSVggWrapper.scala 52:94]
  wire [2095:0] _T_414; // @[AWSVggWrapper.scala 52:94]
  wire [2111:0] _T_415; // @[AWSVggWrapper.scala 52:94]
  wire [2127:0] _T_416; // @[AWSVggWrapper.scala 52:94]
  wire [2143:0] _T_417; // @[AWSVggWrapper.scala 52:94]
  wire [2159:0] _T_418; // @[AWSVggWrapper.scala 52:94]
  wire [2175:0] _T_419; // @[AWSVggWrapper.scala 52:94]
  wire [2191:0] _T_420; // @[AWSVggWrapper.scala 52:94]
  wire [2207:0] _T_421; // @[AWSVggWrapper.scala 52:94]
  wire [2223:0] _T_422; // @[AWSVggWrapper.scala 52:94]
  wire [2239:0] _T_423; // @[AWSVggWrapper.scala 52:94]
  wire [2255:0] _T_424; // @[AWSVggWrapper.scala 52:94]
  wire [2271:0] _T_425; // @[AWSVggWrapper.scala 52:94]
  wire [2287:0] _T_426; // @[AWSVggWrapper.scala 52:94]
  wire [2303:0] _T_427; // @[AWSVggWrapper.scala 52:94]
  wire [2319:0] _T_428; // @[AWSVggWrapper.scala 52:94]
  wire [2335:0] _T_429; // @[AWSVggWrapper.scala 52:94]
  wire [2351:0] _T_430; // @[AWSVggWrapper.scala 52:94]
  wire [2367:0] _T_431; // @[AWSVggWrapper.scala 52:94]
  wire [2383:0] _T_432; // @[AWSVggWrapper.scala 52:94]
  wire [2399:0] _T_433; // @[AWSVggWrapper.scala 52:94]
  wire [2415:0] _T_434; // @[AWSVggWrapper.scala 52:94]
  wire [2431:0] _T_435; // @[AWSVggWrapper.scala 52:94]
  wire [2447:0] _T_436; // @[AWSVggWrapper.scala 52:94]
  wire [2463:0] _T_437; // @[AWSVggWrapper.scala 52:94]
  wire [2479:0] _T_438; // @[AWSVggWrapper.scala 52:94]
  wire [2495:0] _T_439; // @[AWSVggWrapper.scala 52:94]
  wire [2511:0] _T_440; // @[AWSVggWrapper.scala 52:94]
  wire [2527:0] _T_441; // @[AWSVggWrapper.scala 52:94]
  wire [2543:0] _T_442; // @[AWSVggWrapper.scala 52:94]
  wire [2559:0] _T_443; // @[AWSVggWrapper.scala 52:94]
  wire [2575:0] _T_444; // @[AWSVggWrapper.scala 52:94]
  wire [2591:0] _T_445; // @[AWSVggWrapper.scala 52:94]
  wire [2607:0] _T_446; // @[AWSVggWrapper.scala 52:94]
  wire [2623:0] _T_447; // @[AWSVggWrapper.scala 52:94]
  wire [2639:0] _T_448; // @[AWSVggWrapper.scala 52:94]
  wire [2655:0] _T_449; // @[AWSVggWrapper.scala 52:94]
  wire [2671:0] _T_450; // @[AWSVggWrapper.scala 52:94]
  wire [2687:0] _T_451; // @[AWSVggWrapper.scala 52:94]
  wire [2703:0] _T_452; // @[AWSVggWrapper.scala 52:94]
  wire [2719:0] _T_453; // @[AWSVggWrapper.scala 52:94]
  wire [2735:0] _T_454; // @[AWSVggWrapper.scala 52:94]
  wire [2751:0] _T_455; // @[AWSVggWrapper.scala 52:94]
  wire [2767:0] _T_456; // @[AWSVggWrapper.scala 52:94]
  wire [2783:0] _T_457; // @[AWSVggWrapper.scala 52:94]
  wire [2799:0] _T_458; // @[AWSVggWrapper.scala 52:94]
  wire [2815:0] _T_459; // @[AWSVggWrapper.scala 52:94]
  wire [2831:0] _T_460; // @[AWSVggWrapper.scala 52:94]
  wire [2847:0] _T_461; // @[AWSVggWrapper.scala 52:94]
  wire [2863:0] _T_462; // @[AWSVggWrapper.scala 52:94]
  wire [2879:0] _T_463; // @[AWSVggWrapper.scala 52:94]
  wire [2895:0] _T_464; // @[AWSVggWrapper.scala 52:94]
  wire [2911:0] _T_465; // @[AWSVggWrapper.scala 52:94]
  wire [2927:0] _T_466; // @[AWSVggWrapper.scala 52:94]
  wire [2943:0] _T_467; // @[AWSVggWrapper.scala 52:94]
  wire [2959:0] _T_468; // @[AWSVggWrapper.scala 52:94]
  wire [2975:0] _T_469; // @[AWSVggWrapper.scala 52:94]
  wire [2991:0] _T_470; // @[AWSVggWrapper.scala 52:94]
  wire [3007:0] _T_471; // @[AWSVggWrapper.scala 52:94]
  wire [3023:0] _T_472; // @[AWSVggWrapper.scala 52:94]
  wire [3039:0] _T_473; // @[AWSVggWrapper.scala 52:94]
  wire [3055:0] _T_474; // @[AWSVggWrapper.scala 52:94]
  wire [3071:0] _T_475; // @[AWSVggWrapper.scala 52:94]
  wire [3087:0] _T_476; // @[AWSVggWrapper.scala 52:94]
  wire [3103:0] _T_477; // @[AWSVggWrapper.scala 52:94]
  wire [3119:0] _T_478; // @[AWSVggWrapper.scala 52:94]
  wire [3135:0] _T_479; // @[AWSVggWrapper.scala 52:94]
  wire [3151:0] _T_480; // @[AWSVggWrapper.scala 52:94]
  wire [3167:0] _T_481; // @[AWSVggWrapper.scala 52:94]
  wire [3183:0] _T_482; // @[AWSVggWrapper.scala 52:94]
  wire [3199:0] _T_483; // @[AWSVggWrapper.scala 52:94]
  wire [3215:0] _T_484; // @[AWSVggWrapper.scala 52:94]
  wire [3231:0] _T_485; // @[AWSVggWrapper.scala 52:94]
  wire [3247:0] _T_486; // @[AWSVggWrapper.scala 52:94]
  wire [3263:0] _T_487; // @[AWSVggWrapper.scala 52:94]
  wire [3279:0] _T_488; // @[AWSVggWrapper.scala 52:94]
  wire [3295:0] _T_489; // @[AWSVggWrapper.scala 52:94]
  wire [3311:0] _T_490; // @[AWSVggWrapper.scala 52:94]
  wire [3327:0] _T_491; // @[AWSVggWrapper.scala 52:94]
  wire [3343:0] _T_492; // @[AWSVggWrapper.scala 52:94]
  wire [3359:0] _T_493; // @[AWSVggWrapper.scala 52:94]
  wire [3375:0] _T_494; // @[AWSVggWrapper.scala 52:94]
  wire [3391:0] _T_495; // @[AWSVggWrapper.scala 52:94]
  wire [3407:0] _T_496; // @[AWSVggWrapper.scala 52:94]
  wire [3423:0] _T_497; // @[AWSVggWrapper.scala 52:94]
  wire [3439:0] _T_498; // @[AWSVggWrapper.scala 52:94]
  wire [3455:0] _T_499; // @[AWSVggWrapper.scala 52:94]
  wire [3471:0] _T_500; // @[AWSVggWrapper.scala 52:94]
  wire [3487:0] _T_501; // @[AWSVggWrapper.scala 52:94]
  wire [3503:0] _T_502; // @[AWSVggWrapper.scala 52:94]
  wire [3519:0] _T_503; // @[AWSVggWrapper.scala 52:94]
  wire [3535:0] _T_504; // @[AWSVggWrapper.scala 52:94]
  wire [3551:0] _T_505; // @[AWSVggWrapper.scala 52:94]
  wire [3567:0] _T_506; // @[AWSVggWrapper.scala 52:94]
  wire [3583:0] _T_507; // @[AWSVggWrapper.scala 52:94]
  wire [3599:0] _T_508; // @[AWSVggWrapper.scala 52:94]
  wire [3615:0] _T_509; // @[AWSVggWrapper.scala 52:94]
  wire [3631:0] _T_510; // @[AWSVggWrapper.scala 52:94]
  wire [3647:0] _T_511; // @[AWSVggWrapper.scala 52:94]
  wire [3663:0] _T_512; // @[AWSVggWrapper.scala 52:94]
  wire [3679:0] _T_513; // @[AWSVggWrapper.scala 52:94]
  wire [3695:0] _T_514; // @[AWSVggWrapper.scala 52:94]
  wire [3711:0] _T_515; // @[AWSVggWrapper.scala 52:94]
  wire [3727:0] _T_516; // @[AWSVggWrapper.scala 52:94]
  wire [3743:0] _T_517; // @[AWSVggWrapper.scala 52:94]
  wire [3759:0] _T_518; // @[AWSVggWrapper.scala 52:94]
  wire [3775:0] _T_519; // @[AWSVggWrapper.scala 52:94]
  wire [3791:0] _T_520; // @[AWSVggWrapper.scala 52:94]
  wire [3807:0] _T_521; // @[AWSVggWrapper.scala 52:94]
  wire [3823:0] _T_522; // @[AWSVggWrapper.scala 52:94]
  wire [3839:0] _T_523; // @[AWSVggWrapper.scala 52:94]
  wire [3855:0] _T_524; // @[AWSVggWrapper.scala 52:94]
  wire [3871:0] _T_525; // @[AWSVggWrapper.scala 52:94]
  wire [3887:0] _T_526; // @[AWSVggWrapper.scala 52:94]
  wire [3903:0] _T_527; // @[AWSVggWrapper.scala 52:94]
  wire [3919:0] _T_528; // @[AWSVggWrapper.scala 52:94]
  wire [3935:0] _T_529; // @[AWSVggWrapper.scala 52:94]
  wire [3951:0] _T_530; // @[AWSVggWrapper.scala 52:94]
  wire [3967:0] _T_531; // @[AWSVggWrapper.scala 52:94]
  wire [3983:0] _T_532; // @[AWSVggWrapper.scala 52:94]
  wire [3999:0] _T_533; // @[AWSVggWrapper.scala 52:94]
  wire [4015:0] _T_534; // @[AWSVggWrapper.scala 52:94]
  wire [4031:0] _T_535; // @[AWSVggWrapper.scala 52:94]
  wire [4047:0] _T_536; // @[AWSVggWrapper.scala 52:94]
  wire [4063:0] _T_537; // @[AWSVggWrapper.scala 52:94]
  wire [4079:0] _T_538; // @[AWSVggWrapper.scala 52:94]
  wire [4095:0] dataInAsUInt; // @[AWSVggWrapper.scala 52:94]
  wire [15:0] _T_1833; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_255; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1835; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_254; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1837; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_253; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1839; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_252; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1841; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_251; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1843; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_250; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1845; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_249; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1847; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_248; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1849; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_247; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1851; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_246; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1853; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_245; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1855; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_244; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1857; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_243; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1859; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_242; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1861; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_241; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1863; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_240; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1865; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_239; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1867; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_238; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1869; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_237; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1871; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_236; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1873; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_235; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1875; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_234; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1877; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_233; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1879; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_232; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1881; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_231; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1883; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_230; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1885; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_229; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1887; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_228; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1889; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_227; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1891; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_226; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1893; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_225; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1895; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_224; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1897; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_223; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1899; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_222; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1901; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_221; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1903; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_220; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1905; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_219; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1907; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_218; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1909; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_217; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1911; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_216; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1913; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_215; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1915; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_214; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1917; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_213; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1919; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_212; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1921; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_211; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1923; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_210; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1925; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_209; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1927; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_208; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1929; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_207; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1931; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_206; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1933; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_205; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1935; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_204; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1937; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_203; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1939; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_202; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1941; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_201; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1943; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_200; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1945; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_199; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1947; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_198; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1949; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_197; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1951; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_196; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1953; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_195; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1955; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_194; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1957; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_193; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1959; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_192; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1961; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_191; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1963; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_190; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1965; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_189; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1967; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_188; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1969; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_187; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1971; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_186; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1973; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_185; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1975; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_184; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1977; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_183; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1979; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_182; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1981; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_181; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1983; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_180; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1985; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_179; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1987; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_178; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1989; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_177; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1991; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_176; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1993; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_175; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1995; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_174; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1997; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_173; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_1999; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_172; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2001; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_171; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2003; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_170; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2005; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_169; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2007; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_168; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2009; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_167; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2011; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_166; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2013; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_165; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2015; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_164; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2017; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_163; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2019; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_162; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2021; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_161; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2023; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_160; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2025; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_159; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2027; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_158; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2029; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_157; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2031; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_156; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2033; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_155; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2035; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_154; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2037; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_153; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2039; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_152; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2041; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_151; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2043; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_150; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2045; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_149; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2047; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_148; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2049; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_147; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2051; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_146; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2053; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_145; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2055; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_144; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2057; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_143; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2059; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_142; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2061; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_141; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2063; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_140; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2065; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_139; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2067; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_138; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2069; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_137; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2071; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_136; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2073; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_135; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2075; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_134; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2077; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_133; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2079; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_132; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2081; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_131; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2083; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_130; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2085; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_129; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2087; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_128; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2089; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_127; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2091; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_126; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2093; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_125; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2095; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_124; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2097; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_123; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2099; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_122; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2101; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_121; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2103; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_120; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2105; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_119; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2107; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_118; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2109; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_117; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2111; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_116; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2113; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_115; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2115; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_114; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2117; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_113; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2119; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_112; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2121; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_111; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2123; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_110; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2125; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_109; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2127; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_108; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2129; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_107; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2131; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_106; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2133; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_105; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2135; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_104; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2137; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_103; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2139; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_102; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2141; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_101; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2143; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_100; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2145; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_99; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2147; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_98; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2149; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_97; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2151; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_96; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2153; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_95; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2155; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_94; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2157; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_93; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2159; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_92; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2161; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_91; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2163; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_90; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2165; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_89; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2167; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_88; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2169; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_87; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2171; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_86; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2173; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_85; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2175; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_84; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2177; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_83; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2179; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_82; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2181; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_81; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2183; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_80; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2185; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_79; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2187; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_78; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2189; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_77; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2191; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_76; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2193; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_75; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2195; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_74; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2197; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_73; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2199; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_72; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2201; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_71; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2203; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_70; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2205; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_69; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2207; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_68; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2209; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_67; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2211; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_66; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2213; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_65; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2215; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_64; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2217; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_63; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2219; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_62; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2221; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_61; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2223; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_60; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2225; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_59; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2227; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_58; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2229; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_57; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2231; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_56; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2233; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_55; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2235; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_54; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2237; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_53; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2239; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_52; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2241; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_51; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2243; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_50; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2245; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_49; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2247; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_48; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2249; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_47; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2251; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_46; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2253; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_45; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2255; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_44; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2257; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_43; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2259; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_42; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2261; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_41; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2263; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_40; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2265; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_39; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2267; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_38; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2269; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_37; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2271; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_36; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2273; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_35; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2275; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_34; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2277; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_33; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2279; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_32; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2281; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_31; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2283; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_30; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2285; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_29; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2287; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_28; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2289; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_27; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2291; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_26; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2293; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_25; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2295; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_24; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2297; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_23; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2299; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_22; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2301; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_21; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2303; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_20; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2305; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_19; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2307; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_18; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2309; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_17; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2311; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_16; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2313; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_15; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2315; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_14; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2317; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_13; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2319; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_12; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2321; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_11; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2323; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_10; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2325; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_9; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2327; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_8; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2329; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_7; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2331; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_6; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2333; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_5; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2335; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_4; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2337; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_3; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2339; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_2; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2341; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_1; // @[AWSVggWrapper.scala 63:110]
  wire [15:0] _T_2343; // @[AWSVggWrapper.scala 63:67]
  wire [15:0] sintOut_0; // @[AWSVggWrapper.scala 63:110]
  wire  queueIOIn_ready; // @[AWSVggWrapper.scala 53:23]
  wire  queueIOIn_valid; // @[AWSVggWrapper.scala 53:23]
  Vgg7 vgg ( // @[AWSVggWrapper.scala 46:27]
    .clock(vgg_clock),
    .reset(vgg_reset),
    .io_dataIn_ready(vgg_io_dataIn_ready),
    .io_dataIn_valid(vgg_io_dataIn_valid),
    .io_dataIn_bits_0(vgg_io_dataIn_bits_0),
    .io_dataIn_bits_1(vgg_io_dataIn_bits_1),
    .io_dataIn_bits_2(vgg_io_dataIn_bits_2),
    .io_dataOut_ready(vgg_io_dataOut_ready),
    .io_dataOut_valid(vgg_io_dataOut_valid),
    .io_dataOut_bits_0(vgg_io_dataOut_bits_0),
    .io_dataOut_bits_1(vgg_io_dataOut_bits_1),
    .io_dataOut_bits_2(vgg_io_dataOut_bits_2),
    .io_dataOut_bits_3(vgg_io_dataOut_bits_3),
    .io_dataOut_bits_4(vgg_io_dataOut_bits_4),
    .io_dataOut_bits_5(vgg_io_dataOut_bits_5),
    .io_dataOut_bits_6(vgg_io_dataOut_bits_6),
    .io_dataOut_bits_7(vgg_io_dataOut_bits_7),
    .io_dataOut_bits_8(vgg_io_dataOut_bits_8),
    .io_dataOut_bits_9(vgg_io_dataOut_bits_9),
    .io_dataOut_bits_10(vgg_io_dataOut_bits_10),
    .io_dataOut_bits_11(vgg_io_dataOut_bits_11),
    .io_dataOut_bits_12(vgg_io_dataOut_bits_12),
    .io_dataOut_bits_13(vgg_io_dataOut_bits_13),
    .io_dataOut_bits_14(vgg_io_dataOut_bits_14),
    .io_dataOut_bits_15(vgg_io_dataOut_bits_15),
    .io_dataOut_bits_16(vgg_io_dataOut_bits_16),
    .io_dataOut_bits_17(vgg_io_dataOut_bits_17),
    .io_dataOut_bits_18(vgg_io_dataOut_bits_18),
    .io_dataOut_bits_19(vgg_io_dataOut_bits_19),
    .io_dataOut_bits_20(vgg_io_dataOut_bits_20),
    .io_dataOut_bits_21(vgg_io_dataOut_bits_21),
    .io_dataOut_bits_22(vgg_io_dataOut_bits_22),
    .io_dataOut_bits_23(vgg_io_dataOut_bits_23),
    .io_dataOut_bits_24(vgg_io_dataOut_bits_24),
    .io_dataOut_bits_25(vgg_io_dataOut_bits_25),
    .io_dataOut_bits_26(vgg_io_dataOut_bits_26),
    .io_dataOut_bits_27(vgg_io_dataOut_bits_27),
    .io_dataOut_bits_28(vgg_io_dataOut_bits_28),
    .io_dataOut_bits_29(vgg_io_dataOut_bits_29),
    .io_dataOut_bits_30(vgg_io_dataOut_bits_30),
    .io_dataOut_bits_31(vgg_io_dataOut_bits_31),
    .io_dataOut_bits_32(vgg_io_dataOut_bits_32),
    .io_dataOut_bits_33(vgg_io_dataOut_bits_33),
    .io_dataOut_bits_34(vgg_io_dataOut_bits_34),
    .io_dataOut_bits_35(vgg_io_dataOut_bits_35),
    .io_dataOut_bits_36(vgg_io_dataOut_bits_36),
    .io_dataOut_bits_37(vgg_io_dataOut_bits_37),
    .io_dataOut_bits_38(vgg_io_dataOut_bits_38),
    .io_dataOut_bits_39(vgg_io_dataOut_bits_39),
    .io_dataOut_bits_40(vgg_io_dataOut_bits_40),
    .io_dataOut_bits_41(vgg_io_dataOut_bits_41),
    .io_dataOut_bits_42(vgg_io_dataOut_bits_42),
    .io_dataOut_bits_43(vgg_io_dataOut_bits_43),
    .io_dataOut_bits_44(vgg_io_dataOut_bits_44),
    .io_dataOut_bits_45(vgg_io_dataOut_bits_45),
    .io_dataOut_bits_46(vgg_io_dataOut_bits_46),
    .io_dataOut_bits_47(vgg_io_dataOut_bits_47),
    .io_dataOut_bits_48(vgg_io_dataOut_bits_48),
    .io_dataOut_bits_49(vgg_io_dataOut_bits_49),
    .io_dataOut_bits_50(vgg_io_dataOut_bits_50),
    .io_dataOut_bits_51(vgg_io_dataOut_bits_51),
    .io_dataOut_bits_52(vgg_io_dataOut_bits_52),
    .io_dataOut_bits_53(vgg_io_dataOut_bits_53),
    .io_dataOut_bits_54(vgg_io_dataOut_bits_54),
    .io_dataOut_bits_55(vgg_io_dataOut_bits_55),
    .io_dataOut_bits_56(vgg_io_dataOut_bits_56),
    .io_dataOut_bits_57(vgg_io_dataOut_bits_57),
    .io_dataOut_bits_58(vgg_io_dataOut_bits_58),
    .io_dataOut_bits_59(vgg_io_dataOut_bits_59),
    .io_dataOut_bits_60(vgg_io_dataOut_bits_60),
    .io_dataOut_bits_61(vgg_io_dataOut_bits_61),
    .io_dataOut_bits_62(vgg_io_dataOut_bits_62),
    .io_dataOut_bits_63(vgg_io_dataOut_bits_63),
    .io_dataOut_bits_64(vgg_io_dataOut_bits_64),
    .io_dataOut_bits_65(vgg_io_dataOut_bits_65),
    .io_dataOut_bits_66(vgg_io_dataOut_bits_66),
    .io_dataOut_bits_67(vgg_io_dataOut_bits_67),
    .io_dataOut_bits_68(vgg_io_dataOut_bits_68),
    .io_dataOut_bits_69(vgg_io_dataOut_bits_69),
    .io_dataOut_bits_70(vgg_io_dataOut_bits_70),
    .io_dataOut_bits_71(vgg_io_dataOut_bits_71),
    .io_dataOut_bits_72(vgg_io_dataOut_bits_72),
    .io_dataOut_bits_73(vgg_io_dataOut_bits_73),
    .io_dataOut_bits_74(vgg_io_dataOut_bits_74),
    .io_dataOut_bits_75(vgg_io_dataOut_bits_75),
    .io_dataOut_bits_76(vgg_io_dataOut_bits_76),
    .io_dataOut_bits_77(vgg_io_dataOut_bits_77),
    .io_dataOut_bits_78(vgg_io_dataOut_bits_78),
    .io_dataOut_bits_79(vgg_io_dataOut_bits_79),
    .io_dataOut_bits_80(vgg_io_dataOut_bits_80),
    .io_dataOut_bits_81(vgg_io_dataOut_bits_81),
    .io_dataOut_bits_82(vgg_io_dataOut_bits_82),
    .io_dataOut_bits_83(vgg_io_dataOut_bits_83),
    .io_dataOut_bits_84(vgg_io_dataOut_bits_84),
    .io_dataOut_bits_85(vgg_io_dataOut_bits_85),
    .io_dataOut_bits_86(vgg_io_dataOut_bits_86),
    .io_dataOut_bits_87(vgg_io_dataOut_bits_87),
    .io_dataOut_bits_88(vgg_io_dataOut_bits_88),
    .io_dataOut_bits_89(vgg_io_dataOut_bits_89),
    .io_dataOut_bits_90(vgg_io_dataOut_bits_90),
    .io_dataOut_bits_91(vgg_io_dataOut_bits_91),
    .io_dataOut_bits_92(vgg_io_dataOut_bits_92),
    .io_dataOut_bits_93(vgg_io_dataOut_bits_93),
    .io_dataOut_bits_94(vgg_io_dataOut_bits_94),
    .io_dataOut_bits_95(vgg_io_dataOut_bits_95),
    .io_dataOut_bits_96(vgg_io_dataOut_bits_96),
    .io_dataOut_bits_97(vgg_io_dataOut_bits_97),
    .io_dataOut_bits_98(vgg_io_dataOut_bits_98),
    .io_dataOut_bits_99(vgg_io_dataOut_bits_99),
    .io_dataOut_bits_100(vgg_io_dataOut_bits_100),
    .io_dataOut_bits_101(vgg_io_dataOut_bits_101),
    .io_dataOut_bits_102(vgg_io_dataOut_bits_102),
    .io_dataOut_bits_103(vgg_io_dataOut_bits_103),
    .io_dataOut_bits_104(vgg_io_dataOut_bits_104),
    .io_dataOut_bits_105(vgg_io_dataOut_bits_105),
    .io_dataOut_bits_106(vgg_io_dataOut_bits_106),
    .io_dataOut_bits_107(vgg_io_dataOut_bits_107),
    .io_dataOut_bits_108(vgg_io_dataOut_bits_108),
    .io_dataOut_bits_109(vgg_io_dataOut_bits_109),
    .io_dataOut_bits_110(vgg_io_dataOut_bits_110),
    .io_dataOut_bits_111(vgg_io_dataOut_bits_111),
    .io_dataOut_bits_112(vgg_io_dataOut_bits_112),
    .io_dataOut_bits_113(vgg_io_dataOut_bits_113),
    .io_dataOut_bits_114(vgg_io_dataOut_bits_114),
    .io_dataOut_bits_115(vgg_io_dataOut_bits_115),
    .io_dataOut_bits_116(vgg_io_dataOut_bits_116),
    .io_dataOut_bits_117(vgg_io_dataOut_bits_117),
    .io_dataOut_bits_118(vgg_io_dataOut_bits_118),
    .io_dataOut_bits_119(vgg_io_dataOut_bits_119),
    .io_dataOut_bits_120(vgg_io_dataOut_bits_120),
    .io_dataOut_bits_121(vgg_io_dataOut_bits_121),
    .io_dataOut_bits_122(vgg_io_dataOut_bits_122),
    .io_dataOut_bits_123(vgg_io_dataOut_bits_123),
    .io_dataOut_bits_124(vgg_io_dataOut_bits_124),
    .io_dataOut_bits_125(vgg_io_dataOut_bits_125),
    .io_dataOut_bits_126(vgg_io_dataOut_bits_126),
    .io_dataOut_bits_127(vgg_io_dataOut_bits_127),
    .io_dataOut_bits_128(vgg_io_dataOut_bits_128),
    .io_dataOut_bits_129(vgg_io_dataOut_bits_129),
    .io_dataOut_bits_130(vgg_io_dataOut_bits_130),
    .io_dataOut_bits_131(vgg_io_dataOut_bits_131),
    .io_dataOut_bits_132(vgg_io_dataOut_bits_132),
    .io_dataOut_bits_133(vgg_io_dataOut_bits_133),
    .io_dataOut_bits_134(vgg_io_dataOut_bits_134),
    .io_dataOut_bits_135(vgg_io_dataOut_bits_135),
    .io_dataOut_bits_136(vgg_io_dataOut_bits_136),
    .io_dataOut_bits_137(vgg_io_dataOut_bits_137),
    .io_dataOut_bits_138(vgg_io_dataOut_bits_138),
    .io_dataOut_bits_139(vgg_io_dataOut_bits_139),
    .io_dataOut_bits_140(vgg_io_dataOut_bits_140),
    .io_dataOut_bits_141(vgg_io_dataOut_bits_141),
    .io_dataOut_bits_142(vgg_io_dataOut_bits_142),
    .io_dataOut_bits_143(vgg_io_dataOut_bits_143),
    .io_dataOut_bits_144(vgg_io_dataOut_bits_144),
    .io_dataOut_bits_145(vgg_io_dataOut_bits_145),
    .io_dataOut_bits_146(vgg_io_dataOut_bits_146),
    .io_dataOut_bits_147(vgg_io_dataOut_bits_147),
    .io_dataOut_bits_148(vgg_io_dataOut_bits_148),
    .io_dataOut_bits_149(vgg_io_dataOut_bits_149),
    .io_dataOut_bits_150(vgg_io_dataOut_bits_150),
    .io_dataOut_bits_151(vgg_io_dataOut_bits_151),
    .io_dataOut_bits_152(vgg_io_dataOut_bits_152),
    .io_dataOut_bits_153(vgg_io_dataOut_bits_153),
    .io_dataOut_bits_154(vgg_io_dataOut_bits_154),
    .io_dataOut_bits_155(vgg_io_dataOut_bits_155),
    .io_dataOut_bits_156(vgg_io_dataOut_bits_156),
    .io_dataOut_bits_157(vgg_io_dataOut_bits_157),
    .io_dataOut_bits_158(vgg_io_dataOut_bits_158),
    .io_dataOut_bits_159(vgg_io_dataOut_bits_159),
    .io_dataOut_bits_160(vgg_io_dataOut_bits_160),
    .io_dataOut_bits_161(vgg_io_dataOut_bits_161),
    .io_dataOut_bits_162(vgg_io_dataOut_bits_162),
    .io_dataOut_bits_163(vgg_io_dataOut_bits_163),
    .io_dataOut_bits_164(vgg_io_dataOut_bits_164),
    .io_dataOut_bits_165(vgg_io_dataOut_bits_165),
    .io_dataOut_bits_166(vgg_io_dataOut_bits_166),
    .io_dataOut_bits_167(vgg_io_dataOut_bits_167),
    .io_dataOut_bits_168(vgg_io_dataOut_bits_168),
    .io_dataOut_bits_169(vgg_io_dataOut_bits_169),
    .io_dataOut_bits_170(vgg_io_dataOut_bits_170),
    .io_dataOut_bits_171(vgg_io_dataOut_bits_171),
    .io_dataOut_bits_172(vgg_io_dataOut_bits_172),
    .io_dataOut_bits_173(vgg_io_dataOut_bits_173),
    .io_dataOut_bits_174(vgg_io_dataOut_bits_174),
    .io_dataOut_bits_175(vgg_io_dataOut_bits_175),
    .io_dataOut_bits_176(vgg_io_dataOut_bits_176),
    .io_dataOut_bits_177(vgg_io_dataOut_bits_177),
    .io_dataOut_bits_178(vgg_io_dataOut_bits_178),
    .io_dataOut_bits_179(vgg_io_dataOut_bits_179),
    .io_dataOut_bits_180(vgg_io_dataOut_bits_180),
    .io_dataOut_bits_181(vgg_io_dataOut_bits_181),
    .io_dataOut_bits_182(vgg_io_dataOut_bits_182),
    .io_dataOut_bits_183(vgg_io_dataOut_bits_183),
    .io_dataOut_bits_184(vgg_io_dataOut_bits_184),
    .io_dataOut_bits_185(vgg_io_dataOut_bits_185),
    .io_dataOut_bits_186(vgg_io_dataOut_bits_186),
    .io_dataOut_bits_187(vgg_io_dataOut_bits_187),
    .io_dataOut_bits_188(vgg_io_dataOut_bits_188),
    .io_dataOut_bits_189(vgg_io_dataOut_bits_189),
    .io_dataOut_bits_190(vgg_io_dataOut_bits_190),
    .io_dataOut_bits_191(vgg_io_dataOut_bits_191),
    .io_dataOut_bits_192(vgg_io_dataOut_bits_192),
    .io_dataOut_bits_193(vgg_io_dataOut_bits_193),
    .io_dataOut_bits_194(vgg_io_dataOut_bits_194),
    .io_dataOut_bits_195(vgg_io_dataOut_bits_195),
    .io_dataOut_bits_196(vgg_io_dataOut_bits_196),
    .io_dataOut_bits_197(vgg_io_dataOut_bits_197),
    .io_dataOut_bits_198(vgg_io_dataOut_bits_198),
    .io_dataOut_bits_199(vgg_io_dataOut_bits_199),
    .io_dataOut_bits_200(vgg_io_dataOut_bits_200),
    .io_dataOut_bits_201(vgg_io_dataOut_bits_201),
    .io_dataOut_bits_202(vgg_io_dataOut_bits_202),
    .io_dataOut_bits_203(vgg_io_dataOut_bits_203),
    .io_dataOut_bits_204(vgg_io_dataOut_bits_204),
    .io_dataOut_bits_205(vgg_io_dataOut_bits_205),
    .io_dataOut_bits_206(vgg_io_dataOut_bits_206),
    .io_dataOut_bits_207(vgg_io_dataOut_bits_207),
    .io_dataOut_bits_208(vgg_io_dataOut_bits_208),
    .io_dataOut_bits_209(vgg_io_dataOut_bits_209),
    .io_dataOut_bits_210(vgg_io_dataOut_bits_210),
    .io_dataOut_bits_211(vgg_io_dataOut_bits_211),
    .io_dataOut_bits_212(vgg_io_dataOut_bits_212),
    .io_dataOut_bits_213(vgg_io_dataOut_bits_213),
    .io_dataOut_bits_214(vgg_io_dataOut_bits_214),
    .io_dataOut_bits_215(vgg_io_dataOut_bits_215),
    .io_dataOut_bits_216(vgg_io_dataOut_bits_216),
    .io_dataOut_bits_217(vgg_io_dataOut_bits_217),
    .io_dataOut_bits_218(vgg_io_dataOut_bits_218),
    .io_dataOut_bits_219(vgg_io_dataOut_bits_219),
    .io_dataOut_bits_220(vgg_io_dataOut_bits_220),
    .io_dataOut_bits_221(vgg_io_dataOut_bits_221),
    .io_dataOut_bits_222(vgg_io_dataOut_bits_222),
    .io_dataOut_bits_223(vgg_io_dataOut_bits_223),
    .io_dataOut_bits_224(vgg_io_dataOut_bits_224),
    .io_dataOut_bits_225(vgg_io_dataOut_bits_225),
    .io_dataOut_bits_226(vgg_io_dataOut_bits_226),
    .io_dataOut_bits_227(vgg_io_dataOut_bits_227),
    .io_dataOut_bits_228(vgg_io_dataOut_bits_228),
    .io_dataOut_bits_229(vgg_io_dataOut_bits_229),
    .io_dataOut_bits_230(vgg_io_dataOut_bits_230),
    .io_dataOut_bits_231(vgg_io_dataOut_bits_231),
    .io_dataOut_bits_232(vgg_io_dataOut_bits_232),
    .io_dataOut_bits_233(vgg_io_dataOut_bits_233),
    .io_dataOut_bits_234(vgg_io_dataOut_bits_234),
    .io_dataOut_bits_235(vgg_io_dataOut_bits_235),
    .io_dataOut_bits_236(vgg_io_dataOut_bits_236),
    .io_dataOut_bits_237(vgg_io_dataOut_bits_237),
    .io_dataOut_bits_238(vgg_io_dataOut_bits_238),
    .io_dataOut_bits_239(vgg_io_dataOut_bits_239),
    .io_dataOut_bits_240(vgg_io_dataOut_bits_240),
    .io_dataOut_bits_241(vgg_io_dataOut_bits_241),
    .io_dataOut_bits_242(vgg_io_dataOut_bits_242),
    .io_dataOut_bits_243(vgg_io_dataOut_bits_243),
    .io_dataOut_bits_244(vgg_io_dataOut_bits_244),
    .io_dataOut_bits_245(vgg_io_dataOut_bits_245),
    .io_dataOut_bits_246(vgg_io_dataOut_bits_246),
    .io_dataOut_bits_247(vgg_io_dataOut_bits_247),
    .io_dataOut_bits_248(vgg_io_dataOut_bits_248),
    .io_dataOut_bits_249(vgg_io_dataOut_bits_249),
    .io_dataOut_bits_250(vgg_io_dataOut_bits_250),
    .io_dataOut_bits_251(vgg_io_dataOut_bits_251),
    .io_dataOut_bits_252(vgg_io_dataOut_bits_252),
    .io_dataOut_bits_253(vgg_io_dataOut_bits_253),
    .io_dataOut_bits_254(vgg_io_dataOut_bits_254),
    .io_dataOut_bits_255(vgg_io_dataOut_bits_255)
  );
  Queue_4096 queueIOOut ( // @[Decoupled.scala 289:19]
    .clock(queueIOOut_clock),
    .reset(queueIOOut_reset),
    .io_enq_ready(queueIOOut_io_enq_ready),
    .io_enq_valid(queueIOOut_io_enq_valid),
    .io_enq_bits(queueIOOut_io_enq_bits),
    .io_deq_ready(queueIOOut_io_deq_ready),
    .io_deq_valid(queueIOOut_io_deq_valid),
    .io_deq_bits(queueIOOut_io_deq_bits)
  );
  MuxLayer muxLyr ( // @[AWSVggWrapper.scala 65:22]
    .clock(muxLyr_clock),
    .reset(muxLyr_reset),
    .io_dataIn_ready(muxLyr_io_dataIn_ready),
    .io_dataIn_valid(muxLyr_io_dataIn_valid),
    .io_dataIn_bits_0(muxLyr_io_dataIn_bits_0),
    .io_dataIn_bits_1(muxLyr_io_dataIn_bits_1),
    .io_dataIn_bits_2(muxLyr_io_dataIn_bits_2),
    .io_dataIn_bits_3(muxLyr_io_dataIn_bits_3),
    .io_dataIn_bits_4(muxLyr_io_dataIn_bits_4),
    .io_dataIn_bits_5(muxLyr_io_dataIn_bits_5),
    .io_dataIn_bits_6(muxLyr_io_dataIn_bits_6),
    .io_dataIn_bits_7(muxLyr_io_dataIn_bits_7),
    .io_dataIn_bits_8(muxLyr_io_dataIn_bits_8),
    .io_dataIn_bits_9(muxLyr_io_dataIn_bits_9),
    .io_dataIn_bits_10(muxLyr_io_dataIn_bits_10),
    .io_dataIn_bits_11(muxLyr_io_dataIn_bits_11),
    .io_dataIn_bits_12(muxLyr_io_dataIn_bits_12),
    .io_dataIn_bits_13(muxLyr_io_dataIn_bits_13),
    .io_dataIn_bits_14(muxLyr_io_dataIn_bits_14),
    .io_dataIn_bits_15(muxLyr_io_dataIn_bits_15),
    .io_dataIn_bits_16(muxLyr_io_dataIn_bits_16),
    .io_dataIn_bits_17(muxLyr_io_dataIn_bits_17),
    .io_dataIn_bits_18(muxLyr_io_dataIn_bits_18),
    .io_dataIn_bits_19(muxLyr_io_dataIn_bits_19),
    .io_dataIn_bits_20(muxLyr_io_dataIn_bits_20),
    .io_dataIn_bits_21(muxLyr_io_dataIn_bits_21),
    .io_dataIn_bits_22(muxLyr_io_dataIn_bits_22),
    .io_dataIn_bits_23(muxLyr_io_dataIn_bits_23),
    .io_dataIn_bits_24(muxLyr_io_dataIn_bits_24),
    .io_dataIn_bits_25(muxLyr_io_dataIn_bits_25),
    .io_dataIn_bits_26(muxLyr_io_dataIn_bits_26),
    .io_dataIn_bits_27(muxLyr_io_dataIn_bits_27),
    .io_dataIn_bits_28(muxLyr_io_dataIn_bits_28),
    .io_dataIn_bits_29(muxLyr_io_dataIn_bits_29),
    .io_dataIn_bits_30(muxLyr_io_dataIn_bits_30),
    .io_dataIn_bits_31(muxLyr_io_dataIn_bits_31),
    .io_dataIn_bits_32(muxLyr_io_dataIn_bits_32),
    .io_dataIn_bits_33(muxLyr_io_dataIn_bits_33),
    .io_dataIn_bits_34(muxLyr_io_dataIn_bits_34),
    .io_dataIn_bits_35(muxLyr_io_dataIn_bits_35),
    .io_dataIn_bits_36(muxLyr_io_dataIn_bits_36),
    .io_dataIn_bits_37(muxLyr_io_dataIn_bits_37),
    .io_dataIn_bits_38(muxLyr_io_dataIn_bits_38),
    .io_dataIn_bits_39(muxLyr_io_dataIn_bits_39),
    .io_dataIn_bits_40(muxLyr_io_dataIn_bits_40),
    .io_dataIn_bits_41(muxLyr_io_dataIn_bits_41),
    .io_dataIn_bits_42(muxLyr_io_dataIn_bits_42),
    .io_dataIn_bits_43(muxLyr_io_dataIn_bits_43),
    .io_dataIn_bits_44(muxLyr_io_dataIn_bits_44),
    .io_dataIn_bits_45(muxLyr_io_dataIn_bits_45),
    .io_dataIn_bits_46(muxLyr_io_dataIn_bits_46),
    .io_dataIn_bits_47(muxLyr_io_dataIn_bits_47),
    .io_dataIn_bits_48(muxLyr_io_dataIn_bits_48),
    .io_dataIn_bits_49(muxLyr_io_dataIn_bits_49),
    .io_dataIn_bits_50(muxLyr_io_dataIn_bits_50),
    .io_dataIn_bits_51(muxLyr_io_dataIn_bits_51),
    .io_dataIn_bits_52(muxLyr_io_dataIn_bits_52),
    .io_dataIn_bits_53(muxLyr_io_dataIn_bits_53),
    .io_dataIn_bits_54(muxLyr_io_dataIn_bits_54),
    .io_dataIn_bits_55(muxLyr_io_dataIn_bits_55),
    .io_dataIn_bits_56(muxLyr_io_dataIn_bits_56),
    .io_dataIn_bits_57(muxLyr_io_dataIn_bits_57),
    .io_dataIn_bits_58(muxLyr_io_dataIn_bits_58),
    .io_dataIn_bits_59(muxLyr_io_dataIn_bits_59),
    .io_dataIn_bits_60(muxLyr_io_dataIn_bits_60),
    .io_dataIn_bits_61(muxLyr_io_dataIn_bits_61),
    .io_dataIn_bits_62(muxLyr_io_dataIn_bits_62),
    .io_dataIn_bits_63(muxLyr_io_dataIn_bits_63),
    .io_dataIn_bits_64(muxLyr_io_dataIn_bits_64),
    .io_dataIn_bits_65(muxLyr_io_dataIn_bits_65),
    .io_dataIn_bits_66(muxLyr_io_dataIn_bits_66),
    .io_dataIn_bits_67(muxLyr_io_dataIn_bits_67),
    .io_dataIn_bits_68(muxLyr_io_dataIn_bits_68),
    .io_dataIn_bits_69(muxLyr_io_dataIn_bits_69),
    .io_dataIn_bits_70(muxLyr_io_dataIn_bits_70),
    .io_dataIn_bits_71(muxLyr_io_dataIn_bits_71),
    .io_dataIn_bits_72(muxLyr_io_dataIn_bits_72),
    .io_dataIn_bits_73(muxLyr_io_dataIn_bits_73),
    .io_dataIn_bits_74(muxLyr_io_dataIn_bits_74),
    .io_dataIn_bits_75(muxLyr_io_dataIn_bits_75),
    .io_dataIn_bits_76(muxLyr_io_dataIn_bits_76),
    .io_dataIn_bits_77(muxLyr_io_dataIn_bits_77),
    .io_dataIn_bits_78(muxLyr_io_dataIn_bits_78),
    .io_dataIn_bits_79(muxLyr_io_dataIn_bits_79),
    .io_dataIn_bits_80(muxLyr_io_dataIn_bits_80),
    .io_dataIn_bits_81(muxLyr_io_dataIn_bits_81),
    .io_dataIn_bits_82(muxLyr_io_dataIn_bits_82),
    .io_dataIn_bits_83(muxLyr_io_dataIn_bits_83),
    .io_dataIn_bits_84(muxLyr_io_dataIn_bits_84),
    .io_dataIn_bits_85(muxLyr_io_dataIn_bits_85),
    .io_dataIn_bits_86(muxLyr_io_dataIn_bits_86),
    .io_dataIn_bits_87(muxLyr_io_dataIn_bits_87),
    .io_dataIn_bits_88(muxLyr_io_dataIn_bits_88),
    .io_dataIn_bits_89(muxLyr_io_dataIn_bits_89),
    .io_dataIn_bits_90(muxLyr_io_dataIn_bits_90),
    .io_dataIn_bits_91(muxLyr_io_dataIn_bits_91),
    .io_dataIn_bits_92(muxLyr_io_dataIn_bits_92),
    .io_dataIn_bits_93(muxLyr_io_dataIn_bits_93),
    .io_dataIn_bits_94(muxLyr_io_dataIn_bits_94),
    .io_dataIn_bits_95(muxLyr_io_dataIn_bits_95),
    .io_dataIn_bits_96(muxLyr_io_dataIn_bits_96),
    .io_dataIn_bits_97(muxLyr_io_dataIn_bits_97),
    .io_dataIn_bits_98(muxLyr_io_dataIn_bits_98),
    .io_dataIn_bits_99(muxLyr_io_dataIn_bits_99),
    .io_dataIn_bits_100(muxLyr_io_dataIn_bits_100),
    .io_dataIn_bits_101(muxLyr_io_dataIn_bits_101),
    .io_dataIn_bits_102(muxLyr_io_dataIn_bits_102),
    .io_dataIn_bits_103(muxLyr_io_dataIn_bits_103),
    .io_dataIn_bits_104(muxLyr_io_dataIn_bits_104),
    .io_dataIn_bits_105(muxLyr_io_dataIn_bits_105),
    .io_dataIn_bits_106(muxLyr_io_dataIn_bits_106),
    .io_dataIn_bits_107(muxLyr_io_dataIn_bits_107),
    .io_dataIn_bits_108(muxLyr_io_dataIn_bits_108),
    .io_dataIn_bits_109(muxLyr_io_dataIn_bits_109),
    .io_dataIn_bits_110(muxLyr_io_dataIn_bits_110),
    .io_dataIn_bits_111(muxLyr_io_dataIn_bits_111),
    .io_dataIn_bits_112(muxLyr_io_dataIn_bits_112),
    .io_dataIn_bits_113(muxLyr_io_dataIn_bits_113),
    .io_dataIn_bits_114(muxLyr_io_dataIn_bits_114),
    .io_dataIn_bits_115(muxLyr_io_dataIn_bits_115),
    .io_dataIn_bits_116(muxLyr_io_dataIn_bits_116),
    .io_dataIn_bits_117(muxLyr_io_dataIn_bits_117),
    .io_dataIn_bits_118(muxLyr_io_dataIn_bits_118),
    .io_dataIn_bits_119(muxLyr_io_dataIn_bits_119),
    .io_dataIn_bits_120(muxLyr_io_dataIn_bits_120),
    .io_dataIn_bits_121(muxLyr_io_dataIn_bits_121),
    .io_dataIn_bits_122(muxLyr_io_dataIn_bits_122),
    .io_dataIn_bits_123(muxLyr_io_dataIn_bits_123),
    .io_dataIn_bits_124(muxLyr_io_dataIn_bits_124),
    .io_dataIn_bits_125(muxLyr_io_dataIn_bits_125),
    .io_dataIn_bits_126(muxLyr_io_dataIn_bits_126),
    .io_dataIn_bits_127(muxLyr_io_dataIn_bits_127),
    .io_dataIn_bits_128(muxLyr_io_dataIn_bits_128),
    .io_dataIn_bits_129(muxLyr_io_dataIn_bits_129),
    .io_dataIn_bits_130(muxLyr_io_dataIn_bits_130),
    .io_dataIn_bits_131(muxLyr_io_dataIn_bits_131),
    .io_dataIn_bits_132(muxLyr_io_dataIn_bits_132),
    .io_dataIn_bits_133(muxLyr_io_dataIn_bits_133),
    .io_dataIn_bits_134(muxLyr_io_dataIn_bits_134),
    .io_dataIn_bits_135(muxLyr_io_dataIn_bits_135),
    .io_dataIn_bits_136(muxLyr_io_dataIn_bits_136),
    .io_dataIn_bits_137(muxLyr_io_dataIn_bits_137),
    .io_dataIn_bits_138(muxLyr_io_dataIn_bits_138),
    .io_dataIn_bits_139(muxLyr_io_dataIn_bits_139),
    .io_dataIn_bits_140(muxLyr_io_dataIn_bits_140),
    .io_dataIn_bits_141(muxLyr_io_dataIn_bits_141),
    .io_dataIn_bits_142(muxLyr_io_dataIn_bits_142),
    .io_dataIn_bits_143(muxLyr_io_dataIn_bits_143),
    .io_dataIn_bits_144(muxLyr_io_dataIn_bits_144),
    .io_dataIn_bits_145(muxLyr_io_dataIn_bits_145),
    .io_dataIn_bits_146(muxLyr_io_dataIn_bits_146),
    .io_dataIn_bits_147(muxLyr_io_dataIn_bits_147),
    .io_dataIn_bits_148(muxLyr_io_dataIn_bits_148),
    .io_dataIn_bits_149(muxLyr_io_dataIn_bits_149),
    .io_dataIn_bits_150(muxLyr_io_dataIn_bits_150),
    .io_dataIn_bits_151(muxLyr_io_dataIn_bits_151),
    .io_dataIn_bits_152(muxLyr_io_dataIn_bits_152),
    .io_dataIn_bits_153(muxLyr_io_dataIn_bits_153),
    .io_dataIn_bits_154(muxLyr_io_dataIn_bits_154),
    .io_dataIn_bits_155(muxLyr_io_dataIn_bits_155),
    .io_dataIn_bits_156(muxLyr_io_dataIn_bits_156),
    .io_dataIn_bits_157(muxLyr_io_dataIn_bits_157),
    .io_dataIn_bits_158(muxLyr_io_dataIn_bits_158),
    .io_dataIn_bits_159(muxLyr_io_dataIn_bits_159),
    .io_dataIn_bits_160(muxLyr_io_dataIn_bits_160),
    .io_dataIn_bits_161(muxLyr_io_dataIn_bits_161),
    .io_dataIn_bits_162(muxLyr_io_dataIn_bits_162),
    .io_dataIn_bits_163(muxLyr_io_dataIn_bits_163),
    .io_dataIn_bits_164(muxLyr_io_dataIn_bits_164),
    .io_dataIn_bits_165(muxLyr_io_dataIn_bits_165),
    .io_dataIn_bits_166(muxLyr_io_dataIn_bits_166),
    .io_dataIn_bits_167(muxLyr_io_dataIn_bits_167),
    .io_dataIn_bits_168(muxLyr_io_dataIn_bits_168),
    .io_dataIn_bits_169(muxLyr_io_dataIn_bits_169),
    .io_dataIn_bits_170(muxLyr_io_dataIn_bits_170),
    .io_dataIn_bits_171(muxLyr_io_dataIn_bits_171),
    .io_dataIn_bits_172(muxLyr_io_dataIn_bits_172),
    .io_dataIn_bits_173(muxLyr_io_dataIn_bits_173),
    .io_dataIn_bits_174(muxLyr_io_dataIn_bits_174),
    .io_dataIn_bits_175(muxLyr_io_dataIn_bits_175),
    .io_dataIn_bits_176(muxLyr_io_dataIn_bits_176),
    .io_dataIn_bits_177(muxLyr_io_dataIn_bits_177),
    .io_dataIn_bits_178(muxLyr_io_dataIn_bits_178),
    .io_dataIn_bits_179(muxLyr_io_dataIn_bits_179),
    .io_dataIn_bits_180(muxLyr_io_dataIn_bits_180),
    .io_dataIn_bits_181(muxLyr_io_dataIn_bits_181),
    .io_dataIn_bits_182(muxLyr_io_dataIn_bits_182),
    .io_dataIn_bits_183(muxLyr_io_dataIn_bits_183),
    .io_dataIn_bits_184(muxLyr_io_dataIn_bits_184),
    .io_dataIn_bits_185(muxLyr_io_dataIn_bits_185),
    .io_dataIn_bits_186(muxLyr_io_dataIn_bits_186),
    .io_dataIn_bits_187(muxLyr_io_dataIn_bits_187),
    .io_dataIn_bits_188(muxLyr_io_dataIn_bits_188),
    .io_dataIn_bits_189(muxLyr_io_dataIn_bits_189),
    .io_dataIn_bits_190(muxLyr_io_dataIn_bits_190),
    .io_dataIn_bits_191(muxLyr_io_dataIn_bits_191),
    .io_dataIn_bits_192(muxLyr_io_dataIn_bits_192),
    .io_dataIn_bits_193(muxLyr_io_dataIn_bits_193),
    .io_dataIn_bits_194(muxLyr_io_dataIn_bits_194),
    .io_dataIn_bits_195(muxLyr_io_dataIn_bits_195),
    .io_dataIn_bits_196(muxLyr_io_dataIn_bits_196),
    .io_dataIn_bits_197(muxLyr_io_dataIn_bits_197),
    .io_dataIn_bits_198(muxLyr_io_dataIn_bits_198),
    .io_dataIn_bits_199(muxLyr_io_dataIn_bits_199),
    .io_dataIn_bits_200(muxLyr_io_dataIn_bits_200),
    .io_dataIn_bits_201(muxLyr_io_dataIn_bits_201),
    .io_dataIn_bits_202(muxLyr_io_dataIn_bits_202),
    .io_dataIn_bits_203(muxLyr_io_dataIn_bits_203),
    .io_dataIn_bits_204(muxLyr_io_dataIn_bits_204),
    .io_dataIn_bits_205(muxLyr_io_dataIn_bits_205),
    .io_dataIn_bits_206(muxLyr_io_dataIn_bits_206),
    .io_dataIn_bits_207(muxLyr_io_dataIn_bits_207),
    .io_dataIn_bits_208(muxLyr_io_dataIn_bits_208),
    .io_dataIn_bits_209(muxLyr_io_dataIn_bits_209),
    .io_dataIn_bits_210(muxLyr_io_dataIn_bits_210),
    .io_dataIn_bits_211(muxLyr_io_dataIn_bits_211),
    .io_dataIn_bits_212(muxLyr_io_dataIn_bits_212),
    .io_dataIn_bits_213(muxLyr_io_dataIn_bits_213),
    .io_dataIn_bits_214(muxLyr_io_dataIn_bits_214),
    .io_dataIn_bits_215(muxLyr_io_dataIn_bits_215),
    .io_dataIn_bits_216(muxLyr_io_dataIn_bits_216),
    .io_dataIn_bits_217(muxLyr_io_dataIn_bits_217),
    .io_dataIn_bits_218(muxLyr_io_dataIn_bits_218),
    .io_dataIn_bits_219(muxLyr_io_dataIn_bits_219),
    .io_dataIn_bits_220(muxLyr_io_dataIn_bits_220),
    .io_dataIn_bits_221(muxLyr_io_dataIn_bits_221),
    .io_dataIn_bits_222(muxLyr_io_dataIn_bits_222),
    .io_dataIn_bits_223(muxLyr_io_dataIn_bits_223),
    .io_dataIn_bits_224(muxLyr_io_dataIn_bits_224),
    .io_dataIn_bits_225(muxLyr_io_dataIn_bits_225),
    .io_dataIn_bits_226(muxLyr_io_dataIn_bits_226),
    .io_dataIn_bits_227(muxLyr_io_dataIn_bits_227),
    .io_dataIn_bits_228(muxLyr_io_dataIn_bits_228),
    .io_dataIn_bits_229(muxLyr_io_dataIn_bits_229),
    .io_dataIn_bits_230(muxLyr_io_dataIn_bits_230),
    .io_dataIn_bits_231(muxLyr_io_dataIn_bits_231),
    .io_dataIn_bits_232(muxLyr_io_dataIn_bits_232),
    .io_dataIn_bits_233(muxLyr_io_dataIn_bits_233),
    .io_dataIn_bits_234(muxLyr_io_dataIn_bits_234),
    .io_dataIn_bits_235(muxLyr_io_dataIn_bits_235),
    .io_dataIn_bits_236(muxLyr_io_dataIn_bits_236),
    .io_dataIn_bits_237(muxLyr_io_dataIn_bits_237),
    .io_dataIn_bits_238(muxLyr_io_dataIn_bits_238),
    .io_dataIn_bits_239(muxLyr_io_dataIn_bits_239),
    .io_dataIn_bits_240(muxLyr_io_dataIn_bits_240),
    .io_dataIn_bits_241(muxLyr_io_dataIn_bits_241),
    .io_dataIn_bits_242(muxLyr_io_dataIn_bits_242),
    .io_dataIn_bits_243(muxLyr_io_dataIn_bits_243),
    .io_dataIn_bits_244(muxLyr_io_dataIn_bits_244),
    .io_dataIn_bits_245(muxLyr_io_dataIn_bits_245),
    .io_dataIn_bits_246(muxLyr_io_dataIn_bits_246),
    .io_dataIn_bits_247(muxLyr_io_dataIn_bits_247),
    .io_dataIn_bits_248(muxLyr_io_dataIn_bits_248),
    .io_dataIn_bits_249(muxLyr_io_dataIn_bits_249),
    .io_dataIn_bits_250(muxLyr_io_dataIn_bits_250),
    .io_dataIn_bits_251(muxLyr_io_dataIn_bits_251),
    .io_dataIn_bits_252(muxLyr_io_dataIn_bits_252),
    .io_dataIn_bits_253(muxLyr_io_dataIn_bits_253),
    .io_dataIn_bits_254(muxLyr_io_dataIn_bits_254),
    .io_dataIn_bits_255(muxLyr_io_dataIn_bits_255),
    .io_dataOut_valid(muxLyr_io_dataOut_valid),
    .io_dataOut_bits_0(muxLyr_io_dataOut_bits_0),
    .io_dataOut_bits_1(muxLyr_io_dataOut_bits_1),
    .io_dataOut_bits_2(muxLyr_io_dataOut_bits_2),
    .io_dataOut_bits_3(muxLyr_io_dataOut_bits_3)
  );
  assign _T_29 = $unsigned(vgg_io_dataOut_bits_0); // @[AWSVggWrapper.scala 52:79]
  assign _T_30 = $unsigned(vgg_io_dataOut_bits_1); // @[AWSVggWrapper.scala 52:79]
  assign _T_31 = $unsigned(vgg_io_dataOut_bits_2); // @[AWSVggWrapper.scala 52:79]
  assign _T_32 = $unsigned(vgg_io_dataOut_bits_3); // @[AWSVggWrapper.scala 52:79]
  assign _T_33 = $unsigned(vgg_io_dataOut_bits_4); // @[AWSVggWrapper.scala 52:79]
  assign _T_34 = $unsigned(vgg_io_dataOut_bits_5); // @[AWSVggWrapper.scala 52:79]
  assign _T_35 = $unsigned(vgg_io_dataOut_bits_6); // @[AWSVggWrapper.scala 52:79]
  assign _T_36 = $unsigned(vgg_io_dataOut_bits_7); // @[AWSVggWrapper.scala 52:79]
  assign _T_37 = $unsigned(vgg_io_dataOut_bits_8); // @[AWSVggWrapper.scala 52:79]
  assign _T_38 = $unsigned(vgg_io_dataOut_bits_9); // @[AWSVggWrapper.scala 52:79]
  assign _T_39 = $unsigned(vgg_io_dataOut_bits_10); // @[AWSVggWrapper.scala 52:79]
  assign _T_40 = $unsigned(vgg_io_dataOut_bits_11); // @[AWSVggWrapper.scala 52:79]
  assign _T_41 = $unsigned(vgg_io_dataOut_bits_12); // @[AWSVggWrapper.scala 52:79]
  assign _T_42 = $unsigned(vgg_io_dataOut_bits_13); // @[AWSVggWrapper.scala 52:79]
  assign _T_43 = $unsigned(vgg_io_dataOut_bits_14); // @[AWSVggWrapper.scala 52:79]
  assign _T_44 = $unsigned(vgg_io_dataOut_bits_15); // @[AWSVggWrapper.scala 52:79]
  assign _T_45 = $unsigned(vgg_io_dataOut_bits_16); // @[AWSVggWrapper.scala 52:79]
  assign _T_46 = $unsigned(vgg_io_dataOut_bits_17); // @[AWSVggWrapper.scala 52:79]
  assign _T_47 = $unsigned(vgg_io_dataOut_bits_18); // @[AWSVggWrapper.scala 52:79]
  assign _T_48 = $unsigned(vgg_io_dataOut_bits_19); // @[AWSVggWrapper.scala 52:79]
  assign _T_49 = $unsigned(vgg_io_dataOut_bits_20); // @[AWSVggWrapper.scala 52:79]
  assign _T_50 = $unsigned(vgg_io_dataOut_bits_21); // @[AWSVggWrapper.scala 52:79]
  assign _T_51 = $unsigned(vgg_io_dataOut_bits_22); // @[AWSVggWrapper.scala 52:79]
  assign _T_52 = $unsigned(vgg_io_dataOut_bits_23); // @[AWSVggWrapper.scala 52:79]
  assign _T_53 = $unsigned(vgg_io_dataOut_bits_24); // @[AWSVggWrapper.scala 52:79]
  assign _T_54 = $unsigned(vgg_io_dataOut_bits_25); // @[AWSVggWrapper.scala 52:79]
  assign _T_55 = $unsigned(vgg_io_dataOut_bits_26); // @[AWSVggWrapper.scala 52:79]
  assign _T_56 = $unsigned(vgg_io_dataOut_bits_27); // @[AWSVggWrapper.scala 52:79]
  assign _T_57 = $unsigned(vgg_io_dataOut_bits_28); // @[AWSVggWrapper.scala 52:79]
  assign _T_58 = $unsigned(vgg_io_dataOut_bits_29); // @[AWSVggWrapper.scala 52:79]
  assign _T_59 = $unsigned(vgg_io_dataOut_bits_30); // @[AWSVggWrapper.scala 52:79]
  assign _T_60 = $unsigned(vgg_io_dataOut_bits_31); // @[AWSVggWrapper.scala 52:79]
  assign _T_61 = $unsigned(vgg_io_dataOut_bits_32); // @[AWSVggWrapper.scala 52:79]
  assign _T_62 = $unsigned(vgg_io_dataOut_bits_33); // @[AWSVggWrapper.scala 52:79]
  assign _T_63 = $unsigned(vgg_io_dataOut_bits_34); // @[AWSVggWrapper.scala 52:79]
  assign _T_64 = $unsigned(vgg_io_dataOut_bits_35); // @[AWSVggWrapper.scala 52:79]
  assign _T_65 = $unsigned(vgg_io_dataOut_bits_36); // @[AWSVggWrapper.scala 52:79]
  assign _T_66 = $unsigned(vgg_io_dataOut_bits_37); // @[AWSVggWrapper.scala 52:79]
  assign _T_67 = $unsigned(vgg_io_dataOut_bits_38); // @[AWSVggWrapper.scala 52:79]
  assign _T_68 = $unsigned(vgg_io_dataOut_bits_39); // @[AWSVggWrapper.scala 52:79]
  assign _T_69 = $unsigned(vgg_io_dataOut_bits_40); // @[AWSVggWrapper.scala 52:79]
  assign _T_70 = $unsigned(vgg_io_dataOut_bits_41); // @[AWSVggWrapper.scala 52:79]
  assign _T_71 = $unsigned(vgg_io_dataOut_bits_42); // @[AWSVggWrapper.scala 52:79]
  assign _T_72 = $unsigned(vgg_io_dataOut_bits_43); // @[AWSVggWrapper.scala 52:79]
  assign _T_73 = $unsigned(vgg_io_dataOut_bits_44); // @[AWSVggWrapper.scala 52:79]
  assign _T_74 = $unsigned(vgg_io_dataOut_bits_45); // @[AWSVggWrapper.scala 52:79]
  assign _T_75 = $unsigned(vgg_io_dataOut_bits_46); // @[AWSVggWrapper.scala 52:79]
  assign _T_76 = $unsigned(vgg_io_dataOut_bits_47); // @[AWSVggWrapper.scala 52:79]
  assign _T_77 = $unsigned(vgg_io_dataOut_bits_48); // @[AWSVggWrapper.scala 52:79]
  assign _T_78 = $unsigned(vgg_io_dataOut_bits_49); // @[AWSVggWrapper.scala 52:79]
  assign _T_79 = $unsigned(vgg_io_dataOut_bits_50); // @[AWSVggWrapper.scala 52:79]
  assign _T_80 = $unsigned(vgg_io_dataOut_bits_51); // @[AWSVggWrapper.scala 52:79]
  assign _T_81 = $unsigned(vgg_io_dataOut_bits_52); // @[AWSVggWrapper.scala 52:79]
  assign _T_82 = $unsigned(vgg_io_dataOut_bits_53); // @[AWSVggWrapper.scala 52:79]
  assign _T_83 = $unsigned(vgg_io_dataOut_bits_54); // @[AWSVggWrapper.scala 52:79]
  assign _T_84 = $unsigned(vgg_io_dataOut_bits_55); // @[AWSVggWrapper.scala 52:79]
  assign _T_85 = $unsigned(vgg_io_dataOut_bits_56); // @[AWSVggWrapper.scala 52:79]
  assign _T_86 = $unsigned(vgg_io_dataOut_bits_57); // @[AWSVggWrapper.scala 52:79]
  assign _T_87 = $unsigned(vgg_io_dataOut_bits_58); // @[AWSVggWrapper.scala 52:79]
  assign _T_88 = $unsigned(vgg_io_dataOut_bits_59); // @[AWSVggWrapper.scala 52:79]
  assign _T_89 = $unsigned(vgg_io_dataOut_bits_60); // @[AWSVggWrapper.scala 52:79]
  assign _T_90 = $unsigned(vgg_io_dataOut_bits_61); // @[AWSVggWrapper.scala 52:79]
  assign _T_91 = $unsigned(vgg_io_dataOut_bits_62); // @[AWSVggWrapper.scala 52:79]
  assign _T_92 = $unsigned(vgg_io_dataOut_bits_63); // @[AWSVggWrapper.scala 52:79]
  assign _T_93 = $unsigned(vgg_io_dataOut_bits_64); // @[AWSVggWrapper.scala 52:79]
  assign _T_94 = $unsigned(vgg_io_dataOut_bits_65); // @[AWSVggWrapper.scala 52:79]
  assign _T_95 = $unsigned(vgg_io_dataOut_bits_66); // @[AWSVggWrapper.scala 52:79]
  assign _T_96 = $unsigned(vgg_io_dataOut_bits_67); // @[AWSVggWrapper.scala 52:79]
  assign _T_97 = $unsigned(vgg_io_dataOut_bits_68); // @[AWSVggWrapper.scala 52:79]
  assign _T_98 = $unsigned(vgg_io_dataOut_bits_69); // @[AWSVggWrapper.scala 52:79]
  assign _T_99 = $unsigned(vgg_io_dataOut_bits_70); // @[AWSVggWrapper.scala 52:79]
  assign _T_100 = $unsigned(vgg_io_dataOut_bits_71); // @[AWSVggWrapper.scala 52:79]
  assign _T_101 = $unsigned(vgg_io_dataOut_bits_72); // @[AWSVggWrapper.scala 52:79]
  assign _T_102 = $unsigned(vgg_io_dataOut_bits_73); // @[AWSVggWrapper.scala 52:79]
  assign _T_103 = $unsigned(vgg_io_dataOut_bits_74); // @[AWSVggWrapper.scala 52:79]
  assign _T_104 = $unsigned(vgg_io_dataOut_bits_75); // @[AWSVggWrapper.scala 52:79]
  assign _T_105 = $unsigned(vgg_io_dataOut_bits_76); // @[AWSVggWrapper.scala 52:79]
  assign _T_106 = $unsigned(vgg_io_dataOut_bits_77); // @[AWSVggWrapper.scala 52:79]
  assign _T_107 = $unsigned(vgg_io_dataOut_bits_78); // @[AWSVggWrapper.scala 52:79]
  assign _T_108 = $unsigned(vgg_io_dataOut_bits_79); // @[AWSVggWrapper.scala 52:79]
  assign _T_109 = $unsigned(vgg_io_dataOut_bits_80); // @[AWSVggWrapper.scala 52:79]
  assign _T_110 = $unsigned(vgg_io_dataOut_bits_81); // @[AWSVggWrapper.scala 52:79]
  assign _T_111 = $unsigned(vgg_io_dataOut_bits_82); // @[AWSVggWrapper.scala 52:79]
  assign _T_112 = $unsigned(vgg_io_dataOut_bits_83); // @[AWSVggWrapper.scala 52:79]
  assign _T_113 = $unsigned(vgg_io_dataOut_bits_84); // @[AWSVggWrapper.scala 52:79]
  assign _T_114 = $unsigned(vgg_io_dataOut_bits_85); // @[AWSVggWrapper.scala 52:79]
  assign _T_115 = $unsigned(vgg_io_dataOut_bits_86); // @[AWSVggWrapper.scala 52:79]
  assign _T_116 = $unsigned(vgg_io_dataOut_bits_87); // @[AWSVggWrapper.scala 52:79]
  assign _T_117 = $unsigned(vgg_io_dataOut_bits_88); // @[AWSVggWrapper.scala 52:79]
  assign _T_118 = $unsigned(vgg_io_dataOut_bits_89); // @[AWSVggWrapper.scala 52:79]
  assign _T_119 = $unsigned(vgg_io_dataOut_bits_90); // @[AWSVggWrapper.scala 52:79]
  assign _T_120 = $unsigned(vgg_io_dataOut_bits_91); // @[AWSVggWrapper.scala 52:79]
  assign _T_121 = $unsigned(vgg_io_dataOut_bits_92); // @[AWSVggWrapper.scala 52:79]
  assign _T_122 = $unsigned(vgg_io_dataOut_bits_93); // @[AWSVggWrapper.scala 52:79]
  assign _T_123 = $unsigned(vgg_io_dataOut_bits_94); // @[AWSVggWrapper.scala 52:79]
  assign _T_124 = $unsigned(vgg_io_dataOut_bits_95); // @[AWSVggWrapper.scala 52:79]
  assign _T_125 = $unsigned(vgg_io_dataOut_bits_96); // @[AWSVggWrapper.scala 52:79]
  assign _T_126 = $unsigned(vgg_io_dataOut_bits_97); // @[AWSVggWrapper.scala 52:79]
  assign _T_127 = $unsigned(vgg_io_dataOut_bits_98); // @[AWSVggWrapper.scala 52:79]
  assign _T_128 = $unsigned(vgg_io_dataOut_bits_99); // @[AWSVggWrapper.scala 52:79]
  assign _T_129 = $unsigned(vgg_io_dataOut_bits_100); // @[AWSVggWrapper.scala 52:79]
  assign _T_130 = $unsigned(vgg_io_dataOut_bits_101); // @[AWSVggWrapper.scala 52:79]
  assign _T_131 = $unsigned(vgg_io_dataOut_bits_102); // @[AWSVggWrapper.scala 52:79]
  assign _T_132 = $unsigned(vgg_io_dataOut_bits_103); // @[AWSVggWrapper.scala 52:79]
  assign _T_133 = $unsigned(vgg_io_dataOut_bits_104); // @[AWSVggWrapper.scala 52:79]
  assign _T_134 = $unsigned(vgg_io_dataOut_bits_105); // @[AWSVggWrapper.scala 52:79]
  assign _T_135 = $unsigned(vgg_io_dataOut_bits_106); // @[AWSVggWrapper.scala 52:79]
  assign _T_136 = $unsigned(vgg_io_dataOut_bits_107); // @[AWSVggWrapper.scala 52:79]
  assign _T_137 = $unsigned(vgg_io_dataOut_bits_108); // @[AWSVggWrapper.scala 52:79]
  assign _T_138 = $unsigned(vgg_io_dataOut_bits_109); // @[AWSVggWrapper.scala 52:79]
  assign _T_139 = $unsigned(vgg_io_dataOut_bits_110); // @[AWSVggWrapper.scala 52:79]
  assign _T_140 = $unsigned(vgg_io_dataOut_bits_111); // @[AWSVggWrapper.scala 52:79]
  assign _T_141 = $unsigned(vgg_io_dataOut_bits_112); // @[AWSVggWrapper.scala 52:79]
  assign _T_142 = $unsigned(vgg_io_dataOut_bits_113); // @[AWSVggWrapper.scala 52:79]
  assign _T_143 = $unsigned(vgg_io_dataOut_bits_114); // @[AWSVggWrapper.scala 52:79]
  assign _T_144 = $unsigned(vgg_io_dataOut_bits_115); // @[AWSVggWrapper.scala 52:79]
  assign _T_145 = $unsigned(vgg_io_dataOut_bits_116); // @[AWSVggWrapper.scala 52:79]
  assign _T_146 = $unsigned(vgg_io_dataOut_bits_117); // @[AWSVggWrapper.scala 52:79]
  assign _T_147 = $unsigned(vgg_io_dataOut_bits_118); // @[AWSVggWrapper.scala 52:79]
  assign _T_148 = $unsigned(vgg_io_dataOut_bits_119); // @[AWSVggWrapper.scala 52:79]
  assign _T_149 = $unsigned(vgg_io_dataOut_bits_120); // @[AWSVggWrapper.scala 52:79]
  assign _T_150 = $unsigned(vgg_io_dataOut_bits_121); // @[AWSVggWrapper.scala 52:79]
  assign _T_151 = $unsigned(vgg_io_dataOut_bits_122); // @[AWSVggWrapper.scala 52:79]
  assign _T_152 = $unsigned(vgg_io_dataOut_bits_123); // @[AWSVggWrapper.scala 52:79]
  assign _T_153 = $unsigned(vgg_io_dataOut_bits_124); // @[AWSVggWrapper.scala 52:79]
  assign _T_154 = $unsigned(vgg_io_dataOut_bits_125); // @[AWSVggWrapper.scala 52:79]
  assign _T_155 = $unsigned(vgg_io_dataOut_bits_126); // @[AWSVggWrapper.scala 52:79]
  assign _T_156 = $unsigned(vgg_io_dataOut_bits_127); // @[AWSVggWrapper.scala 52:79]
  assign _T_157 = $unsigned(vgg_io_dataOut_bits_128); // @[AWSVggWrapper.scala 52:79]
  assign _T_158 = $unsigned(vgg_io_dataOut_bits_129); // @[AWSVggWrapper.scala 52:79]
  assign _T_159 = $unsigned(vgg_io_dataOut_bits_130); // @[AWSVggWrapper.scala 52:79]
  assign _T_160 = $unsigned(vgg_io_dataOut_bits_131); // @[AWSVggWrapper.scala 52:79]
  assign _T_161 = $unsigned(vgg_io_dataOut_bits_132); // @[AWSVggWrapper.scala 52:79]
  assign _T_162 = $unsigned(vgg_io_dataOut_bits_133); // @[AWSVggWrapper.scala 52:79]
  assign _T_163 = $unsigned(vgg_io_dataOut_bits_134); // @[AWSVggWrapper.scala 52:79]
  assign _T_164 = $unsigned(vgg_io_dataOut_bits_135); // @[AWSVggWrapper.scala 52:79]
  assign _T_165 = $unsigned(vgg_io_dataOut_bits_136); // @[AWSVggWrapper.scala 52:79]
  assign _T_166 = $unsigned(vgg_io_dataOut_bits_137); // @[AWSVggWrapper.scala 52:79]
  assign _T_167 = $unsigned(vgg_io_dataOut_bits_138); // @[AWSVggWrapper.scala 52:79]
  assign _T_168 = $unsigned(vgg_io_dataOut_bits_139); // @[AWSVggWrapper.scala 52:79]
  assign _T_169 = $unsigned(vgg_io_dataOut_bits_140); // @[AWSVggWrapper.scala 52:79]
  assign _T_170 = $unsigned(vgg_io_dataOut_bits_141); // @[AWSVggWrapper.scala 52:79]
  assign _T_171 = $unsigned(vgg_io_dataOut_bits_142); // @[AWSVggWrapper.scala 52:79]
  assign _T_172 = $unsigned(vgg_io_dataOut_bits_143); // @[AWSVggWrapper.scala 52:79]
  assign _T_173 = $unsigned(vgg_io_dataOut_bits_144); // @[AWSVggWrapper.scala 52:79]
  assign _T_174 = $unsigned(vgg_io_dataOut_bits_145); // @[AWSVggWrapper.scala 52:79]
  assign _T_175 = $unsigned(vgg_io_dataOut_bits_146); // @[AWSVggWrapper.scala 52:79]
  assign _T_176 = $unsigned(vgg_io_dataOut_bits_147); // @[AWSVggWrapper.scala 52:79]
  assign _T_177 = $unsigned(vgg_io_dataOut_bits_148); // @[AWSVggWrapper.scala 52:79]
  assign _T_178 = $unsigned(vgg_io_dataOut_bits_149); // @[AWSVggWrapper.scala 52:79]
  assign _T_179 = $unsigned(vgg_io_dataOut_bits_150); // @[AWSVggWrapper.scala 52:79]
  assign _T_180 = $unsigned(vgg_io_dataOut_bits_151); // @[AWSVggWrapper.scala 52:79]
  assign _T_181 = $unsigned(vgg_io_dataOut_bits_152); // @[AWSVggWrapper.scala 52:79]
  assign _T_182 = $unsigned(vgg_io_dataOut_bits_153); // @[AWSVggWrapper.scala 52:79]
  assign _T_183 = $unsigned(vgg_io_dataOut_bits_154); // @[AWSVggWrapper.scala 52:79]
  assign _T_184 = $unsigned(vgg_io_dataOut_bits_155); // @[AWSVggWrapper.scala 52:79]
  assign _T_185 = $unsigned(vgg_io_dataOut_bits_156); // @[AWSVggWrapper.scala 52:79]
  assign _T_186 = $unsigned(vgg_io_dataOut_bits_157); // @[AWSVggWrapper.scala 52:79]
  assign _T_187 = $unsigned(vgg_io_dataOut_bits_158); // @[AWSVggWrapper.scala 52:79]
  assign _T_188 = $unsigned(vgg_io_dataOut_bits_159); // @[AWSVggWrapper.scala 52:79]
  assign _T_189 = $unsigned(vgg_io_dataOut_bits_160); // @[AWSVggWrapper.scala 52:79]
  assign _T_190 = $unsigned(vgg_io_dataOut_bits_161); // @[AWSVggWrapper.scala 52:79]
  assign _T_191 = $unsigned(vgg_io_dataOut_bits_162); // @[AWSVggWrapper.scala 52:79]
  assign _T_192 = $unsigned(vgg_io_dataOut_bits_163); // @[AWSVggWrapper.scala 52:79]
  assign _T_193 = $unsigned(vgg_io_dataOut_bits_164); // @[AWSVggWrapper.scala 52:79]
  assign _T_194 = $unsigned(vgg_io_dataOut_bits_165); // @[AWSVggWrapper.scala 52:79]
  assign _T_195 = $unsigned(vgg_io_dataOut_bits_166); // @[AWSVggWrapper.scala 52:79]
  assign _T_196 = $unsigned(vgg_io_dataOut_bits_167); // @[AWSVggWrapper.scala 52:79]
  assign _T_197 = $unsigned(vgg_io_dataOut_bits_168); // @[AWSVggWrapper.scala 52:79]
  assign _T_198 = $unsigned(vgg_io_dataOut_bits_169); // @[AWSVggWrapper.scala 52:79]
  assign _T_199 = $unsigned(vgg_io_dataOut_bits_170); // @[AWSVggWrapper.scala 52:79]
  assign _T_200 = $unsigned(vgg_io_dataOut_bits_171); // @[AWSVggWrapper.scala 52:79]
  assign _T_201 = $unsigned(vgg_io_dataOut_bits_172); // @[AWSVggWrapper.scala 52:79]
  assign _T_202 = $unsigned(vgg_io_dataOut_bits_173); // @[AWSVggWrapper.scala 52:79]
  assign _T_203 = $unsigned(vgg_io_dataOut_bits_174); // @[AWSVggWrapper.scala 52:79]
  assign _T_204 = $unsigned(vgg_io_dataOut_bits_175); // @[AWSVggWrapper.scala 52:79]
  assign _T_205 = $unsigned(vgg_io_dataOut_bits_176); // @[AWSVggWrapper.scala 52:79]
  assign _T_206 = $unsigned(vgg_io_dataOut_bits_177); // @[AWSVggWrapper.scala 52:79]
  assign _T_207 = $unsigned(vgg_io_dataOut_bits_178); // @[AWSVggWrapper.scala 52:79]
  assign _T_208 = $unsigned(vgg_io_dataOut_bits_179); // @[AWSVggWrapper.scala 52:79]
  assign _T_209 = $unsigned(vgg_io_dataOut_bits_180); // @[AWSVggWrapper.scala 52:79]
  assign _T_210 = $unsigned(vgg_io_dataOut_bits_181); // @[AWSVggWrapper.scala 52:79]
  assign _T_211 = $unsigned(vgg_io_dataOut_bits_182); // @[AWSVggWrapper.scala 52:79]
  assign _T_212 = $unsigned(vgg_io_dataOut_bits_183); // @[AWSVggWrapper.scala 52:79]
  assign _T_213 = $unsigned(vgg_io_dataOut_bits_184); // @[AWSVggWrapper.scala 52:79]
  assign _T_214 = $unsigned(vgg_io_dataOut_bits_185); // @[AWSVggWrapper.scala 52:79]
  assign _T_215 = $unsigned(vgg_io_dataOut_bits_186); // @[AWSVggWrapper.scala 52:79]
  assign _T_216 = $unsigned(vgg_io_dataOut_bits_187); // @[AWSVggWrapper.scala 52:79]
  assign _T_217 = $unsigned(vgg_io_dataOut_bits_188); // @[AWSVggWrapper.scala 52:79]
  assign _T_218 = $unsigned(vgg_io_dataOut_bits_189); // @[AWSVggWrapper.scala 52:79]
  assign _T_219 = $unsigned(vgg_io_dataOut_bits_190); // @[AWSVggWrapper.scala 52:79]
  assign _T_220 = $unsigned(vgg_io_dataOut_bits_191); // @[AWSVggWrapper.scala 52:79]
  assign _T_221 = $unsigned(vgg_io_dataOut_bits_192); // @[AWSVggWrapper.scala 52:79]
  assign _T_222 = $unsigned(vgg_io_dataOut_bits_193); // @[AWSVggWrapper.scala 52:79]
  assign _T_223 = $unsigned(vgg_io_dataOut_bits_194); // @[AWSVggWrapper.scala 52:79]
  assign _T_224 = $unsigned(vgg_io_dataOut_bits_195); // @[AWSVggWrapper.scala 52:79]
  assign _T_225 = $unsigned(vgg_io_dataOut_bits_196); // @[AWSVggWrapper.scala 52:79]
  assign _T_226 = $unsigned(vgg_io_dataOut_bits_197); // @[AWSVggWrapper.scala 52:79]
  assign _T_227 = $unsigned(vgg_io_dataOut_bits_198); // @[AWSVggWrapper.scala 52:79]
  assign _T_228 = $unsigned(vgg_io_dataOut_bits_199); // @[AWSVggWrapper.scala 52:79]
  assign _T_229 = $unsigned(vgg_io_dataOut_bits_200); // @[AWSVggWrapper.scala 52:79]
  assign _T_230 = $unsigned(vgg_io_dataOut_bits_201); // @[AWSVggWrapper.scala 52:79]
  assign _T_231 = $unsigned(vgg_io_dataOut_bits_202); // @[AWSVggWrapper.scala 52:79]
  assign _T_232 = $unsigned(vgg_io_dataOut_bits_203); // @[AWSVggWrapper.scala 52:79]
  assign _T_233 = $unsigned(vgg_io_dataOut_bits_204); // @[AWSVggWrapper.scala 52:79]
  assign _T_234 = $unsigned(vgg_io_dataOut_bits_205); // @[AWSVggWrapper.scala 52:79]
  assign _T_235 = $unsigned(vgg_io_dataOut_bits_206); // @[AWSVggWrapper.scala 52:79]
  assign _T_236 = $unsigned(vgg_io_dataOut_bits_207); // @[AWSVggWrapper.scala 52:79]
  assign _T_237 = $unsigned(vgg_io_dataOut_bits_208); // @[AWSVggWrapper.scala 52:79]
  assign _T_238 = $unsigned(vgg_io_dataOut_bits_209); // @[AWSVggWrapper.scala 52:79]
  assign _T_239 = $unsigned(vgg_io_dataOut_bits_210); // @[AWSVggWrapper.scala 52:79]
  assign _T_240 = $unsigned(vgg_io_dataOut_bits_211); // @[AWSVggWrapper.scala 52:79]
  assign _T_241 = $unsigned(vgg_io_dataOut_bits_212); // @[AWSVggWrapper.scala 52:79]
  assign _T_242 = $unsigned(vgg_io_dataOut_bits_213); // @[AWSVggWrapper.scala 52:79]
  assign _T_243 = $unsigned(vgg_io_dataOut_bits_214); // @[AWSVggWrapper.scala 52:79]
  assign _T_244 = $unsigned(vgg_io_dataOut_bits_215); // @[AWSVggWrapper.scala 52:79]
  assign _T_245 = $unsigned(vgg_io_dataOut_bits_216); // @[AWSVggWrapper.scala 52:79]
  assign _T_246 = $unsigned(vgg_io_dataOut_bits_217); // @[AWSVggWrapper.scala 52:79]
  assign _T_247 = $unsigned(vgg_io_dataOut_bits_218); // @[AWSVggWrapper.scala 52:79]
  assign _T_248 = $unsigned(vgg_io_dataOut_bits_219); // @[AWSVggWrapper.scala 52:79]
  assign _T_249 = $unsigned(vgg_io_dataOut_bits_220); // @[AWSVggWrapper.scala 52:79]
  assign _T_250 = $unsigned(vgg_io_dataOut_bits_221); // @[AWSVggWrapper.scala 52:79]
  assign _T_251 = $unsigned(vgg_io_dataOut_bits_222); // @[AWSVggWrapper.scala 52:79]
  assign _T_252 = $unsigned(vgg_io_dataOut_bits_223); // @[AWSVggWrapper.scala 52:79]
  assign _T_253 = $unsigned(vgg_io_dataOut_bits_224); // @[AWSVggWrapper.scala 52:79]
  assign _T_254 = $unsigned(vgg_io_dataOut_bits_225); // @[AWSVggWrapper.scala 52:79]
  assign _T_255 = $unsigned(vgg_io_dataOut_bits_226); // @[AWSVggWrapper.scala 52:79]
  assign _T_256 = $unsigned(vgg_io_dataOut_bits_227); // @[AWSVggWrapper.scala 52:79]
  assign _T_257 = $unsigned(vgg_io_dataOut_bits_228); // @[AWSVggWrapper.scala 52:79]
  assign _T_258 = $unsigned(vgg_io_dataOut_bits_229); // @[AWSVggWrapper.scala 52:79]
  assign _T_259 = $unsigned(vgg_io_dataOut_bits_230); // @[AWSVggWrapper.scala 52:79]
  assign _T_260 = $unsigned(vgg_io_dataOut_bits_231); // @[AWSVggWrapper.scala 52:79]
  assign _T_261 = $unsigned(vgg_io_dataOut_bits_232); // @[AWSVggWrapper.scala 52:79]
  assign _T_262 = $unsigned(vgg_io_dataOut_bits_233); // @[AWSVggWrapper.scala 52:79]
  assign _T_263 = $unsigned(vgg_io_dataOut_bits_234); // @[AWSVggWrapper.scala 52:79]
  assign _T_264 = $unsigned(vgg_io_dataOut_bits_235); // @[AWSVggWrapper.scala 52:79]
  assign _T_265 = $unsigned(vgg_io_dataOut_bits_236); // @[AWSVggWrapper.scala 52:79]
  assign _T_266 = $unsigned(vgg_io_dataOut_bits_237); // @[AWSVggWrapper.scala 52:79]
  assign _T_267 = $unsigned(vgg_io_dataOut_bits_238); // @[AWSVggWrapper.scala 52:79]
  assign _T_268 = $unsigned(vgg_io_dataOut_bits_239); // @[AWSVggWrapper.scala 52:79]
  assign _T_269 = $unsigned(vgg_io_dataOut_bits_240); // @[AWSVggWrapper.scala 52:79]
  assign _T_270 = $unsigned(vgg_io_dataOut_bits_241); // @[AWSVggWrapper.scala 52:79]
  assign _T_271 = $unsigned(vgg_io_dataOut_bits_242); // @[AWSVggWrapper.scala 52:79]
  assign _T_272 = $unsigned(vgg_io_dataOut_bits_243); // @[AWSVggWrapper.scala 52:79]
  assign _T_273 = $unsigned(vgg_io_dataOut_bits_244); // @[AWSVggWrapper.scala 52:79]
  assign _T_274 = $unsigned(vgg_io_dataOut_bits_245); // @[AWSVggWrapper.scala 52:79]
  assign _T_275 = $unsigned(vgg_io_dataOut_bits_246); // @[AWSVggWrapper.scala 52:79]
  assign _T_276 = $unsigned(vgg_io_dataOut_bits_247); // @[AWSVggWrapper.scala 52:79]
  assign _T_277 = $unsigned(vgg_io_dataOut_bits_248); // @[AWSVggWrapper.scala 52:79]
  assign _T_278 = $unsigned(vgg_io_dataOut_bits_249); // @[AWSVggWrapper.scala 52:79]
  assign _T_279 = $unsigned(vgg_io_dataOut_bits_250); // @[AWSVggWrapper.scala 52:79]
  assign _T_280 = $unsigned(vgg_io_dataOut_bits_251); // @[AWSVggWrapper.scala 52:79]
  assign _T_281 = $unsigned(vgg_io_dataOut_bits_252); // @[AWSVggWrapper.scala 52:79]
  assign _T_282 = $unsigned(vgg_io_dataOut_bits_253); // @[AWSVggWrapper.scala 52:79]
  assign _T_283 = $unsigned(vgg_io_dataOut_bits_254); // @[AWSVggWrapper.scala 52:79]
  assign _T_284 = $unsigned(vgg_io_dataOut_bits_255); // @[AWSVggWrapper.scala 52:79]
  assign _T_285 = {_T_29,_T_30}; // @[AWSVggWrapper.scala 52:94]
  assign _T_286 = {_T_285,_T_31}; // @[AWSVggWrapper.scala 52:94]
  assign _T_287 = {_T_286,_T_32}; // @[AWSVggWrapper.scala 52:94]
  assign _T_288 = {_T_287,_T_33}; // @[AWSVggWrapper.scala 52:94]
  assign _T_289 = {_T_288,_T_34}; // @[AWSVggWrapper.scala 52:94]
  assign _T_290 = {_T_289,_T_35}; // @[AWSVggWrapper.scala 52:94]
  assign _T_291 = {_T_290,_T_36}; // @[AWSVggWrapper.scala 52:94]
  assign _T_292 = {_T_291,_T_37}; // @[AWSVggWrapper.scala 52:94]
  assign _T_293 = {_T_292,_T_38}; // @[AWSVggWrapper.scala 52:94]
  assign _T_294 = {_T_293,_T_39}; // @[AWSVggWrapper.scala 52:94]
  assign _T_295 = {_T_294,_T_40}; // @[AWSVggWrapper.scala 52:94]
  assign _T_296 = {_T_295,_T_41}; // @[AWSVggWrapper.scala 52:94]
  assign _T_297 = {_T_296,_T_42}; // @[AWSVggWrapper.scala 52:94]
  assign _T_298 = {_T_297,_T_43}; // @[AWSVggWrapper.scala 52:94]
  assign _T_299 = {_T_298,_T_44}; // @[AWSVggWrapper.scala 52:94]
  assign _T_300 = {_T_299,_T_45}; // @[AWSVggWrapper.scala 52:94]
  assign _T_301 = {_T_300,_T_46}; // @[AWSVggWrapper.scala 52:94]
  assign _T_302 = {_T_301,_T_47}; // @[AWSVggWrapper.scala 52:94]
  assign _T_303 = {_T_302,_T_48}; // @[AWSVggWrapper.scala 52:94]
  assign _T_304 = {_T_303,_T_49}; // @[AWSVggWrapper.scala 52:94]
  assign _T_305 = {_T_304,_T_50}; // @[AWSVggWrapper.scala 52:94]
  assign _T_306 = {_T_305,_T_51}; // @[AWSVggWrapper.scala 52:94]
  assign _T_307 = {_T_306,_T_52}; // @[AWSVggWrapper.scala 52:94]
  assign _T_308 = {_T_307,_T_53}; // @[AWSVggWrapper.scala 52:94]
  assign _T_309 = {_T_308,_T_54}; // @[AWSVggWrapper.scala 52:94]
  assign _T_310 = {_T_309,_T_55}; // @[AWSVggWrapper.scala 52:94]
  assign _T_311 = {_T_310,_T_56}; // @[AWSVggWrapper.scala 52:94]
  assign _T_312 = {_T_311,_T_57}; // @[AWSVggWrapper.scala 52:94]
  assign _T_313 = {_T_312,_T_58}; // @[AWSVggWrapper.scala 52:94]
  assign _T_314 = {_T_313,_T_59}; // @[AWSVggWrapper.scala 52:94]
  assign _T_315 = {_T_314,_T_60}; // @[AWSVggWrapper.scala 52:94]
  assign _T_316 = {_T_315,_T_61}; // @[AWSVggWrapper.scala 52:94]
  assign _T_317 = {_T_316,_T_62}; // @[AWSVggWrapper.scala 52:94]
  assign _T_318 = {_T_317,_T_63}; // @[AWSVggWrapper.scala 52:94]
  assign _T_319 = {_T_318,_T_64}; // @[AWSVggWrapper.scala 52:94]
  assign _T_320 = {_T_319,_T_65}; // @[AWSVggWrapper.scala 52:94]
  assign _T_321 = {_T_320,_T_66}; // @[AWSVggWrapper.scala 52:94]
  assign _T_322 = {_T_321,_T_67}; // @[AWSVggWrapper.scala 52:94]
  assign _T_323 = {_T_322,_T_68}; // @[AWSVggWrapper.scala 52:94]
  assign _T_324 = {_T_323,_T_69}; // @[AWSVggWrapper.scala 52:94]
  assign _T_325 = {_T_324,_T_70}; // @[AWSVggWrapper.scala 52:94]
  assign _T_326 = {_T_325,_T_71}; // @[AWSVggWrapper.scala 52:94]
  assign _T_327 = {_T_326,_T_72}; // @[AWSVggWrapper.scala 52:94]
  assign _T_328 = {_T_327,_T_73}; // @[AWSVggWrapper.scala 52:94]
  assign _T_329 = {_T_328,_T_74}; // @[AWSVggWrapper.scala 52:94]
  assign _T_330 = {_T_329,_T_75}; // @[AWSVggWrapper.scala 52:94]
  assign _T_331 = {_T_330,_T_76}; // @[AWSVggWrapper.scala 52:94]
  assign _T_332 = {_T_331,_T_77}; // @[AWSVggWrapper.scala 52:94]
  assign _T_333 = {_T_332,_T_78}; // @[AWSVggWrapper.scala 52:94]
  assign _T_334 = {_T_333,_T_79}; // @[AWSVggWrapper.scala 52:94]
  assign _T_335 = {_T_334,_T_80}; // @[AWSVggWrapper.scala 52:94]
  assign _T_336 = {_T_335,_T_81}; // @[AWSVggWrapper.scala 52:94]
  assign _T_337 = {_T_336,_T_82}; // @[AWSVggWrapper.scala 52:94]
  assign _T_338 = {_T_337,_T_83}; // @[AWSVggWrapper.scala 52:94]
  assign _T_339 = {_T_338,_T_84}; // @[AWSVggWrapper.scala 52:94]
  assign _T_340 = {_T_339,_T_85}; // @[AWSVggWrapper.scala 52:94]
  assign _T_341 = {_T_340,_T_86}; // @[AWSVggWrapper.scala 52:94]
  assign _T_342 = {_T_341,_T_87}; // @[AWSVggWrapper.scala 52:94]
  assign _T_343 = {_T_342,_T_88}; // @[AWSVggWrapper.scala 52:94]
  assign _T_344 = {_T_343,_T_89}; // @[AWSVggWrapper.scala 52:94]
  assign _T_345 = {_T_344,_T_90}; // @[AWSVggWrapper.scala 52:94]
  assign _T_346 = {_T_345,_T_91}; // @[AWSVggWrapper.scala 52:94]
  assign _T_347 = {_T_346,_T_92}; // @[AWSVggWrapper.scala 52:94]
  assign _T_348 = {_T_347,_T_93}; // @[AWSVggWrapper.scala 52:94]
  assign _T_349 = {_T_348,_T_94}; // @[AWSVggWrapper.scala 52:94]
  assign _T_350 = {_T_349,_T_95}; // @[AWSVggWrapper.scala 52:94]
  assign _T_351 = {_T_350,_T_96}; // @[AWSVggWrapper.scala 52:94]
  assign _T_352 = {_T_351,_T_97}; // @[AWSVggWrapper.scala 52:94]
  assign _T_353 = {_T_352,_T_98}; // @[AWSVggWrapper.scala 52:94]
  assign _T_354 = {_T_353,_T_99}; // @[AWSVggWrapper.scala 52:94]
  assign _T_355 = {_T_354,_T_100}; // @[AWSVggWrapper.scala 52:94]
  assign _T_356 = {_T_355,_T_101}; // @[AWSVggWrapper.scala 52:94]
  assign _T_357 = {_T_356,_T_102}; // @[AWSVggWrapper.scala 52:94]
  assign _T_358 = {_T_357,_T_103}; // @[AWSVggWrapper.scala 52:94]
  assign _T_359 = {_T_358,_T_104}; // @[AWSVggWrapper.scala 52:94]
  assign _T_360 = {_T_359,_T_105}; // @[AWSVggWrapper.scala 52:94]
  assign _T_361 = {_T_360,_T_106}; // @[AWSVggWrapper.scala 52:94]
  assign _T_362 = {_T_361,_T_107}; // @[AWSVggWrapper.scala 52:94]
  assign _T_363 = {_T_362,_T_108}; // @[AWSVggWrapper.scala 52:94]
  assign _T_364 = {_T_363,_T_109}; // @[AWSVggWrapper.scala 52:94]
  assign _T_365 = {_T_364,_T_110}; // @[AWSVggWrapper.scala 52:94]
  assign _T_366 = {_T_365,_T_111}; // @[AWSVggWrapper.scala 52:94]
  assign _T_367 = {_T_366,_T_112}; // @[AWSVggWrapper.scala 52:94]
  assign _T_368 = {_T_367,_T_113}; // @[AWSVggWrapper.scala 52:94]
  assign _T_369 = {_T_368,_T_114}; // @[AWSVggWrapper.scala 52:94]
  assign _T_370 = {_T_369,_T_115}; // @[AWSVggWrapper.scala 52:94]
  assign _T_371 = {_T_370,_T_116}; // @[AWSVggWrapper.scala 52:94]
  assign _T_372 = {_T_371,_T_117}; // @[AWSVggWrapper.scala 52:94]
  assign _T_373 = {_T_372,_T_118}; // @[AWSVggWrapper.scala 52:94]
  assign _T_374 = {_T_373,_T_119}; // @[AWSVggWrapper.scala 52:94]
  assign _T_375 = {_T_374,_T_120}; // @[AWSVggWrapper.scala 52:94]
  assign _T_376 = {_T_375,_T_121}; // @[AWSVggWrapper.scala 52:94]
  assign _T_377 = {_T_376,_T_122}; // @[AWSVggWrapper.scala 52:94]
  assign _T_378 = {_T_377,_T_123}; // @[AWSVggWrapper.scala 52:94]
  assign _T_379 = {_T_378,_T_124}; // @[AWSVggWrapper.scala 52:94]
  assign _T_380 = {_T_379,_T_125}; // @[AWSVggWrapper.scala 52:94]
  assign _T_381 = {_T_380,_T_126}; // @[AWSVggWrapper.scala 52:94]
  assign _T_382 = {_T_381,_T_127}; // @[AWSVggWrapper.scala 52:94]
  assign _T_383 = {_T_382,_T_128}; // @[AWSVggWrapper.scala 52:94]
  assign _T_384 = {_T_383,_T_129}; // @[AWSVggWrapper.scala 52:94]
  assign _T_385 = {_T_384,_T_130}; // @[AWSVggWrapper.scala 52:94]
  assign _T_386 = {_T_385,_T_131}; // @[AWSVggWrapper.scala 52:94]
  assign _T_387 = {_T_386,_T_132}; // @[AWSVggWrapper.scala 52:94]
  assign _T_388 = {_T_387,_T_133}; // @[AWSVggWrapper.scala 52:94]
  assign _T_389 = {_T_388,_T_134}; // @[AWSVggWrapper.scala 52:94]
  assign _T_390 = {_T_389,_T_135}; // @[AWSVggWrapper.scala 52:94]
  assign _T_391 = {_T_390,_T_136}; // @[AWSVggWrapper.scala 52:94]
  assign _T_392 = {_T_391,_T_137}; // @[AWSVggWrapper.scala 52:94]
  assign _T_393 = {_T_392,_T_138}; // @[AWSVggWrapper.scala 52:94]
  assign _T_394 = {_T_393,_T_139}; // @[AWSVggWrapper.scala 52:94]
  assign _T_395 = {_T_394,_T_140}; // @[AWSVggWrapper.scala 52:94]
  assign _T_396 = {_T_395,_T_141}; // @[AWSVggWrapper.scala 52:94]
  assign _T_397 = {_T_396,_T_142}; // @[AWSVggWrapper.scala 52:94]
  assign _T_398 = {_T_397,_T_143}; // @[AWSVggWrapper.scala 52:94]
  assign _T_399 = {_T_398,_T_144}; // @[AWSVggWrapper.scala 52:94]
  assign _T_400 = {_T_399,_T_145}; // @[AWSVggWrapper.scala 52:94]
  assign _T_401 = {_T_400,_T_146}; // @[AWSVggWrapper.scala 52:94]
  assign _T_402 = {_T_401,_T_147}; // @[AWSVggWrapper.scala 52:94]
  assign _T_403 = {_T_402,_T_148}; // @[AWSVggWrapper.scala 52:94]
  assign _T_404 = {_T_403,_T_149}; // @[AWSVggWrapper.scala 52:94]
  assign _T_405 = {_T_404,_T_150}; // @[AWSVggWrapper.scala 52:94]
  assign _T_406 = {_T_405,_T_151}; // @[AWSVggWrapper.scala 52:94]
  assign _T_407 = {_T_406,_T_152}; // @[AWSVggWrapper.scala 52:94]
  assign _T_408 = {_T_407,_T_153}; // @[AWSVggWrapper.scala 52:94]
  assign _T_409 = {_T_408,_T_154}; // @[AWSVggWrapper.scala 52:94]
  assign _T_410 = {_T_409,_T_155}; // @[AWSVggWrapper.scala 52:94]
  assign _T_411 = {_T_410,_T_156}; // @[AWSVggWrapper.scala 52:94]
  assign _T_412 = {_T_411,_T_157}; // @[AWSVggWrapper.scala 52:94]
  assign _T_413 = {_T_412,_T_158}; // @[AWSVggWrapper.scala 52:94]
  assign _T_414 = {_T_413,_T_159}; // @[AWSVggWrapper.scala 52:94]
  assign _T_415 = {_T_414,_T_160}; // @[AWSVggWrapper.scala 52:94]
  assign _T_416 = {_T_415,_T_161}; // @[AWSVggWrapper.scala 52:94]
  assign _T_417 = {_T_416,_T_162}; // @[AWSVggWrapper.scala 52:94]
  assign _T_418 = {_T_417,_T_163}; // @[AWSVggWrapper.scala 52:94]
  assign _T_419 = {_T_418,_T_164}; // @[AWSVggWrapper.scala 52:94]
  assign _T_420 = {_T_419,_T_165}; // @[AWSVggWrapper.scala 52:94]
  assign _T_421 = {_T_420,_T_166}; // @[AWSVggWrapper.scala 52:94]
  assign _T_422 = {_T_421,_T_167}; // @[AWSVggWrapper.scala 52:94]
  assign _T_423 = {_T_422,_T_168}; // @[AWSVggWrapper.scala 52:94]
  assign _T_424 = {_T_423,_T_169}; // @[AWSVggWrapper.scala 52:94]
  assign _T_425 = {_T_424,_T_170}; // @[AWSVggWrapper.scala 52:94]
  assign _T_426 = {_T_425,_T_171}; // @[AWSVggWrapper.scala 52:94]
  assign _T_427 = {_T_426,_T_172}; // @[AWSVggWrapper.scala 52:94]
  assign _T_428 = {_T_427,_T_173}; // @[AWSVggWrapper.scala 52:94]
  assign _T_429 = {_T_428,_T_174}; // @[AWSVggWrapper.scala 52:94]
  assign _T_430 = {_T_429,_T_175}; // @[AWSVggWrapper.scala 52:94]
  assign _T_431 = {_T_430,_T_176}; // @[AWSVggWrapper.scala 52:94]
  assign _T_432 = {_T_431,_T_177}; // @[AWSVggWrapper.scala 52:94]
  assign _T_433 = {_T_432,_T_178}; // @[AWSVggWrapper.scala 52:94]
  assign _T_434 = {_T_433,_T_179}; // @[AWSVggWrapper.scala 52:94]
  assign _T_435 = {_T_434,_T_180}; // @[AWSVggWrapper.scala 52:94]
  assign _T_436 = {_T_435,_T_181}; // @[AWSVggWrapper.scala 52:94]
  assign _T_437 = {_T_436,_T_182}; // @[AWSVggWrapper.scala 52:94]
  assign _T_438 = {_T_437,_T_183}; // @[AWSVggWrapper.scala 52:94]
  assign _T_439 = {_T_438,_T_184}; // @[AWSVggWrapper.scala 52:94]
  assign _T_440 = {_T_439,_T_185}; // @[AWSVggWrapper.scala 52:94]
  assign _T_441 = {_T_440,_T_186}; // @[AWSVggWrapper.scala 52:94]
  assign _T_442 = {_T_441,_T_187}; // @[AWSVggWrapper.scala 52:94]
  assign _T_443 = {_T_442,_T_188}; // @[AWSVggWrapper.scala 52:94]
  assign _T_444 = {_T_443,_T_189}; // @[AWSVggWrapper.scala 52:94]
  assign _T_445 = {_T_444,_T_190}; // @[AWSVggWrapper.scala 52:94]
  assign _T_446 = {_T_445,_T_191}; // @[AWSVggWrapper.scala 52:94]
  assign _T_447 = {_T_446,_T_192}; // @[AWSVggWrapper.scala 52:94]
  assign _T_448 = {_T_447,_T_193}; // @[AWSVggWrapper.scala 52:94]
  assign _T_449 = {_T_448,_T_194}; // @[AWSVggWrapper.scala 52:94]
  assign _T_450 = {_T_449,_T_195}; // @[AWSVggWrapper.scala 52:94]
  assign _T_451 = {_T_450,_T_196}; // @[AWSVggWrapper.scala 52:94]
  assign _T_452 = {_T_451,_T_197}; // @[AWSVggWrapper.scala 52:94]
  assign _T_453 = {_T_452,_T_198}; // @[AWSVggWrapper.scala 52:94]
  assign _T_454 = {_T_453,_T_199}; // @[AWSVggWrapper.scala 52:94]
  assign _T_455 = {_T_454,_T_200}; // @[AWSVggWrapper.scala 52:94]
  assign _T_456 = {_T_455,_T_201}; // @[AWSVggWrapper.scala 52:94]
  assign _T_457 = {_T_456,_T_202}; // @[AWSVggWrapper.scala 52:94]
  assign _T_458 = {_T_457,_T_203}; // @[AWSVggWrapper.scala 52:94]
  assign _T_459 = {_T_458,_T_204}; // @[AWSVggWrapper.scala 52:94]
  assign _T_460 = {_T_459,_T_205}; // @[AWSVggWrapper.scala 52:94]
  assign _T_461 = {_T_460,_T_206}; // @[AWSVggWrapper.scala 52:94]
  assign _T_462 = {_T_461,_T_207}; // @[AWSVggWrapper.scala 52:94]
  assign _T_463 = {_T_462,_T_208}; // @[AWSVggWrapper.scala 52:94]
  assign _T_464 = {_T_463,_T_209}; // @[AWSVggWrapper.scala 52:94]
  assign _T_465 = {_T_464,_T_210}; // @[AWSVggWrapper.scala 52:94]
  assign _T_466 = {_T_465,_T_211}; // @[AWSVggWrapper.scala 52:94]
  assign _T_467 = {_T_466,_T_212}; // @[AWSVggWrapper.scala 52:94]
  assign _T_468 = {_T_467,_T_213}; // @[AWSVggWrapper.scala 52:94]
  assign _T_469 = {_T_468,_T_214}; // @[AWSVggWrapper.scala 52:94]
  assign _T_470 = {_T_469,_T_215}; // @[AWSVggWrapper.scala 52:94]
  assign _T_471 = {_T_470,_T_216}; // @[AWSVggWrapper.scala 52:94]
  assign _T_472 = {_T_471,_T_217}; // @[AWSVggWrapper.scala 52:94]
  assign _T_473 = {_T_472,_T_218}; // @[AWSVggWrapper.scala 52:94]
  assign _T_474 = {_T_473,_T_219}; // @[AWSVggWrapper.scala 52:94]
  assign _T_475 = {_T_474,_T_220}; // @[AWSVggWrapper.scala 52:94]
  assign _T_476 = {_T_475,_T_221}; // @[AWSVggWrapper.scala 52:94]
  assign _T_477 = {_T_476,_T_222}; // @[AWSVggWrapper.scala 52:94]
  assign _T_478 = {_T_477,_T_223}; // @[AWSVggWrapper.scala 52:94]
  assign _T_479 = {_T_478,_T_224}; // @[AWSVggWrapper.scala 52:94]
  assign _T_480 = {_T_479,_T_225}; // @[AWSVggWrapper.scala 52:94]
  assign _T_481 = {_T_480,_T_226}; // @[AWSVggWrapper.scala 52:94]
  assign _T_482 = {_T_481,_T_227}; // @[AWSVggWrapper.scala 52:94]
  assign _T_483 = {_T_482,_T_228}; // @[AWSVggWrapper.scala 52:94]
  assign _T_484 = {_T_483,_T_229}; // @[AWSVggWrapper.scala 52:94]
  assign _T_485 = {_T_484,_T_230}; // @[AWSVggWrapper.scala 52:94]
  assign _T_486 = {_T_485,_T_231}; // @[AWSVggWrapper.scala 52:94]
  assign _T_487 = {_T_486,_T_232}; // @[AWSVggWrapper.scala 52:94]
  assign _T_488 = {_T_487,_T_233}; // @[AWSVggWrapper.scala 52:94]
  assign _T_489 = {_T_488,_T_234}; // @[AWSVggWrapper.scala 52:94]
  assign _T_490 = {_T_489,_T_235}; // @[AWSVggWrapper.scala 52:94]
  assign _T_491 = {_T_490,_T_236}; // @[AWSVggWrapper.scala 52:94]
  assign _T_492 = {_T_491,_T_237}; // @[AWSVggWrapper.scala 52:94]
  assign _T_493 = {_T_492,_T_238}; // @[AWSVggWrapper.scala 52:94]
  assign _T_494 = {_T_493,_T_239}; // @[AWSVggWrapper.scala 52:94]
  assign _T_495 = {_T_494,_T_240}; // @[AWSVggWrapper.scala 52:94]
  assign _T_496 = {_T_495,_T_241}; // @[AWSVggWrapper.scala 52:94]
  assign _T_497 = {_T_496,_T_242}; // @[AWSVggWrapper.scala 52:94]
  assign _T_498 = {_T_497,_T_243}; // @[AWSVggWrapper.scala 52:94]
  assign _T_499 = {_T_498,_T_244}; // @[AWSVggWrapper.scala 52:94]
  assign _T_500 = {_T_499,_T_245}; // @[AWSVggWrapper.scala 52:94]
  assign _T_501 = {_T_500,_T_246}; // @[AWSVggWrapper.scala 52:94]
  assign _T_502 = {_T_501,_T_247}; // @[AWSVggWrapper.scala 52:94]
  assign _T_503 = {_T_502,_T_248}; // @[AWSVggWrapper.scala 52:94]
  assign _T_504 = {_T_503,_T_249}; // @[AWSVggWrapper.scala 52:94]
  assign _T_505 = {_T_504,_T_250}; // @[AWSVggWrapper.scala 52:94]
  assign _T_506 = {_T_505,_T_251}; // @[AWSVggWrapper.scala 52:94]
  assign _T_507 = {_T_506,_T_252}; // @[AWSVggWrapper.scala 52:94]
  assign _T_508 = {_T_507,_T_253}; // @[AWSVggWrapper.scala 52:94]
  assign _T_509 = {_T_508,_T_254}; // @[AWSVggWrapper.scala 52:94]
  assign _T_510 = {_T_509,_T_255}; // @[AWSVggWrapper.scala 52:94]
  assign _T_511 = {_T_510,_T_256}; // @[AWSVggWrapper.scala 52:94]
  assign _T_512 = {_T_511,_T_257}; // @[AWSVggWrapper.scala 52:94]
  assign _T_513 = {_T_512,_T_258}; // @[AWSVggWrapper.scala 52:94]
  assign _T_514 = {_T_513,_T_259}; // @[AWSVggWrapper.scala 52:94]
  assign _T_515 = {_T_514,_T_260}; // @[AWSVggWrapper.scala 52:94]
  assign _T_516 = {_T_515,_T_261}; // @[AWSVggWrapper.scala 52:94]
  assign _T_517 = {_T_516,_T_262}; // @[AWSVggWrapper.scala 52:94]
  assign _T_518 = {_T_517,_T_263}; // @[AWSVggWrapper.scala 52:94]
  assign _T_519 = {_T_518,_T_264}; // @[AWSVggWrapper.scala 52:94]
  assign _T_520 = {_T_519,_T_265}; // @[AWSVggWrapper.scala 52:94]
  assign _T_521 = {_T_520,_T_266}; // @[AWSVggWrapper.scala 52:94]
  assign _T_522 = {_T_521,_T_267}; // @[AWSVggWrapper.scala 52:94]
  assign _T_523 = {_T_522,_T_268}; // @[AWSVggWrapper.scala 52:94]
  assign _T_524 = {_T_523,_T_269}; // @[AWSVggWrapper.scala 52:94]
  assign _T_525 = {_T_524,_T_270}; // @[AWSVggWrapper.scala 52:94]
  assign _T_526 = {_T_525,_T_271}; // @[AWSVggWrapper.scala 52:94]
  assign _T_527 = {_T_526,_T_272}; // @[AWSVggWrapper.scala 52:94]
  assign _T_528 = {_T_527,_T_273}; // @[AWSVggWrapper.scala 52:94]
  assign _T_529 = {_T_528,_T_274}; // @[AWSVggWrapper.scala 52:94]
  assign _T_530 = {_T_529,_T_275}; // @[AWSVggWrapper.scala 52:94]
  assign _T_531 = {_T_530,_T_276}; // @[AWSVggWrapper.scala 52:94]
  assign _T_532 = {_T_531,_T_277}; // @[AWSVggWrapper.scala 52:94]
  assign _T_533 = {_T_532,_T_278}; // @[AWSVggWrapper.scala 52:94]
  assign _T_534 = {_T_533,_T_279}; // @[AWSVggWrapper.scala 52:94]
  assign _T_535 = {_T_534,_T_280}; // @[AWSVggWrapper.scala 52:94]
  assign _T_536 = {_T_535,_T_281}; // @[AWSVggWrapper.scala 52:94]
  assign _T_537 = {_T_536,_T_282}; // @[AWSVggWrapper.scala 52:94]
  assign _T_538 = {_T_537,_T_283}; // @[AWSVggWrapper.scala 52:94]
  assign dataInAsUInt = {_T_538,_T_284}; // @[AWSVggWrapper.scala 52:94]
  assign _T_1833 = queueIOOut_io_deq_bits[15:0]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_255 = $signed(_T_1833); // @[AWSVggWrapper.scala 63:110]
  assign _T_1835 = queueIOOut_io_deq_bits[31:16]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_254 = $signed(_T_1835); // @[AWSVggWrapper.scala 63:110]
  assign _T_1837 = queueIOOut_io_deq_bits[47:32]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_253 = $signed(_T_1837); // @[AWSVggWrapper.scala 63:110]
  assign _T_1839 = queueIOOut_io_deq_bits[63:48]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_252 = $signed(_T_1839); // @[AWSVggWrapper.scala 63:110]
  assign _T_1841 = queueIOOut_io_deq_bits[79:64]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_251 = $signed(_T_1841); // @[AWSVggWrapper.scala 63:110]
  assign _T_1843 = queueIOOut_io_deq_bits[95:80]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_250 = $signed(_T_1843); // @[AWSVggWrapper.scala 63:110]
  assign _T_1845 = queueIOOut_io_deq_bits[111:96]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_249 = $signed(_T_1845); // @[AWSVggWrapper.scala 63:110]
  assign _T_1847 = queueIOOut_io_deq_bits[127:112]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_248 = $signed(_T_1847); // @[AWSVggWrapper.scala 63:110]
  assign _T_1849 = queueIOOut_io_deq_bits[143:128]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_247 = $signed(_T_1849); // @[AWSVggWrapper.scala 63:110]
  assign _T_1851 = queueIOOut_io_deq_bits[159:144]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_246 = $signed(_T_1851); // @[AWSVggWrapper.scala 63:110]
  assign _T_1853 = queueIOOut_io_deq_bits[175:160]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_245 = $signed(_T_1853); // @[AWSVggWrapper.scala 63:110]
  assign _T_1855 = queueIOOut_io_deq_bits[191:176]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_244 = $signed(_T_1855); // @[AWSVggWrapper.scala 63:110]
  assign _T_1857 = queueIOOut_io_deq_bits[207:192]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_243 = $signed(_T_1857); // @[AWSVggWrapper.scala 63:110]
  assign _T_1859 = queueIOOut_io_deq_bits[223:208]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_242 = $signed(_T_1859); // @[AWSVggWrapper.scala 63:110]
  assign _T_1861 = queueIOOut_io_deq_bits[239:224]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_241 = $signed(_T_1861); // @[AWSVggWrapper.scala 63:110]
  assign _T_1863 = queueIOOut_io_deq_bits[255:240]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_240 = $signed(_T_1863); // @[AWSVggWrapper.scala 63:110]
  assign _T_1865 = queueIOOut_io_deq_bits[271:256]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_239 = $signed(_T_1865); // @[AWSVggWrapper.scala 63:110]
  assign _T_1867 = queueIOOut_io_deq_bits[287:272]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_238 = $signed(_T_1867); // @[AWSVggWrapper.scala 63:110]
  assign _T_1869 = queueIOOut_io_deq_bits[303:288]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_237 = $signed(_T_1869); // @[AWSVggWrapper.scala 63:110]
  assign _T_1871 = queueIOOut_io_deq_bits[319:304]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_236 = $signed(_T_1871); // @[AWSVggWrapper.scala 63:110]
  assign _T_1873 = queueIOOut_io_deq_bits[335:320]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_235 = $signed(_T_1873); // @[AWSVggWrapper.scala 63:110]
  assign _T_1875 = queueIOOut_io_deq_bits[351:336]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_234 = $signed(_T_1875); // @[AWSVggWrapper.scala 63:110]
  assign _T_1877 = queueIOOut_io_deq_bits[367:352]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_233 = $signed(_T_1877); // @[AWSVggWrapper.scala 63:110]
  assign _T_1879 = queueIOOut_io_deq_bits[383:368]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_232 = $signed(_T_1879); // @[AWSVggWrapper.scala 63:110]
  assign _T_1881 = queueIOOut_io_deq_bits[399:384]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_231 = $signed(_T_1881); // @[AWSVggWrapper.scala 63:110]
  assign _T_1883 = queueIOOut_io_deq_bits[415:400]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_230 = $signed(_T_1883); // @[AWSVggWrapper.scala 63:110]
  assign _T_1885 = queueIOOut_io_deq_bits[431:416]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_229 = $signed(_T_1885); // @[AWSVggWrapper.scala 63:110]
  assign _T_1887 = queueIOOut_io_deq_bits[447:432]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_228 = $signed(_T_1887); // @[AWSVggWrapper.scala 63:110]
  assign _T_1889 = queueIOOut_io_deq_bits[463:448]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_227 = $signed(_T_1889); // @[AWSVggWrapper.scala 63:110]
  assign _T_1891 = queueIOOut_io_deq_bits[479:464]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_226 = $signed(_T_1891); // @[AWSVggWrapper.scala 63:110]
  assign _T_1893 = queueIOOut_io_deq_bits[495:480]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_225 = $signed(_T_1893); // @[AWSVggWrapper.scala 63:110]
  assign _T_1895 = queueIOOut_io_deq_bits[511:496]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_224 = $signed(_T_1895); // @[AWSVggWrapper.scala 63:110]
  assign _T_1897 = queueIOOut_io_deq_bits[527:512]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_223 = $signed(_T_1897); // @[AWSVggWrapper.scala 63:110]
  assign _T_1899 = queueIOOut_io_deq_bits[543:528]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_222 = $signed(_T_1899); // @[AWSVggWrapper.scala 63:110]
  assign _T_1901 = queueIOOut_io_deq_bits[559:544]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_221 = $signed(_T_1901); // @[AWSVggWrapper.scala 63:110]
  assign _T_1903 = queueIOOut_io_deq_bits[575:560]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_220 = $signed(_T_1903); // @[AWSVggWrapper.scala 63:110]
  assign _T_1905 = queueIOOut_io_deq_bits[591:576]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_219 = $signed(_T_1905); // @[AWSVggWrapper.scala 63:110]
  assign _T_1907 = queueIOOut_io_deq_bits[607:592]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_218 = $signed(_T_1907); // @[AWSVggWrapper.scala 63:110]
  assign _T_1909 = queueIOOut_io_deq_bits[623:608]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_217 = $signed(_T_1909); // @[AWSVggWrapper.scala 63:110]
  assign _T_1911 = queueIOOut_io_deq_bits[639:624]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_216 = $signed(_T_1911); // @[AWSVggWrapper.scala 63:110]
  assign _T_1913 = queueIOOut_io_deq_bits[655:640]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_215 = $signed(_T_1913); // @[AWSVggWrapper.scala 63:110]
  assign _T_1915 = queueIOOut_io_deq_bits[671:656]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_214 = $signed(_T_1915); // @[AWSVggWrapper.scala 63:110]
  assign _T_1917 = queueIOOut_io_deq_bits[687:672]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_213 = $signed(_T_1917); // @[AWSVggWrapper.scala 63:110]
  assign _T_1919 = queueIOOut_io_deq_bits[703:688]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_212 = $signed(_T_1919); // @[AWSVggWrapper.scala 63:110]
  assign _T_1921 = queueIOOut_io_deq_bits[719:704]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_211 = $signed(_T_1921); // @[AWSVggWrapper.scala 63:110]
  assign _T_1923 = queueIOOut_io_deq_bits[735:720]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_210 = $signed(_T_1923); // @[AWSVggWrapper.scala 63:110]
  assign _T_1925 = queueIOOut_io_deq_bits[751:736]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_209 = $signed(_T_1925); // @[AWSVggWrapper.scala 63:110]
  assign _T_1927 = queueIOOut_io_deq_bits[767:752]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_208 = $signed(_T_1927); // @[AWSVggWrapper.scala 63:110]
  assign _T_1929 = queueIOOut_io_deq_bits[783:768]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_207 = $signed(_T_1929); // @[AWSVggWrapper.scala 63:110]
  assign _T_1931 = queueIOOut_io_deq_bits[799:784]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_206 = $signed(_T_1931); // @[AWSVggWrapper.scala 63:110]
  assign _T_1933 = queueIOOut_io_deq_bits[815:800]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_205 = $signed(_T_1933); // @[AWSVggWrapper.scala 63:110]
  assign _T_1935 = queueIOOut_io_deq_bits[831:816]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_204 = $signed(_T_1935); // @[AWSVggWrapper.scala 63:110]
  assign _T_1937 = queueIOOut_io_deq_bits[847:832]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_203 = $signed(_T_1937); // @[AWSVggWrapper.scala 63:110]
  assign _T_1939 = queueIOOut_io_deq_bits[863:848]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_202 = $signed(_T_1939); // @[AWSVggWrapper.scala 63:110]
  assign _T_1941 = queueIOOut_io_deq_bits[879:864]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_201 = $signed(_T_1941); // @[AWSVggWrapper.scala 63:110]
  assign _T_1943 = queueIOOut_io_deq_bits[895:880]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_200 = $signed(_T_1943); // @[AWSVggWrapper.scala 63:110]
  assign _T_1945 = queueIOOut_io_deq_bits[911:896]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_199 = $signed(_T_1945); // @[AWSVggWrapper.scala 63:110]
  assign _T_1947 = queueIOOut_io_deq_bits[927:912]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_198 = $signed(_T_1947); // @[AWSVggWrapper.scala 63:110]
  assign _T_1949 = queueIOOut_io_deq_bits[943:928]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_197 = $signed(_T_1949); // @[AWSVggWrapper.scala 63:110]
  assign _T_1951 = queueIOOut_io_deq_bits[959:944]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_196 = $signed(_T_1951); // @[AWSVggWrapper.scala 63:110]
  assign _T_1953 = queueIOOut_io_deq_bits[975:960]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_195 = $signed(_T_1953); // @[AWSVggWrapper.scala 63:110]
  assign _T_1955 = queueIOOut_io_deq_bits[991:976]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_194 = $signed(_T_1955); // @[AWSVggWrapper.scala 63:110]
  assign _T_1957 = queueIOOut_io_deq_bits[1007:992]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_193 = $signed(_T_1957); // @[AWSVggWrapper.scala 63:110]
  assign _T_1959 = queueIOOut_io_deq_bits[1023:1008]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_192 = $signed(_T_1959); // @[AWSVggWrapper.scala 63:110]
  assign _T_1961 = queueIOOut_io_deq_bits[1039:1024]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_191 = $signed(_T_1961); // @[AWSVggWrapper.scala 63:110]
  assign _T_1963 = queueIOOut_io_deq_bits[1055:1040]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_190 = $signed(_T_1963); // @[AWSVggWrapper.scala 63:110]
  assign _T_1965 = queueIOOut_io_deq_bits[1071:1056]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_189 = $signed(_T_1965); // @[AWSVggWrapper.scala 63:110]
  assign _T_1967 = queueIOOut_io_deq_bits[1087:1072]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_188 = $signed(_T_1967); // @[AWSVggWrapper.scala 63:110]
  assign _T_1969 = queueIOOut_io_deq_bits[1103:1088]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_187 = $signed(_T_1969); // @[AWSVggWrapper.scala 63:110]
  assign _T_1971 = queueIOOut_io_deq_bits[1119:1104]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_186 = $signed(_T_1971); // @[AWSVggWrapper.scala 63:110]
  assign _T_1973 = queueIOOut_io_deq_bits[1135:1120]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_185 = $signed(_T_1973); // @[AWSVggWrapper.scala 63:110]
  assign _T_1975 = queueIOOut_io_deq_bits[1151:1136]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_184 = $signed(_T_1975); // @[AWSVggWrapper.scala 63:110]
  assign _T_1977 = queueIOOut_io_deq_bits[1167:1152]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_183 = $signed(_T_1977); // @[AWSVggWrapper.scala 63:110]
  assign _T_1979 = queueIOOut_io_deq_bits[1183:1168]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_182 = $signed(_T_1979); // @[AWSVggWrapper.scala 63:110]
  assign _T_1981 = queueIOOut_io_deq_bits[1199:1184]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_181 = $signed(_T_1981); // @[AWSVggWrapper.scala 63:110]
  assign _T_1983 = queueIOOut_io_deq_bits[1215:1200]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_180 = $signed(_T_1983); // @[AWSVggWrapper.scala 63:110]
  assign _T_1985 = queueIOOut_io_deq_bits[1231:1216]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_179 = $signed(_T_1985); // @[AWSVggWrapper.scala 63:110]
  assign _T_1987 = queueIOOut_io_deq_bits[1247:1232]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_178 = $signed(_T_1987); // @[AWSVggWrapper.scala 63:110]
  assign _T_1989 = queueIOOut_io_deq_bits[1263:1248]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_177 = $signed(_T_1989); // @[AWSVggWrapper.scala 63:110]
  assign _T_1991 = queueIOOut_io_deq_bits[1279:1264]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_176 = $signed(_T_1991); // @[AWSVggWrapper.scala 63:110]
  assign _T_1993 = queueIOOut_io_deq_bits[1295:1280]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_175 = $signed(_T_1993); // @[AWSVggWrapper.scala 63:110]
  assign _T_1995 = queueIOOut_io_deq_bits[1311:1296]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_174 = $signed(_T_1995); // @[AWSVggWrapper.scala 63:110]
  assign _T_1997 = queueIOOut_io_deq_bits[1327:1312]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_173 = $signed(_T_1997); // @[AWSVggWrapper.scala 63:110]
  assign _T_1999 = queueIOOut_io_deq_bits[1343:1328]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_172 = $signed(_T_1999); // @[AWSVggWrapper.scala 63:110]
  assign _T_2001 = queueIOOut_io_deq_bits[1359:1344]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_171 = $signed(_T_2001); // @[AWSVggWrapper.scala 63:110]
  assign _T_2003 = queueIOOut_io_deq_bits[1375:1360]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_170 = $signed(_T_2003); // @[AWSVggWrapper.scala 63:110]
  assign _T_2005 = queueIOOut_io_deq_bits[1391:1376]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_169 = $signed(_T_2005); // @[AWSVggWrapper.scala 63:110]
  assign _T_2007 = queueIOOut_io_deq_bits[1407:1392]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_168 = $signed(_T_2007); // @[AWSVggWrapper.scala 63:110]
  assign _T_2009 = queueIOOut_io_deq_bits[1423:1408]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_167 = $signed(_T_2009); // @[AWSVggWrapper.scala 63:110]
  assign _T_2011 = queueIOOut_io_deq_bits[1439:1424]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_166 = $signed(_T_2011); // @[AWSVggWrapper.scala 63:110]
  assign _T_2013 = queueIOOut_io_deq_bits[1455:1440]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_165 = $signed(_T_2013); // @[AWSVggWrapper.scala 63:110]
  assign _T_2015 = queueIOOut_io_deq_bits[1471:1456]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_164 = $signed(_T_2015); // @[AWSVggWrapper.scala 63:110]
  assign _T_2017 = queueIOOut_io_deq_bits[1487:1472]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_163 = $signed(_T_2017); // @[AWSVggWrapper.scala 63:110]
  assign _T_2019 = queueIOOut_io_deq_bits[1503:1488]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_162 = $signed(_T_2019); // @[AWSVggWrapper.scala 63:110]
  assign _T_2021 = queueIOOut_io_deq_bits[1519:1504]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_161 = $signed(_T_2021); // @[AWSVggWrapper.scala 63:110]
  assign _T_2023 = queueIOOut_io_deq_bits[1535:1520]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_160 = $signed(_T_2023); // @[AWSVggWrapper.scala 63:110]
  assign _T_2025 = queueIOOut_io_deq_bits[1551:1536]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_159 = $signed(_T_2025); // @[AWSVggWrapper.scala 63:110]
  assign _T_2027 = queueIOOut_io_deq_bits[1567:1552]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_158 = $signed(_T_2027); // @[AWSVggWrapper.scala 63:110]
  assign _T_2029 = queueIOOut_io_deq_bits[1583:1568]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_157 = $signed(_T_2029); // @[AWSVggWrapper.scala 63:110]
  assign _T_2031 = queueIOOut_io_deq_bits[1599:1584]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_156 = $signed(_T_2031); // @[AWSVggWrapper.scala 63:110]
  assign _T_2033 = queueIOOut_io_deq_bits[1615:1600]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_155 = $signed(_T_2033); // @[AWSVggWrapper.scala 63:110]
  assign _T_2035 = queueIOOut_io_deq_bits[1631:1616]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_154 = $signed(_T_2035); // @[AWSVggWrapper.scala 63:110]
  assign _T_2037 = queueIOOut_io_deq_bits[1647:1632]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_153 = $signed(_T_2037); // @[AWSVggWrapper.scala 63:110]
  assign _T_2039 = queueIOOut_io_deq_bits[1663:1648]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_152 = $signed(_T_2039); // @[AWSVggWrapper.scala 63:110]
  assign _T_2041 = queueIOOut_io_deq_bits[1679:1664]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_151 = $signed(_T_2041); // @[AWSVggWrapper.scala 63:110]
  assign _T_2043 = queueIOOut_io_deq_bits[1695:1680]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_150 = $signed(_T_2043); // @[AWSVggWrapper.scala 63:110]
  assign _T_2045 = queueIOOut_io_deq_bits[1711:1696]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_149 = $signed(_T_2045); // @[AWSVggWrapper.scala 63:110]
  assign _T_2047 = queueIOOut_io_deq_bits[1727:1712]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_148 = $signed(_T_2047); // @[AWSVggWrapper.scala 63:110]
  assign _T_2049 = queueIOOut_io_deq_bits[1743:1728]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_147 = $signed(_T_2049); // @[AWSVggWrapper.scala 63:110]
  assign _T_2051 = queueIOOut_io_deq_bits[1759:1744]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_146 = $signed(_T_2051); // @[AWSVggWrapper.scala 63:110]
  assign _T_2053 = queueIOOut_io_deq_bits[1775:1760]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_145 = $signed(_T_2053); // @[AWSVggWrapper.scala 63:110]
  assign _T_2055 = queueIOOut_io_deq_bits[1791:1776]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_144 = $signed(_T_2055); // @[AWSVggWrapper.scala 63:110]
  assign _T_2057 = queueIOOut_io_deq_bits[1807:1792]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_143 = $signed(_T_2057); // @[AWSVggWrapper.scala 63:110]
  assign _T_2059 = queueIOOut_io_deq_bits[1823:1808]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_142 = $signed(_T_2059); // @[AWSVggWrapper.scala 63:110]
  assign _T_2061 = queueIOOut_io_deq_bits[1839:1824]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_141 = $signed(_T_2061); // @[AWSVggWrapper.scala 63:110]
  assign _T_2063 = queueIOOut_io_deq_bits[1855:1840]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_140 = $signed(_T_2063); // @[AWSVggWrapper.scala 63:110]
  assign _T_2065 = queueIOOut_io_deq_bits[1871:1856]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_139 = $signed(_T_2065); // @[AWSVggWrapper.scala 63:110]
  assign _T_2067 = queueIOOut_io_deq_bits[1887:1872]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_138 = $signed(_T_2067); // @[AWSVggWrapper.scala 63:110]
  assign _T_2069 = queueIOOut_io_deq_bits[1903:1888]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_137 = $signed(_T_2069); // @[AWSVggWrapper.scala 63:110]
  assign _T_2071 = queueIOOut_io_deq_bits[1919:1904]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_136 = $signed(_T_2071); // @[AWSVggWrapper.scala 63:110]
  assign _T_2073 = queueIOOut_io_deq_bits[1935:1920]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_135 = $signed(_T_2073); // @[AWSVggWrapper.scala 63:110]
  assign _T_2075 = queueIOOut_io_deq_bits[1951:1936]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_134 = $signed(_T_2075); // @[AWSVggWrapper.scala 63:110]
  assign _T_2077 = queueIOOut_io_deq_bits[1967:1952]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_133 = $signed(_T_2077); // @[AWSVggWrapper.scala 63:110]
  assign _T_2079 = queueIOOut_io_deq_bits[1983:1968]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_132 = $signed(_T_2079); // @[AWSVggWrapper.scala 63:110]
  assign _T_2081 = queueIOOut_io_deq_bits[1999:1984]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_131 = $signed(_T_2081); // @[AWSVggWrapper.scala 63:110]
  assign _T_2083 = queueIOOut_io_deq_bits[2015:2000]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_130 = $signed(_T_2083); // @[AWSVggWrapper.scala 63:110]
  assign _T_2085 = queueIOOut_io_deq_bits[2031:2016]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_129 = $signed(_T_2085); // @[AWSVggWrapper.scala 63:110]
  assign _T_2087 = queueIOOut_io_deq_bits[2047:2032]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_128 = $signed(_T_2087); // @[AWSVggWrapper.scala 63:110]
  assign _T_2089 = queueIOOut_io_deq_bits[2063:2048]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_127 = $signed(_T_2089); // @[AWSVggWrapper.scala 63:110]
  assign _T_2091 = queueIOOut_io_deq_bits[2079:2064]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_126 = $signed(_T_2091); // @[AWSVggWrapper.scala 63:110]
  assign _T_2093 = queueIOOut_io_deq_bits[2095:2080]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_125 = $signed(_T_2093); // @[AWSVggWrapper.scala 63:110]
  assign _T_2095 = queueIOOut_io_deq_bits[2111:2096]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_124 = $signed(_T_2095); // @[AWSVggWrapper.scala 63:110]
  assign _T_2097 = queueIOOut_io_deq_bits[2127:2112]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_123 = $signed(_T_2097); // @[AWSVggWrapper.scala 63:110]
  assign _T_2099 = queueIOOut_io_deq_bits[2143:2128]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_122 = $signed(_T_2099); // @[AWSVggWrapper.scala 63:110]
  assign _T_2101 = queueIOOut_io_deq_bits[2159:2144]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_121 = $signed(_T_2101); // @[AWSVggWrapper.scala 63:110]
  assign _T_2103 = queueIOOut_io_deq_bits[2175:2160]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_120 = $signed(_T_2103); // @[AWSVggWrapper.scala 63:110]
  assign _T_2105 = queueIOOut_io_deq_bits[2191:2176]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_119 = $signed(_T_2105); // @[AWSVggWrapper.scala 63:110]
  assign _T_2107 = queueIOOut_io_deq_bits[2207:2192]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_118 = $signed(_T_2107); // @[AWSVggWrapper.scala 63:110]
  assign _T_2109 = queueIOOut_io_deq_bits[2223:2208]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_117 = $signed(_T_2109); // @[AWSVggWrapper.scala 63:110]
  assign _T_2111 = queueIOOut_io_deq_bits[2239:2224]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_116 = $signed(_T_2111); // @[AWSVggWrapper.scala 63:110]
  assign _T_2113 = queueIOOut_io_deq_bits[2255:2240]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_115 = $signed(_T_2113); // @[AWSVggWrapper.scala 63:110]
  assign _T_2115 = queueIOOut_io_deq_bits[2271:2256]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_114 = $signed(_T_2115); // @[AWSVggWrapper.scala 63:110]
  assign _T_2117 = queueIOOut_io_deq_bits[2287:2272]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_113 = $signed(_T_2117); // @[AWSVggWrapper.scala 63:110]
  assign _T_2119 = queueIOOut_io_deq_bits[2303:2288]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_112 = $signed(_T_2119); // @[AWSVggWrapper.scala 63:110]
  assign _T_2121 = queueIOOut_io_deq_bits[2319:2304]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_111 = $signed(_T_2121); // @[AWSVggWrapper.scala 63:110]
  assign _T_2123 = queueIOOut_io_deq_bits[2335:2320]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_110 = $signed(_T_2123); // @[AWSVggWrapper.scala 63:110]
  assign _T_2125 = queueIOOut_io_deq_bits[2351:2336]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_109 = $signed(_T_2125); // @[AWSVggWrapper.scala 63:110]
  assign _T_2127 = queueIOOut_io_deq_bits[2367:2352]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_108 = $signed(_T_2127); // @[AWSVggWrapper.scala 63:110]
  assign _T_2129 = queueIOOut_io_deq_bits[2383:2368]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_107 = $signed(_T_2129); // @[AWSVggWrapper.scala 63:110]
  assign _T_2131 = queueIOOut_io_deq_bits[2399:2384]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_106 = $signed(_T_2131); // @[AWSVggWrapper.scala 63:110]
  assign _T_2133 = queueIOOut_io_deq_bits[2415:2400]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_105 = $signed(_T_2133); // @[AWSVggWrapper.scala 63:110]
  assign _T_2135 = queueIOOut_io_deq_bits[2431:2416]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_104 = $signed(_T_2135); // @[AWSVggWrapper.scala 63:110]
  assign _T_2137 = queueIOOut_io_deq_bits[2447:2432]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_103 = $signed(_T_2137); // @[AWSVggWrapper.scala 63:110]
  assign _T_2139 = queueIOOut_io_deq_bits[2463:2448]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_102 = $signed(_T_2139); // @[AWSVggWrapper.scala 63:110]
  assign _T_2141 = queueIOOut_io_deq_bits[2479:2464]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_101 = $signed(_T_2141); // @[AWSVggWrapper.scala 63:110]
  assign _T_2143 = queueIOOut_io_deq_bits[2495:2480]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_100 = $signed(_T_2143); // @[AWSVggWrapper.scala 63:110]
  assign _T_2145 = queueIOOut_io_deq_bits[2511:2496]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_99 = $signed(_T_2145); // @[AWSVggWrapper.scala 63:110]
  assign _T_2147 = queueIOOut_io_deq_bits[2527:2512]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_98 = $signed(_T_2147); // @[AWSVggWrapper.scala 63:110]
  assign _T_2149 = queueIOOut_io_deq_bits[2543:2528]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_97 = $signed(_T_2149); // @[AWSVggWrapper.scala 63:110]
  assign _T_2151 = queueIOOut_io_deq_bits[2559:2544]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_96 = $signed(_T_2151); // @[AWSVggWrapper.scala 63:110]
  assign _T_2153 = queueIOOut_io_deq_bits[2575:2560]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_95 = $signed(_T_2153); // @[AWSVggWrapper.scala 63:110]
  assign _T_2155 = queueIOOut_io_deq_bits[2591:2576]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_94 = $signed(_T_2155); // @[AWSVggWrapper.scala 63:110]
  assign _T_2157 = queueIOOut_io_deq_bits[2607:2592]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_93 = $signed(_T_2157); // @[AWSVggWrapper.scala 63:110]
  assign _T_2159 = queueIOOut_io_deq_bits[2623:2608]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_92 = $signed(_T_2159); // @[AWSVggWrapper.scala 63:110]
  assign _T_2161 = queueIOOut_io_deq_bits[2639:2624]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_91 = $signed(_T_2161); // @[AWSVggWrapper.scala 63:110]
  assign _T_2163 = queueIOOut_io_deq_bits[2655:2640]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_90 = $signed(_T_2163); // @[AWSVggWrapper.scala 63:110]
  assign _T_2165 = queueIOOut_io_deq_bits[2671:2656]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_89 = $signed(_T_2165); // @[AWSVggWrapper.scala 63:110]
  assign _T_2167 = queueIOOut_io_deq_bits[2687:2672]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_88 = $signed(_T_2167); // @[AWSVggWrapper.scala 63:110]
  assign _T_2169 = queueIOOut_io_deq_bits[2703:2688]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_87 = $signed(_T_2169); // @[AWSVggWrapper.scala 63:110]
  assign _T_2171 = queueIOOut_io_deq_bits[2719:2704]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_86 = $signed(_T_2171); // @[AWSVggWrapper.scala 63:110]
  assign _T_2173 = queueIOOut_io_deq_bits[2735:2720]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_85 = $signed(_T_2173); // @[AWSVggWrapper.scala 63:110]
  assign _T_2175 = queueIOOut_io_deq_bits[2751:2736]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_84 = $signed(_T_2175); // @[AWSVggWrapper.scala 63:110]
  assign _T_2177 = queueIOOut_io_deq_bits[2767:2752]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_83 = $signed(_T_2177); // @[AWSVggWrapper.scala 63:110]
  assign _T_2179 = queueIOOut_io_deq_bits[2783:2768]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_82 = $signed(_T_2179); // @[AWSVggWrapper.scala 63:110]
  assign _T_2181 = queueIOOut_io_deq_bits[2799:2784]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_81 = $signed(_T_2181); // @[AWSVggWrapper.scala 63:110]
  assign _T_2183 = queueIOOut_io_deq_bits[2815:2800]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_80 = $signed(_T_2183); // @[AWSVggWrapper.scala 63:110]
  assign _T_2185 = queueIOOut_io_deq_bits[2831:2816]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_79 = $signed(_T_2185); // @[AWSVggWrapper.scala 63:110]
  assign _T_2187 = queueIOOut_io_deq_bits[2847:2832]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_78 = $signed(_T_2187); // @[AWSVggWrapper.scala 63:110]
  assign _T_2189 = queueIOOut_io_deq_bits[2863:2848]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_77 = $signed(_T_2189); // @[AWSVggWrapper.scala 63:110]
  assign _T_2191 = queueIOOut_io_deq_bits[2879:2864]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_76 = $signed(_T_2191); // @[AWSVggWrapper.scala 63:110]
  assign _T_2193 = queueIOOut_io_deq_bits[2895:2880]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_75 = $signed(_T_2193); // @[AWSVggWrapper.scala 63:110]
  assign _T_2195 = queueIOOut_io_deq_bits[2911:2896]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_74 = $signed(_T_2195); // @[AWSVggWrapper.scala 63:110]
  assign _T_2197 = queueIOOut_io_deq_bits[2927:2912]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_73 = $signed(_T_2197); // @[AWSVggWrapper.scala 63:110]
  assign _T_2199 = queueIOOut_io_deq_bits[2943:2928]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_72 = $signed(_T_2199); // @[AWSVggWrapper.scala 63:110]
  assign _T_2201 = queueIOOut_io_deq_bits[2959:2944]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_71 = $signed(_T_2201); // @[AWSVggWrapper.scala 63:110]
  assign _T_2203 = queueIOOut_io_deq_bits[2975:2960]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_70 = $signed(_T_2203); // @[AWSVggWrapper.scala 63:110]
  assign _T_2205 = queueIOOut_io_deq_bits[2991:2976]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_69 = $signed(_T_2205); // @[AWSVggWrapper.scala 63:110]
  assign _T_2207 = queueIOOut_io_deq_bits[3007:2992]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_68 = $signed(_T_2207); // @[AWSVggWrapper.scala 63:110]
  assign _T_2209 = queueIOOut_io_deq_bits[3023:3008]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_67 = $signed(_T_2209); // @[AWSVggWrapper.scala 63:110]
  assign _T_2211 = queueIOOut_io_deq_bits[3039:3024]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_66 = $signed(_T_2211); // @[AWSVggWrapper.scala 63:110]
  assign _T_2213 = queueIOOut_io_deq_bits[3055:3040]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_65 = $signed(_T_2213); // @[AWSVggWrapper.scala 63:110]
  assign _T_2215 = queueIOOut_io_deq_bits[3071:3056]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_64 = $signed(_T_2215); // @[AWSVggWrapper.scala 63:110]
  assign _T_2217 = queueIOOut_io_deq_bits[3087:3072]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_63 = $signed(_T_2217); // @[AWSVggWrapper.scala 63:110]
  assign _T_2219 = queueIOOut_io_deq_bits[3103:3088]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_62 = $signed(_T_2219); // @[AWSVggWrapper.scala 63:110]
  assign _T_2221 = queueIOOut_io_deq_bits[3119:3104]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_61 = $signed(_T_2221); // @[AWSVggWrapper.scala 63:110]
  assign _T_2223 = queueIOOut_io_deq_bits[3135:3120]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_60 = $signed(_T_2223); // @[AWSVggWrapper.scala 63:110]
  assign _T_2225 = queueIOOut_io_deq_bits[3151:3136]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_59 = $signed(_T_2225); // @[AWSVggWrapper.scala 63:110]
  assign _T_2227 = queueIOOut_io_deq_bits[3167:3152]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_58 = $signed(_T_2227); // @[AWSVggWrapper.scala 63:110]
  assign _T_2229 = queueIOOut_io_deq_bits[3183:3168]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_57 = $signed(_T_2229); // @[AWSVggWrapper.scala 63:110]
  assign _T_2231 = queueIOOut_io_deq_bits[3199:3184]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_56 = $signed(_T_2231); // @[AWSVggWrapper.scala 63:110]
  assign _T_2233 = queueIOOut_io_deq_bits[3215:3200]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_55 = $signed(_T_2233); // @[AWSVggWrapper.scala 63:110]
  assign _T_2235 = queueIOOut_io_deq_bits[3231:3216]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_54 = $signed(_T_2235); // @[AWSVggWrapper.scala 63:110]
  assign _T_2237 = queueIOOut_io_deq_bits[3247:3232]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_53 = $signed(_T_2237); // @[AWSVggWrapper.scala 63:110]
  assign _T_2239 = queueIOOut_io_deq_bits[3263:3248]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_52 = $signed(_T_2239); // @[AWSVggWrapper.scala 63:110]
  assign _T_2241 = queueIOOut_io_deq_bits[3279:3264]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_51 = $signed(_T_2241); // @[AWSVggWrapper.scala 63:110]
  assign _T_2243 = queueIOOut_io_deq_bits[3295:3280]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_50 = $signed(_T_2243); // @[AWSVggWrapper.scala 63:110]
  assign _T_2245 = queueIOOut_io_deq_bits[3311:3296]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_49 = $signed(_T_2245); // @[AWSVggWrapper.scala 63:110]
  assign _T_2247 = queueIOOut_io_deq_bits[3327:3312]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_48 = $signed(_T_2247); // @[AWSVggWrapper.scala 63:110]
  assign _T_2249 = queueIOOut_io_deq_bits[3343:3328]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_47 = $signed(_T_2249); // @[AWSVggWrapper.scala 63:110]
  assign _T_2251 = queueIOOut_io_deq_bits[3359:3344]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_46 = $signed(_T_2251); // @[AWSVggWrapper.scala 63:110]
  assign _T_2253 = queueIOOut_io_deq_bits[3375:3360]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_45 = $signed(_T_2253); // @[AWSVggWrapper.scala 63:110]
  assign _T_2255 = queueIOOut_io_deq_bits[3391:3376]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_44 = $signed(_T_2255); // @[AWSVggWrapper.scala 63:110]
  assign _T_2257 = queueIOOut_io_deq_bits[3407:3392]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_43 = $signed(_T_2257); // @[AWSVggWrapper.scala 63:110]
  assign _T_2259 = queueIOOut_io_deq_bits[3423:3408]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_42 = $signed(_T_2259); // @[AWSVggWrapper.scala 63:110]
  assign _T_2261 = queueIOOut_io_deq_bits[3439:3424]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_41 = $signed(_T_2261); // @[AWSVggWrapper.scala 63:110]
  assign _T_2263 = queueIOOut_io_deq_bits[3455:3440]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_40 = $signed(_T_2263); // @[AWSVggWrapper.scala 63:110]
  assign _T_2265 = queueIOOut_io_deq_bits[3471:3456]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_39 = $signed(_T_2265); // @[AWSVggWrapper.scala 63:110]
  assign _T_2267 = queueIOOut_io_deq_bits[3487:3472]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_38 = $signed(_T_2267); // @[AWSVggWrapper.scala 63:110]
  assign _T_2269 = queueIOOut_io_deq_bits[3503:3488]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_37 = $signed(_T_2269); // @[AWSVggWrapper.scala 63:110]
  assign _T_2271 = queueIOOut_io_deq_bits[3519:3504]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_36 = $signed(_T_2271); // @[AWSVggWrapper.scala 63:110]
  assign _T_2273 = queueIOOut_io_deq_bits[3535:3520]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_35 = $signed(_T_2273); // @[AWSVggWrapper.scala 63:110]
  assign _T_2275 = queueIOOut_io_deq_bits[3551:3536]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_34 = $signed(_T_2275); // @[AWSVggWrapper.scala 63:110]
  assign _T_2277 = queueIOOut_io_deq_bits[3567:3552]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_33 = $signed(_T_2277); // @[AWSVggWrapper.scala 63:110]
  assign _T_2279 = queueIOOut_io_deq_bits[3583:3568]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_32 = $signed(_T_2279); // @[AWSVggWrapper.scala 63:110]
  assign _T_2281 = queueIOOut_io_deq_bits[3599:3584]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_31 = $signed(_T_2281); // @[AWSVggWrapper.scala 63:110]
  assign _T_2283 = queueIOOut_io_deq_bits[3615:3600]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_30 = $signed(_T_2283); // @[AWSVggWrapper.scala 63:110]
  assign _T_2285 = queueIOOut_io_deq_bits[3631:3616]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_29 = $signed(_T_2285); // @[AWSVggWrapper.scala 63:110]
  assign _T_2287 = queueIOOut_io_deq_bits[3647:3632]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_28 = $signed(_T_2287); // @[AWSVggWrapper.scala 63:110]
  assign _T_2289 = queueIOOut_io_deq_bits[3663:3648]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_27 = $signed(_T_2289); // @[AWSVggWrapper.scala 63:110]
  assign _T_2291 = queueIOOut_io_deq_bits[3679:3664]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_26 = $signed(_T_2291); // @[AWSVggWrapper.scala 63:110]
  assign _T_2293 = queueIOOut_io_deq_bits[3695:3680]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_25 = $signed(_T_2293); // @[AWSVggWrapper.scala 63:110]
  assign _T_2295 = queueIOOut_io_deq_bits[3711:3696]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_24 = $signed(_T_2295); // @[AWSVggWrapper.scala 63:110]
  assign _T_2297 = queueIOOut_io_deq_bits[3727:3712]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_23 = $signed(_T_2297); // @[AWSVggWrapper.scala 63:110]
  assign _T_2299 = queueIOOut_io_deq_bits[3743:3728]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_22 = $signed(_T_2299); // @[AWSVggWrapper.scala 63:110]
  assign _T_2301 = queueIOOut_io_deq_bits[3759:3744]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_21 = $signed(_T_2301); // @[AWSVggWrapper.scala 63:110]
  assign _T_2303 = queueIOOut_io_deq_bits[3775:3760]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_20 = $signed(_T_2303); // @[AWSVggWrapper.scala 63:110]
  assign _T_2305 = queueIOOut_io_deq_bits[3791:3776]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_19 = $signed(_T_2305); // @[AWSVggWrapper.scala 63:110]
  assign _T_2307 = queueIOOut_io_deq_bits[3807:3792]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_18 = $signed(_T_2307); // @[AWSVggWrapper.scala 63:110]
  assign _T_2309 = queueIOOut_io_deq_bits[3823:3808]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_17 = $signed(_T_2309); // @[AWSVggWrapper.scala 63:110]
  assign _T_2311 = queueIOOut_io_deq_bits[3839:3824]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_16 = $signed(_T_2311); // @[AWSVggWrapper.scala 63:110]
  assign _T_2313 = queueIOOut_io_deq_bits[3855:3840]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_15 = $signed(_T_2313); // @[AWSVggWrapper.scala 63:110]
  assign _T_2315 = queueIOOut_io_deq_bits[3871:3856]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_14 = $signed(_T_2315); // @[AWSVggWrapper.scala 63:110]
  assign _T_2317 = queueIOOut_io_deq_bits[3887:3872]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_13 = $signed(_T_2317); // @[AWSVggWrapper.scala 63:110]
  assign _T_2319 = queueIOOut_io_deq_bits[3903:3888]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_12 = $signed(_T_2319); // @[AWSVggWrapper.scala 63:110]
  assign _T_2321 = queueIOOut_io_deq_bits[3919:3904]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_11 = $signed(_T_2321); // @[AWSVggWrapper.scala 63:110]
  assign _T_2323 = queueIOOut_io_deq_bits[3935:3920]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_10 = $signed(_T_2323); // @[AWSVggWrapper.scala 63:110]
  assign _T_2325 = queueIOOut_io_deq_bits[3951:3936]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_9 = $signed(_T_2325); // @[AWSVggWrapper.scala 63:110]
  assign _T_2327 = queueIOOut_io_deq_bits[3967:3952]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_8 = $signed(_T_2327); // @[AWSVggWrapper.scala 63:110]
  assign _T_2329 = queueIOOut_io_deq_bits[3983:3968]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_7 = $signed(_T_2329); // @[AWSVggWrapper.scala 63:110]
  assign _T_2331 = queueIOOut_io_deq_bits[3999:3984]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_6 = $signed(_T_2331); // @[AWSVggWrapper.scala 63:110]
  assign _T_2333 = queueIOOut_io_deq_bits[4015:4000]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_5 = $signed(_T_2333); // @[AWSVggWrapper.scala 63:110]
  assign _T_2335 = queueIOOut_io_deq_bits[4031:4016]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_4 = $signed(_T_2335); // @[AWSVggWrapper.scala 63:110]
  assign _T_2337 = queueIOOut_io_deq_bits[4047:4032]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_3 = $signed(_T_2337); // @[AWSVggWrapper.scala 63:110]
  assign _T_2339 = queueIOOut_io_deq_bits[4063:4048]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_2 = $signed(_T_2339); // @[AWSVggWrapper.scala 63:110]
  assign _T_2341 = queueIOOut_io_deq_bits[4079:4064]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_1 = $signed(_T_2341); // @[AWSVggWrapper.scala 63:110]
  assign _T_2343 = queueIOOut_io_deq_bits[4095:4080]; // @[AWSVggWrapper.scala 63:67]
  assign sintOut_0 = $signed(_T_2343); // @[AWSVggWrapper.scala 63:110]
  assign queueIOIn_ready = queueIOOut_io_enq_ready; // @[AWSVggWrapper.scala 53:23]
  assign queueIOIn_valid = vgg_io_dataOut_valid; // @[AWSVggWrapper.scala 53:23]
  assign io_dataIn_ready = vgg_io_dataIn_ready;
  assign io_dataOut_valid = muxLyr_io_dataOut_valid;
  assign io_dataOut_bits_0 = muxLyr_io_dataOut_bits_0;
  assign io_dataOut_bits_1 = muxLyr_io_dataOut_bits_1;
  assign io_dataOut_bits_2 = muxLyr_io_dataOut_bits_2;
  assign io_dataOut_bits_3 = muxLyr_io_dataOut_bits_3;
  assign vgg_clock = clock;
  assign vgg_reset = reset;
  assign vgg_io_dataIn_valid = io_dataIn_valid;
  assign vgg_io_dataIn_bits_0 = io_dataIn_bits_0;
  assign vgg_io_dataIn_bits_1 = io_dataIn_bits_1;
  assign vgg_io_dataIn_bits_2 = io_dataIn_bits_2;
  assign vgg_io_dataOut_ready = queueIOIn_ready;
  assign queueIOOut_clock = clock;
  assign queueIOOut_reset = reset;
  assign queueIOOut_io_enq_valid = queueIOIn_valid;
  assign queueIOOut_io_enq_bits = dataInAsUInt;
  assign queueIOOut_io_deq_ready = muxLyr_io_dataIn_ready;
  assign muxLyr_clock = clock;
  assign muxLyr_reset = reset;
  assign muxLyr_io_dataIn_valid = queueIOOut_io_deq_valid;
  assign muxLyr_io_dataIn_bits_0 = sintOut_0;
  assign muxLyr_io_dataIn_bits_1 = sintOut_1;
  assign muxLyr_io_dataIn_bits_2 = sintOut_2;
  assign muxLyr_io_dataIn_bits_3 = sintOut_3;
  assign muxLyr_io_dataIn_bits_4 = sintOut_4;
  assign muxLyr_io_dataIn_bits_5 = sintOut_5;
  assign muxLyr_io_dataIn_bits_6 = sintOut_6;
  assign muxLyr_io_dataIn_bits_7 = sintOut_7;
  assign muxLyr_io_dataIn_bits_8 = sintOut_8;
  assign muxLyr_io_dataIn_bits_9 = sintOut_9;
  assign muxLyr_io_dataIn_bits_10 = sintOut_10;
  assign muxLyr_io_dataIn_bits_11 = sintOut_11;
  assign muxLyr_io_dataIn_bits_12 = sintOut_12;
  assign muxLyr_io_dataIn_bits_13 = sintOut_13;
  assign muxLyr_io_dataIn_bits_14 = sintOut_14;
  assign muxLyr_io_dataIn_bits_15 = sintOut_15;
  assign muxLyr_io_dataIn_bits_16 = sintOut_16;
  assign muxLyr_io_dataIn_bits_17 = sintOut_17;
  assign muxLyr_io_dataIn_bits_18 = sintOut_18;
  assign muxLyr_io_dataIn_bits_19 = sintOut_19;
  assign muxLyr_io_dataIn_bits_20 = sintOut_20;
  assign muxLyr_io_dataIn_bits_21 = sintOut_21;
  assign muxLyr_io_dataIn_bits_22 = sintOut_22;
  assign muxLyr_io_dataIn_bits_23 = sintOut_23;
  assign muxLyr_io_dataIn_bits_24 = sintOut_24;
  assign muxLyr_io_dataIn_bits_25 = sintOut_25;
  assign muxLyr_io_dataIn_bits_26 = sintOut_26;
  assign muxLyr_io_dataIn_bits_27 = sintOut_27;
  assign muxLyr_io_dataIn_bits_28 = sintOut_28;
  assign muxLyr_io_dataIn_bits_29 = sintOut_29;
  assign muxLyr_io_dataIn_bits_30 = sintOut_30;
  assign muxLyr_io_dataIn_bits_31 = sintOut_31;
  assign muxLyr_io_dataIn_bits_32 = sintOut_32;
  assign muxLyr_io_dataIn_bits_33 = sintOut_33;
  assign muxLyr_io_dataIn_bits_34 = sintOut_34;
  assign muxLyr_io_dataIn_bits_35 = sintOut_35;
  assign muxLyr_io_dataIn_bits_36 = sintOut_36;
  assign muxLyr_io_dataIn_bits_37 = sintOut_37;
  assign muxLyr_io_dataIn_bits_38 = sintOut_38;
  assign muxLyr_io_dataIn_bits_39 = sintOut_39;
  assign muxLyr_io_dataIn_bits_40 = sintOut_40;
  assign muxLyr_io_dataIn_bits_41 = sintOut_41;
  assign muxLyr_io_dataIn_bits_42 = sintOut_42;
  assign muxLyr_io_dataIn_bits_43 = sintOut_43;
  assign muxLyr_io_dataIn_bits_44 = sintOut_44;
  assign muxLyr_io_dataIn_bits_45 = sintOut_45;
  assign muxLyr_io_dataIn_bits_46 = sintOut_46;
  assign muxLyr_io_dataIn_bits_47 = sintOut_47;
  assign muxLyr_io_dataIn_bits_48 = sintOut_48;
  assign muxLyr_io_dataIn_bits_49 = sintOut_49;
  assign muxLyr_io_dataIn_bits_50 = sintOut_50;
  assign muxLyr_io_dataIn_bits_51 = sintOut_51;
  assign muxLyr_io_dataIn_bits_52 = sintOut_52;
  assign muxLyr_io_dataIn_bits_53 = sintOut_53;
  assign muxLyr_io_dataIn_bits_54 = sintOut_54;
  assign muxLyr_io_dataIn_bits_55 = sintOut_55;
  assign muxLyr_io_dataIn_bits_56 = sintOut_56;
  assign muxLyr_io_dataIn_bits_57 = sintOut_57;
  assign muxLyr_io_dataIn_bits_58 = sintOut_58;
  assign muxLyr_io_dataIn_bits_59 = sintOut_59;
  assign muxLyr_io_dataIn_bits_60 = sintOut_60;
  assign muxLyr_io_dataIn_bits_61 = sintOut_61;
  assign muxLyr_io_dataIn_bits_62 = sintOut_62;
  assign muxLyr_io_dataIn_bits_63 = sintOut_63;
  assign muxLyr_io_dataIn_bits_64 = sintOut_64;
  assign muxLyr_io_dataIn_bits_65 = sintOut_65;
  assign muxLyr_io_dataIn_bits_66 = sintOut_66;
  assign muxLyr_io_dataIn_bits_67 = sintOut_67;
  assign muxLyr_io_dataIn_bits_68 = sintOut_68;
  assign muxLyr_io_dataIn_bits_69 = sintOut_69;
  assign muxLyr_io_dataIn_bits_70 = sintOut_70;
  assign muxLyr_io_dataIn_bits_71 = sintOut_71;
  assign muxLyr_io_dataIn_bits_72 = sintOut_72;
  assign muxLyr_io_dataIn_bits_73 = sintOut_73;
  assign muxLyr_io_dataIn_bits_74 = sintOut_74;
  assign muxLyr_io_dataIn_bits_75 = sintOut_75;
  assign muxLyr_io_dataIn_bits_76 = sintOut_76;
  assign muxLyr_io_dataIn_bits_77 = sintOut_77;
  assign muxLyr_io_dataIn_bits_78 = sintOut_78;
  assign muxLyr_io_dataIn_bits_79 = sintOut_79;
  assign muxLyr_io_dataIn_bits_80 = sintOut_80;
  assign muxLyr_io_dataIn_bits_81 = sintOut_81;
  assign muxLyr_io_dataIn_bits_82 = sintOut_82;
  assign muxLyr_io_dataIn_bits_83 = sintOut_83;
  assign muxLyr_io_dataIn_bits_84 = sintOut_84;
  assign muxLyr_io_dataIn_bits_85 = sintOut_85;
  assign muxLyr_io_dataIn_bits_86 = sintOut_86;
  assign muxLyr_io_dataIn_bits_87 = sintOut_87;
  assign muxLyr_io_dataIn_bits_88 = sintOut_88;
  assign muxLyr_io_dataIn_bits_89 = sintOut_89;
  assign muxLyr_io_dataIn_bits_90 = sintOut_90;
  assign muxLyr_io_dataIn_bits_91 = sintOut_91;
  assign muxLyr_io_dataIn_bits_92 = sintOut_92;
  assign muxLyr_io_dataIn_bits_93 = sintOut_93;
  assign muxLyr_io_dataIn_bits_94 = sintOut_94;
  assign muxLyr_io_dataIn_bits_95 = sintOut_95;
  assign muxLyr_io_dataIn_bits_96 = sintOut_96;
  assign muxLyr_io_dataIn_bits_97 = sintOut_97;
  assign muxLyr_io_dataIn_bits_98 = sintOut_98;
  assign muxLyr_io_dataIn_bits_99 = sintOut_99;
  assign muxLyr_io_dataIn_bits_100 = sintOut_100;
  assign muxLyr_io_dataIn_bits_101 = sintOut_101;
  assign muxLyr_io_dataIn_bits_102 = sintOut_102;
  assign muxLyr_io_dataIn_bits_103 = sintOut_103;
  assign muxLyr_io_dataIn_bits_104 = sintOut_104;
  assign muxLyr_io_dataIn_bits_105 = sintOut_105;
  assign muxLyr_io_dataIn_bits_106 = sintOut_106;
  assign muxLyr_io_dataIn_bits_107 = sintOut_107;
  assign muxLyr_io_dataIn_bits_108 = sintOut_108;
  assign muxLyr_io_dataIn_bits_109 = sintOut_109;
  assign muxLyr_io_dataIn_bits_110 = sintOut_110;
  assign muxLyr_io_dataIn_bits_111 = sintOut_111;
  assign muxLyr_io_dataIn_bits_112 = sintOut_112;
  assign muxLyr_io_dataIn_bits_113 = sintOut_113;
  assign muxLyr_io_dataIn_bits_114 = sintOut_114;
  assign muxLyr_io_dataIn_bits_115 = sintOut_115;
  assign muxLyr_io_dataIn_bits_116 = sintOut_116;
  assign muxLyr_io_dataIn_bits_117 = sintOut_117;
  assign muxLyr_io_dataIn_bits_118 = sintOut_118;
  assign muxLyr_io_dataIn_bits_119 = sintOut_119;
  assign muxLyr_io_dataIn_bits_120 = sintOut_120;
  assign muxLyr_io_dataIn_bits_121 = sintOut_121;
  assign muxLyr_io_dataIn_bits_122 = sintOut_122;
  assign muxLyr_io_dataIn_bits_123 = sintOut_123;
  assign muxLyr_io_dataIn_bits_124 = sintOut_124;
  assign muxLyr_io_dataIn_bits_125 = sintOut_125;
  assign muxLyr_io_dataIn_bits_126 = sintOut_126;
  assign muxLyr_io_dataIn_bits_127 = sintOut_127;
  assign muxLyr_io_dataIn_bits_128 = sintOut_128;
  assign muxLyr_io_dataIn_bits_129 = sintOut_129;
  assign muxLyr_io_dataIn_bits_130 = sintOut_130;
  assign muxLyr_io_dataIn_bits_131 = sintOut_131;
  assign muxLyr_io_dataIn_bits_132 = sintOut_132;
  assign muxLyr_io_dataIn_bits_133 = sintOut_133;
  assign muxLyr_io_dataIn_bits_134 = sintOut_134;
  assign muxLyr_io_dataIn_bits_135 = sintOut_135;
  assign muxLyr_io_dataIn_bits_136 = sintOut_136;
  assign muxLyr_io_dataIn_bits_137 = sintOut_137;
  assign muxLyr_io_dataIn_bits_138 = sintOut_138;
  assign muxLyr_io_dataIn_bits_139 = sintOut_139;
  assign muxLyr_io_dataIn_bits_140 = sintOut_140;
  assign muxLyr_io_dataIn_bits_141 = sintOut_141;
  assign muxLyr_io_dataIn_bits_142 = sintOut_142;
  assign muxLyr_io_dataIn_bits_143 = sintOut_143;
  assign muxLyr_io_dataIn_bits_144 = sintOut_144;
  assign muxLyr_io_dataIn_bits_145 = sintOut_145;
  assign muxLyr_io_dataIn_bits_146 = sintOut_146;
  assign muxLyr_io_dataIn_bits_147 = sintOut_147;
  assign muxLyr_io_dataIn_bits_148 = sintOut_148;
  assign muxLyr_io_dataIn_bits_149 = sintOut_149;
  assign muxLyr_io_dataIn_bits_150 = sintOut_150;
  assign muxLyr_io_dataIn_bits_151 = sintOut_151;
  assign muxLyr_io_dataIn_bits_152 = sintOut_152;
  assign muxLyr_io_dataIn_bits_153 = sintOut_153;
  assign muxLyr_io_dataIn_bits_154 = sintOut_154;
  assign muxLyr_io_dataIn_bits_155 = sintOut_155;
  assign muxLyr_io_dataIn_bits_156 = sintOut_156;
  assign muxLyr_io_dataIn_bits_157 = sintOut_157;
  assign muxLyr_io_dataIn_bits_158 = sintOut_158;
  assign muxLyr_io_dataIn_bits_159 = sintOut_159;
  assign muxLyr_io_dataIn_bits_160 = sintOut_160;
  assign muxLyr_io_dataIn_bits_161 = sintOut_161;
  assign muxLyr_io_dataIn_bits_162 = sintOut_162;
  assign muxLyr_io_dataIn_bits_163 = sintOut_163;
  assign muxLyr_io_dataIn_bits_164 = sintOut_164;
  assign muxLyr_io_dataIn_bits_165 = sintOut_165;
  assign muxLyr_io_dataIn_bits_166 = sintOut_166;
  assign muxLyr_io_dataIn_bits_167 = sintOut_167;
  assign muxLyr_io_dataIn_bits_168 = sintOut_168;
  assign muxLyr_io_dataIn_bits_169 = sintOut_169;
  assign muxLyr_io_dataIn_bits_170 = sintOut_170;
  assign muxLyr_io_dataIn_bits_171 = sintOut_171;
  assign muxLyr_io_dataIn_bits_172 = sintOut_172;
  assign muxLyr_io_dataIn_bits_173 = sintOut_173;
  assign muxLyr_io_dataIn_bits_174 = sintOut_174;
  assign muxLyr_io_dataIn_bits_175 = sintOut_175;
  assign muxLyr_io_dataIn_bits_176 = sintOut_176;
  assign muxLyr_io_dataIn_bits_177 = sintOut_177;
  assign muxLyr_io_dataIn_bits_178 = sintOut_178;
  assign muxLyr_io_dataIn_bits_179 = sintOut_179;
  assign muxLyr_io_dataIn_bits_180 = sintOut_180;
  assign muxLyr_io_dataIn_bits_181 = sintOut_181;
  assign muxLyr_io_dataIn_bits_182 = sintOut_182;
  assign muxLyr_io_dataIn_bits_183 = sintOut_183;
  assign muxLyr_io_dataIn_bits_184 = sintOut_184;
  assign muxLyr_io_dataIn_bits_185 = sintOut_185;
  assign muxLyr_io_dataIn_bits_186 = sintOut_186;
  assign muxLyr_io_dataIn_bits_187 = sintOut_187;
  assign muxLyr_io_dataIn_bits_188 = sintOut_188;
  assign muxLyr_io_dataIn_bits_189 = sintOut_189;
  assign muxLyr_io_dataIn_bits_190 = sintOut_190;
  assign muxLyr_io_dataIn_bits_191 = sintOut_191;
  assign muxLyr_io_dataIn_bits_192 = sintOut_192;
  assign muxLyr_io_dataIn_bits_193 = sintOut_193;
  assign muxLyr_io_dataIn_bits_194 = sintOut_194;
  assign muxLyr_io_dataIn_bits_195 = sintOut_195;
  assign muxLyr_io_dataIn_bits_196 = sintOut_196;
  assign muxLyr_io_dataIn_bits_197 = sintOut_197;
  assign muxLyr_io_dataIn_bits_198 = sintOut_198;
  assign muxLyr_io_dataIn_bits_199 = sintOut_199;
  assign muxLyr_io_dataIn_bits_200 = sintOut_200;
  assign muxLyr_io_dataIn_bits_201 = sintOut_201;
  assign muxLyr_io_dataIn_bits_202 = sintOut_202;
  assign muxLyr_io_dataIn_bits_203 = sintOut_203;
  assign muxLyr_io_dataIn_bits_204 = sintOut_204;
  assign muxLyr_io_dataIn_bits_205 = sintOut_205;
  assign muxLyr_io_dataIn_bits_206 = sintOut_206;
  assign muxLyr_io_dataIn_bits_207 = sintOut_207;
  assign muxLyr_io_dataIn_bits_208 = sintOut_208;
  assign muxLyr_io_dataIn_bits_209 = sintOut_209;
  assign muxLyr_io_dataIn_bits_210 = sintOut_210;
  assign muxLyr_io_dataIn_bits_211 = sintOut_211;
  assign muxLyr_io_dataIn_bits_212 = sintOut_212;
  assign muxLyr_io_dataIn_bits_213 = sintOut_213;
  assign muxLyr_io_dataIn_bits_214 = sintOut_214;
  assign muxLyr_io_dataIn_bits_215 = sintOut_215;
  assign muxLyr_io_dataIn_bits_216 = sintOut_216;
  assign muxLyr_io_dataIn_bits_217 = sintOut_217;
  assign muxLyr_io_dataIn_bits_218 = sintOut_218;
  assign muxLyr_io_dataIn_bits_219 = sintOut_219;
  assign muxLyr_io_dataIn_bits_220 = sintOut_220;
  assign muxLyr_io_dataIn_bits_221 = sintOut_221;
  assign muxLyr_io_dataIn_bits_222 = sintOut_222;
  assign muxLyr_io_dataIn_bits_223 = sintOut_223;
  assign muxLyr_io_dataIn_bits_224 = sintOut_224;
  assign muxLyr_io_dataIn_bits_225 = sintOut_225;
  assign muxLyr_io_dataIn_bits_226 = sintOut_226;
  assign muxLyr_io_dataIn_bits_227 = sintOut_227;
  assign muxLyr_io_dataIn_bits_228 = sintOut_228;
  assign muxLyr_io_dataIn_bits_229 = sintOut_229;
  assign muxLyr_io_dataIn_bits_230 = sintOut_230;
  assign muxLyr_io_dataIn_bits_231 = sintOut_231;
  assign muxLyr_io_dataIn_bits_232 = sintOut_232;
  assign muxLyr_io_dataIn_bits_233 = sintOut_233;
  assign muxLyr_io_dataIn_bits_234 = sintOut_234;
  assign muxLyr_io_dataIn_bits_235 = sintOut_235;
  assign muxLyr_io_dataIn_bits_236 = sintOut_236;
  assign muxLyr_io_dataIn_bits_237 = sintOut_237;
  assign muxLyr_io_dataIn_bits_238 = sintOut_238;
  assign muxLyr_io_dataIn_bits_239 = sintOut_239;
  assign muxLyr_io_dataIn_bits_240 = sintOut_240;
  assign muxLyr_io_dataIn_bits_241 = sintOut_241;
  assign muxLyr_io_dataIn_bits_242 = sintOut_242;
  assign muxLyr_io_dataIn_bits_243 = sintOut_243;
  assign muxLyr_io_dataIn_bits_244 = sintOut_244;
  assign muxLyr_io_dataIn_bits_245 = sintOut_245;
  assign muxLyr_io_dataIn_bits_246 = sintOut_246;
  assign muxLyr_io_dataIn_bits_247 = sintOut_247;
  assign muxLyr_io_dataIn_bits_248 = sintOut_248;
  assign muxLyr_io_dataIn_bits_249 = sintOut_249;
  assign muxLyr_io_dataIn_bits_250 = sintOut_250;
  assign muxLyr_io_dataIn_bits_251 = sintOut_251;
  assign muxLyr_io_dataIn_bits_252 = sintOut_252;
  assign muxLyr_io_dataIn_bits_253 = sintOut_253;
  assign muxLyr_io_dataIn_bits_254 = sintOut_254;
  assign muxLyr_io_dataIn_bits_255 = sintOut_255;
endmodule
