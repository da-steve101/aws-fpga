module MuxLayer(
  input         clock,
  input         reset,
  output        io_dataIn_ready,
  input         io_dataIn_valid,
  input  [15:0] io_dataIn_bits_0,
  input  [15:0] io_dataIn_bits_1,
  input  [15:0] io_dataIn_bits_2,
  input  [15:0] io_dataIn_bits_3,
  input  [15:0] io_dataIn_bits_4,
  input  [15:0] io_dataIn_bits_5,
  input  [15:0] io_dataIn_bits_6,
  input  [15:0] io_dataIn_bits_7,
  input  [15:0] io_dataIn_bits_8,
  input  [15:0] io_dataIn_bits_9,
  input  [15:0] io_dataIn_bits_10,
  input  [15:0] io_dataIn_bits_11,
  input  [15:0] io_dataIn_bits_12,
  input  [15:0] io_dataIn_bits_13,
  input  [15:0] io_dataIn_bits_14,
  input  [15:0] io_dataIn_bits_15,
  input  [15:0] io_dataIn_bits_16,
  input  [15:0] io_dataIn_bits_17,
  input  [15:0] io_dataIn_bits_18,
  input  [15:0] io_dataIn_bits_19,
  input  [15:0] io_dataIn_bits_20,
  input  [15:0] io_dataIn_bits_21,
  input  [15:0] io_dataIn_bits_22,
  input  [15:0] io_dataIn_bits_23,
  input  [15:0] io_dataIn_bits_24,
  input  [15:0] io_dataIn_bits_25,
  input  [15:0] io_dataIn_bits_26,
  input  [15:0] io_dataIn_bits_27,
  input  [15:0] io_dataIn_bits_28,
  input  [15:0] io_dataIn_bits_29,
  input  [15:0] io_dataIn_bits_30,
  input  [15:0] io_dataIn_bits_31,
  input  [15:0] io_dataIn_bits_32,
  input  [15:0] io_dataIn_bits_33,
  input  [15:0] io_dataIn_bits_34,
  input  [15:0] io_dataIn_bits_35,
  input  [15:0] io_dataIn_bits_36,
  input  [15:0] io_dataIn_bits_37,
  input  [15:0] io_dataIn_bits_38,
  input  [15:0] io_dataIn_bits_39,
  input  [15:0] io_dataIn_bits_40,
  input  [15:0] io_dataIn_bits_41,
  input  [15:0] io_dataIn_bits_42,
  input  [15:0] io_dataIn_bits_43,
  input  [15:0] io_dataIn_bits_44,
  input  [15:0] io_dataIn_bits_45,
  input  [15:0] io_dataIn_bits_46,
  input  [15:0] io_dataIn_bits_47,
  input  [15:0] io_dataIn_bits_48,
  input  [15:0] io_dataIn_bits_49,
  input  [15:0] io_dataIn_bits_50,
  input  [15:0] io_dataIn_bits_51,
  input  [15:0] io_dataIn_bits_52,
  input  [15:0] io_dataIn_bits_53,
  input  [15:0] io_dataIn_bits_54,
  input  [15:0] io_dataIn_bits_55,
  input  [15:0] io_dataIn_bits_56,
  input  [15:0] io_dataIn_bits_57,
  input  [15:0] io_dataIn_bits_58,
  input  [15:0] io_dataIn_bits_59,
  input  [15:0] io_dataIn_bits_60,
  input  [15:0] io_dataIn_bits_61,
  input  [15:0] io_dataIn_bits_62,
  input  [15:0] io_dataIn_bits_63,
  input  [15:0] io_dataIn_bits_64,
  input  [15:0] io_dataIn_bits_65,
  input  [15:0] io_dataIn_bits_66,
  input  [15:0] io_dataIn_bits_67,
  input  [15:0] io_dataIn_bits_68,
  input  [15:0] io_dataIn_bits_69,
  input  [15:0] io_dataIn_bits_70,
  input  [15:0] io_dataIn_bits_71,
  input  [15:0] io_dataIn_bits_72,
  input  [15:0] io_dataIn_bits_73,
  input  [15:0] io_dataIn_bits_74,
  input  [15:0] io_dataIn_bits_75,
  input  [15:0] io_dataIn_bits_76,
  input  [15:0] io_dataIn_bits_77,
  input  [15:0] io_dataIn_bits_78,
  input  [15:0] io_dataIn_bits_79,
  input  [15:0] io_dataIn_bits_80,
  input  [15:0] io_dataIn_bits_81,
  input  [15:0] io_dataIn_bits_82,
  input  [15:0] io_dataIn_bits_83,
  input  [15:0] io_dataIn_bits_84,
  input  [15:0] io_dataIn_bits_85,
  input  [15:0] io_dataIn_bits_86,
  input  [15:0] io_dataIn_bits_87,
  input  [15:0] io_dataIn_bits_88,
  input  [15:0] io_dataIn_bits_89,
  input  [15:0] io_dataIn_bits_90,
  input  [15:0] io_dataIn_bits_91,
  input  [15:0] io_dataIn_bits_92,
  input  [15:0] io_dataIn_bits_93,
  input  [15:0] io_dataIn_bits_94,
  input  [15:0] io_dataIn_bits_95,
  input  [15:0] io_dataIn_bits_96,
  input  [15:0] io_dataIn_bits_97,
  input  [15:0] io_dataIn_bits_98,
  input  [15:0] io_dataIn_bits_99,
  input  [15:0] io_dataIn_bits_100,
  input  [15:0] io_dataIn_bits_101,
  input  [15:0] io_dataIn_bits_102,
  input  [15:0] io_dataIn_bits_103,
  input  [15:0] io_dataIn_bits_104,
  input  [15:0] io_dataIn_bits_105,
  input  [15:0] io_dataIn_bits_106,
  input  [15:0] io_dataIn_bits_107,
  input  [15:0] io_dataIn_bits_108,
  input  [15:0] io_dataIn_bits_109,
  input  [15:0] io_dataIn_bits_110,
  input  [15:0] io_dataIn_bits_111,
  input  [15:0] io_dataIn_bits_112,
  input  [15:0] io_dataIn_bits_113,
  input  [15:0] io_dataIn_bits_114,
  input  [15:0] io_dataIn_bits_115,
  input  [15:0] io_dataIn_bits_116,
  input  [15:0] io_dataIn_bits_117,
  input  [15:0] io_dataIn_bits_118,
  input  [15:0] io_dataIn_bits_119,
  input  [15:0] io_dataIn_bits_120,
  input  [15:0] io_dataIn_bits_121,
  input  [15:0] io_dataIn_bits_122,
  input  [15:0] io_dataIn_bits_123,
  input  [15:0] io_dataIn_bits_124,
  input  [15:0] io_dataIn_bits_125,
  input  [15:0] io_dataIn_bits_126,
  input  [15:0] io_dataIn_bits_127,
  input  [15:0] io_dataIn_bits_128,
  input  [15:0] io_dataIn_bits_129,
  input  [15:0] io_dataIn_bits_130,
  input  [15:0] io_dataIn_bits_131,
  input  [15:0] io_dataIn_bits_132,
  input  [15:0] io_dataIn_bits_133,
  input  [15:0] io_dataIn_bits_134,
  input  [15:0] io_dataIn_bits_135,
  input  [15:0] io_dataIn_bits_136,
  input  [15:0] io_dataIn_bits_137,
  input  [15:0] io_dataIn_bits_138,
  input  [15:0] io_dataIn_bits_139,
  input  [15:0] io_dataIn_bits_140,
  input  [15:0] io_dataIn_bits_141,
  input  [15:0] io_dataIn_bits_142,
  input  [15:0] io_dataIn_bits_143,
  input  [15:0] io_dataIn_bits_144,
  input  [15:0] io_dataIn_bits_145,
  input  [15:0] io_dataIn_bits_146,
  input  [15:0] io_dataIn_bits_147,
  input  [15:0] io_dataIn_bits_148,
  input  [15:0] io_dataIn_bits_149,
  input  [15:0] io_dataIn_bits_150,
  input  [15:0] io_dataIn_bits_151,
  input  [15:0] io_dataIn_bits_152,
  input  [15:0] io_dataIn_bits_153,
  input  [15:0] io_dataIn_bits_154,
  input  [15:0] io_dataIn_bits_155,
  input  [15:0] io_dataIn_bits_156,
  input  [15:0] io_dataIn_bits_157,
  input  [15:0] io_dataIn_bits_158,
  input  [15:0] io_dataIn_bits_159,
  input  [15:0] io_dataIn_bits_160,
  input  [15:0] io_dataIn_bits_161,
  input  [15:0] io_dataIn_bits_162,
  input  [15:0] io_dataIn_bits_163,
  input  [15:0] io_dataIn_bits_164,
  input  [15:0] io_dataIn_bits_165,
  input  [15:0] io_dataIn_bits_166,
  input  [15:0] io_dataIn_bits_167,
  input  [15:0] io_dataIn_bits_168,
  input  [15:0] io_dataIn_bits_169,
  input  [15:0] io_dataIn_bits_170,
  input  [15:0] io_dataIn_bits_171,
  input  [15:0] io_dataIn_bits_172,
  input  [15:0] io_dataIn_bits_173,
  input  [15:0] io_dataIn_bits_174,
  input  [15:0] io_dataIn_bits_175,
  input  [15:0] io_dataIn_bits_176,
  input  [15:0] io_dataIn_bits_177,
  input  [15:0] io_dataIn_bits_178,
  input  [15:0] io_dataIn_bits_179,
  input  [15:0] io_dataIn_bits_180,
  input  [15:0] io_dataIn_bits_181,
  input  [15:0] io_dataIn_bits_182,
  input  [15:0] io_dataIn_bits_183,
  input  [15:0] io_dataIn_bits_184,
  input  [15:0] io_dataIn_bits_185,
  input  [15:0] io_dataIn_bits_186,
  input  [15:0] io_dataIn_bits_187,
  input  [15:0] io_dataIn_bits_188,
  input  [15:0] io_dataIn_bits_189,
  input  [15:0] io_dataIn_bits_190,
  input  [15:0] io_dataIn_bits_191,
  input  [15:0] io_dataIn_bits_192,
  input  [15:0] io_dataIn_bits_193,
  input  [15:0] io_dataIn_bits_194,
  input  [15:0] io_dataIn_bits_195,
  input  [15:0] io_dataIn_bits_196,
  input  [15:0] io_dataIn_bits_197,
  input  [15:0] io_dataIn_bits_198,
  input  [15:0] io_dataIn_bits_199,
  input  [15:0] io_dataIn_bits_200,
  input  [15:0] io_dataIn_bits_201,
  input  [15:0] io_dataIn_bits_202,
  input  [15:0] io_dataIn_bits_203,
  input  [15:0] io_dataIn_bits_204,
  input  [15:0] io_dataIn_bits_205,
  input  [15:0] io_dataIn_bits_206,
  input  [15:0] io_dataIn_bits_207,
  input  [15:0] io_dataIn_bits_208,
  input  [15:0] io_dataIn_bits_209,
  input  [15:0] io_dataIn_bits_210,
  input  [15:0] io_dataIn_bits_211,
  input  [15:0] io_dataIn_bits_212,
  input  [15:0] io_dataIn_bits_213,
  input  [15:0] io_dataIn_bits_214,
  input  [15:0] io_dataIn_bits_215,
  input  [15:0] io_dataIn_bits_216,
  input  [15:0] io_dataIn_bits_217,
  input  [15:0] io_dataIn_bits_218,
  input  [15:0] io_dataIn_bits_219,
  input  [15:0] io_dataIn_bits_220,
  input  [15:0] io_dataIn_bits_221,
  input  [15:0] io_dataIn_bits_222,
  input  [15:0] io_dataIn_bits_223,
  input  [15:0] io_dataIn_bits_224,
  input  [15:0] io_dataIn_bits_225,
  input  [15:0] io_dataIn_bits_226,
  input  [15:0] io_dataIn_bits_227,
  input  [15:0] io_dataIn_bits_228,
  input  [15:0] io_dataIn_bits_229,
  input  [15:0] io_dataIn_bits_230,
  input  [15:0] io_dataIn_bits_231,
  input  [15:0] io_dataIn_bits_232,
  input  [15:0] io_dataIn_bits_233,
  input  [15:0] io_dataIn_bits_234,
  input  [15:0] io_dataIn_bits_235,
  input  [15:0] io_dataIn_bits_236,
  input  [15:0] io_dataIn_bits_237,
  input  [15:0] io_dataIn_bits_238,
  input  [15:0] io_dataIn_bits_239,
  input  [15:0] io_dataIn_bits_240,
  input  [15:0] io_dataIn_bits_241,
  input  [15:0] io_dataIn_bits_242,
  input  [15:0] io_dataIn_bits_243,
  input  [15:0] io_dataIn_bits_244,
  input  [15:0] io_dataIn_bits_245,
  input  [15:0] io_dataIn_bits_246,
  input  [15:0] io_dataIn_bits_247,
  input  [15:0] io_dataIn_bits_248,
  input  [15:0] io_dataIn_bits_249,
  input  [15:0] io_dataIn_bits_250,
  input  [15:0] io_dataIn_bits_251,
  input  [15:0] io_dataIn_bits_252,
  input  [15:0] io_dataIn_bits_253,
  input  [15:0] io_dataIn_bits_254,
  input  [15:0] io_dataIn_bits_255,
  output        io_dataOut_valid,
  output [15:0] io_dataOut_bits_0,
  output [15:0] io_dataOut_bits_1,
  output [15:0] io_dataOut_bits_2,
  output [15:0] io_dataOut_bits_3
);
  reg  rdyReg; // @[MuxLayer.scala 14:23]
  reg [31:0] _RAND_0;
  reg [5:0] cntr; // @[MuxLayer.scala 17:21]
  reg [31:0] _RAND_1;
  reg [15:0] buffers_0_0_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_2;
  reg [15:0] buffers_0_0_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_3;
  reg [15:0] buffers_0_0_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_4;
  reg [15:0] buffers_0_0_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_5;
  reg [15:0] buffers_0_1_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_6;
  reg [15:0] buffers_0_1_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_7;
  reg [15:0] buffers_0_1_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_8;
  reg [15:0] buffers_0_1_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_9;
  reg [15:0] buffers_0_2_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_10;
  reg [15:0] buffers_0_2_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_11;
  reg [15:0] buffers_0_2_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_12;
  reg [15:0] buffers_0_2_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_13;
  reg [15:0] buffers_0_3_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_14;
  reg [15:0] buffers_0_3_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_15;
  reg [15:0] buffers_0_3_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_16;
  reg [15:0] buffers_0_3_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_17;
  reg [15:0] buffers_0_4_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_18;
  reg [15:0] buffers_0_4_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_19;
  reg [15:0] buffers_0_4_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_20;
  reg [15:0] buffers_0_4_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_21;
  reg [15:0] buffers_0_5_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_22;
  reg [15:0] buffers_0_5_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_23;
  reg [15:0] buffers_0_5_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_24;
  reg [15:0] buffers_0_5_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_25;
  reg [15:0] buffers_0_6_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_26;
  reg [15:0] buffers_0_6_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_27;
  reg [15:0] buffers_0_6_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_28;
  reg [15:0] buffers_0_6_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_29;
  reg [15:0] buffers_0_7_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_30;
  reg [15:0] buffers_0_7_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_31;
  reg [15:0] buffers_0_7_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_32;
  reg [15:0] buffers_0_7_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_33;
  reg [15:0] buffers_0_8_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_34;
  reg [15:0] buffers_0_8_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_35;
  reg [15:0] buffers_0_8_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_36;
  reg [15:0] buffers_0_8_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_37;
  reg [15:0] buffers_0_9_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_38;
  reg [15:0] buffers_0_9_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_39;
  reg [15:0] buffers_0_9_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_40;
  reg [15:0] buffers_0_9_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_41;
  reg [15:0] buffers_0_10_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_42;
  reg [15:0] buffers_0_10_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_43;
  reg [15:0] buffers_0_10_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_44;
  reg [15:0] buffers_0_10_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_45;
  reg [15:0] buffers_0_11_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_46;
  reg [15:0] buffers_0_11_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_47;
  reg [15:0] buffers_0_11_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_48;
  reg [15:0] buffers_0_11_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_49;
  reg [15:0] buffers_0_12_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_50;
  reg [15:0] buffers_0_12_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_51;
  reg [15:0] buffers_0_12_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_52;
  reg [15:0] buffers_0_12_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_53;
  reg [15:0] buffers_0_13_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_54;
  reg [15:0] buffers_0_13_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_55;
  reg [15:0] buffers_0_13_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_56;
  reg [15:0] buffers_0_13_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_57;
  reg [15:0] buffers_0_14_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_58;
  reg [15:0] buffers_0_14_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_59;
  reg [15:0] buffers_0_14_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_60;
  reg [15:0] buffers_0_14_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_61;
  reg [15:0] buffers_0_15_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_62;
  reg [15:0] buffers_0_15_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_63;
  reg [15:0] buffers_0_15_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_64;
  reg [15:0] buffers_0_15_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_65;
  reg [15:0] buffers_0_16_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_66;
  reg [15:0] buffers_0_16_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_67;
  reg [15:0] buffers_0_16_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_68;
  reg [15:0] buffers_0_16_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_69;
  reg [15:0] buffers_0_17_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_70;
  reg [15:0] buffers_0_17_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_71;
  reg [15:0] buffers_0_17_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_72;
  reg [15:0] buffers_0_17_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_73;
  reg [15:0] buffers_0_18_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_74;
  reg [15:0] buffers_0_18_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_75;
  reg [15:0] buffers_0_18_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_76;
  reg [15:0] buffers_0_18_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_77;
  reg [15:0] buffers_0_19_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_78;
  reg [15:0] buffers_0_19_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_79;
  reg [15:0] buffers_0_19_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_80;
  reg [15:0] buffers_0_19_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_81;
  reg [15:0] buffers_0_20_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_82;
  reg [15:0] buffers_0_20_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_83;
  reg [15:0] buffers_0_20_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_84;
  reg [15:0] buffers_0_20_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_85;
  reg [15:0] buffers_0_21_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_86;
  reg [15:0] buffers_0_21_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_87;
  reg [15:0] buffers_0_21_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_88;
  reg [15:0] buffers_0_21_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_89;
  reg [15:0] buffers_0_22_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_90;
  reg [15:0] buffers_0_22_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_91;
  reg [15:0] buffers_0_22_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_92;
  reg [15:0] buffers_0_22_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_93;
  reg [15:0] buffers_0_23_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_94;
  reg [15:0] buffers_0_23_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_95;
  reg [15:0] buffers_0_23_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_96;
  reg [15:0] buffers_0_23_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_97;
  reg [15:0] buffers_0_24_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_98;
  reg [15:0] buffers_0_24_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_99;
  reg [15:0] buffers_0_24_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_100;
  reg [15:0] buffers_0_24_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_101;
  reg [15:0] buffers_0_25_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_102;
  reg [15:0] buffers_0_25_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_103;
  reg [15:0] buffers_0_25_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_104;
  reg [15:0] buffers_0_25_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_105;
  reg [15:0] buffers_0_26_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_106;
  reg [15:0] buffers_0_26_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_107;
  reg [15:0] buffers_0_26_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_108;
  reg [15:0] buffers_0_26_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_109;
  reg [15:0] buffers_0_27_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_110;
  reg [15:0] buffers_0_27_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_111;
  reg [15:0] buffers_0_27_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_112;
  reg [15:0] buffers_0_27_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_113;
  reg [15:0] buffers_0_28_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_114;
  reg [15:0] buffers_0_28_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_115;
  reg [15:0] buffers_0_28_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_116;
  reg [15:0] buffers_0_28_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_117;
  reg [15:0] buffers_0_29_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_118;
  reg [15:0] buffers_0_29_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_119;
  reg [15:0] buffers_0_29_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_120;
  reg [15:0] buffers_0_29_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_121;
  reg [15:0] buffers_0_30_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_122;
  reg [15:0] buffers_0_30_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_123;
  reg [15:0] buffers_0_30_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_124;
  reg [15:0] buffers_0_30_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_125;
  reg [15:0] buffers_0_31_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_126;
  reg [15:0] buffers_0_31_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_127;
  reg [15:0] buffers_0_31_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_128;
  reg [15:0] buffers_0_31_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_129;
  reg [15:0] buffers_0_32_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_130;
  reg [15:0] buffers_0_32_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_131;
  reg [15:0] buffers_0_32_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_132;
  reg [15:0] buffers_0_32_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_133;
  reg [15:0] buffers_0_33_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_134;
  reg [15:0] buffers_0_33_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_135;
  reg [15:0] buffers_0_33_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_136;
  reg [15:0] buffers_0_33_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_137;
  reg [15:0] buffers_0_34_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_138;
  reg [15:0] buffers_0_34_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_139;
  reg [15:0] buffers_0_34_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_140;
  reg [15:0] buffers_0_34_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_141;
  reg [15:0] buffers_0_35_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_142;
  reg [15:0] buffers_0_35_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_143;
  reg [15:0] buffers_0_35_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_144;
  reg [15:0] buffers_0_35_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_145;
  reg [15:0] buffers_0_36_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_146;
  reg [15:0] buffers_0_36_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_147;
  reg [15:0] buffers_0_36_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_148;
  reg [15:0] buffers_0_36_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_149;
  reg [15:0] buffers_0_37_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_150;
  reg [15:0] buffers_0_37_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_151;
  reg [15:0] buffers_0_37_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_152;
  reg [15:0] buffers_0_37_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_153;
  reg [15:0] buffers_0_38_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_154;
  reg [15:0] buffers_0_38_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_155;
  reg [15:0] buffers_0_38_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_156;
  reg [15:0] buffers_0_38_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_157;
  reg [15:0] buffers_0_39_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_158;
  reg [15:0] buffers_0_39_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_159;
  reg [15:0] buffers_0_39_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_160;
  reg [15:0] buffers_0_39_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_161;
  reg [15:0] buffers_0_40_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_162;
  reg [15:0] buffers_0_40_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_163;
  reg [15:0] buffers_0_40_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_164;
  reg [15:0] buffers_0_40_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_165;
  reg [15:0] buffers_0_41_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_166;
  reg [15:0] buffers_0_41_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_167;
  reg [15:0] buffers_0_41_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_168;
  reg [15:0] buffers_0_41_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_169;
  reg [15:0] buffers_0_42_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_170;
  reg [15:0] buffers_0_42_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_171;
  reg [15:0] buffers_0_42_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_172;
  reg [15:0] buffers_0_42_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_173;
  reg [15:0] buffers_0_43_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_174;
  reg [15:0] buffers_0_43_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_175;
  reg [15:0] buffers_0_43_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_176;
  reg [15:0] buffers_0_43_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_177;
  reg [15:0] buffers_0_44_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_178;
  reg [15:0] buffers_0_44_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_179;
  reg [15:0] buffers_0_44_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_180;
  reg [15:0] buffers_0_44_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_181;
  reg [15:0] buffers_0_45_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_182;
  reg [15:0] buffers_0_45_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_183;
  reg [15:0] buffers_0_45_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_184;
  reg [15:0] buffers_0_45_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_185;
  reg [15:0] buffers_0_46_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_186;
  reg [15:0] buffers_0_46_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_187;
  reg [15:0] buffers_0_46_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_188;
  reg [15:0] buffers_0_46_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_189;
  reg [15:0] buffers_0_47_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_190;
  reg [15:0] buffers_0_47_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_191;
  reg [15:0] buffers_0_47_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_192;
  reg [15:0] buffers_0_47_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_193;
  reg [15:0] buffers_0_48_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_194;
  reg [15:0] buffers_0_48_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_195;
  reg [15:0] buffers_0_48_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_196;
  reg [15:0] buffers_0_48_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_197;
  reg [15:0] buffers_0_49_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_198;
  reg [15:0] buffers_0_49_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_199;
  reg [15:0] buffers_0_49_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_200;
  reg [15:0] buffers_0_49_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_201;
  reg [15:0] buffers_0_50_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_202;
  reg [15:0] buffers_0_50_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_203;
  reg [15:0] buffers_0_50_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_204;
  reg [15:0] buffers_0_50_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_205;
  reg [15:0] buffers_0_51_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_206;
  reg [15:0] buffers_0_51_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_207;
  reg [15:0] buffers_0_51_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_208;
  reg [15:0] buffers_0_51_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_209;
  reg [15:0] buffers_0_52_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_210;
  reg [15:0] buffers_0_52_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_211;
  reg [15:0] buffers_0_52_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_212;
  reg [15:0] buffers_0_52_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_213;
  reg [15:0] buffers_0_53_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_214;
  reg [15:0] buffers_0_53_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_215;
  reg [15:0] buffers_0_53_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_216;
  reg [15:0] buffers_0_53_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_217;
  reg [15:0] buffers_0_54_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_218;
  reg [15:0] buffers_0_54_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_219;
  reg [15:0] buffers_0_54_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_220;
  reg [15:0] buffers_0_54_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_221;
  reg [15:0] buffers_0_55_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_222;
  reg [15:0] buffers_0_55_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_223;
  reg [15:0] buffers_0_55_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_224;
  reg [15:0] buffers_0_55_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_225;
  reg [15:0] buffers_0_56_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_226;
  reg [15:0] buffers_0_56_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_227;
  reg [15:0] buffers_0_56_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_228;
  reg [15:0] buffers_0_56_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_229;
  reg [15:0] buffers_0_57_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_230;
  reg [15:0] buffers_0_57_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_231;
  reg [15:0] buffers_0_57_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_232;
  reg [15:0] buffers_0_57_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_233;
  reg [15:0] buffers_0_58_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_234;
  reg [15:0] buffers_0_58_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_235;
  reg [15:0] buffers_0_58_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_236;
  reg [15:0] buffers_0_58_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_237;
  reg [15:0] buffers_0_59_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_238;
  reg [15:0] buffers_0_59_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_239;
  reg [15:0] buffers_0_59_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_240;
  reg [15:0] buffers_0_59_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_241;
  reg [15:0] buffers_0_60_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_242;
  reg [15:0] buffers_0_60_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_243;
  reg [15:0] buffers_0_60_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_244;
  reg [15:0] buffers_0_60_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_245;
  reg [15:0] buffers_0_61_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_246;
  reg [15:0] buffers_0_61_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_247;
  reg [15:0] buffers_0_61_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_248;
  reg [15:0] buffers_0_61_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_249;
  reg [15:0] buffers_0_62_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_250;
  reg [15:0] buffers_0_62_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_251;
  reg [15:0] buffers_0_62_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_252;
  reg [15:0] buffers_0_62_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_253;
  reg [15:0] buffers_0_63_0; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_254;
  reg [15:0] buffers_0_63_1; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_255;
  reg [15:0] buffers_0_63_2; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_256;
  reg [15:0] buffers_0_63_3; // @[MuxLayer.scala 18:45]
  reg [31:0] _RAND_257;
  reg [1:0] cntrs_0; // @[Reg.scala 11:16]
  reg [31:0] _RAND_258;
  reg [1:0] _T_1071; // @[Reg.scala 11:16]
  reg [31:0] _RAND_259;
  reg [1:0] cntrs_1; // @[Reg.scala 11:16]
  reg [31:0] _RAND_260;
  reg [1:0] _T_1076; // @[Reg.scala 11:16]
  reg [31:0] _RAND_261;
  reg [1:0] _T_1078; // @[Reg.scala 11:16]
  reg [31:0] _RAND_262;
  reg [1:0] cntrs_2; // @[Reg.scala 11:16]
  reg [31:0] _RAND_263;
  reg [15:0] buffers_1_0_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_264;
  reg [15:0] buffers_1_0_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_265;
  reg [15:0] buffers_1_0_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_266;
  reg [15:0] buffers_1_0_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_267;
  reg [15:0] buffers_1_1_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_268;
  reg [15:0] buffers_1_1_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_269;
  reg [15:0] buffers_1_1_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_270;
  reg [15:0] buffers_1_1_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_271;
  reg [15:0] buffers_1_2_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_272;
  reg [15:0] buffers_1_2_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_273;
  reg [15:0] buffers_1_2_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_274;
  reg [15:0] buffers_1_2_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_275;
  reg [15:0] buffers_1_3_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_276;
  reg [15:0] buffers_1_3_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_277;
  reg [15:0] buffers_1_3_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_278;
  reg [15:0] buffers_1_3_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_279;
  reg [15:0] buffers_1_4_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_280;
  reg [15:0] buffers_1_4_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_281;
  reg [15:0] buffers_1_4_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_282;
  reg [15:0] buffers_1_4_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_283;
  reg [15:0] buffers_1_5_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_284;
  reg [15:0] buffers_1_5_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_285;
  reg [15:0] buffers_1_5_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_286;
  reg [15:0] buffers_1_5_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_287;
  reg [15:0] buffers_1_6_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_288;
  reg [15:0] buffers_1_6_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_289;
  reg [15:0] buffers_1_6_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_290;
  reg [15:0] buffers_1_6_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_291;
  reg [15:0] buffers_1_7_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_292;
  reg [15:0] buffers_1_7_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_293;
  reg [15:0] buffers_1_7_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_294;
  reg [15:0] buffers_1_7_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_295;
  reg [15:0] buffers_1_8_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_296;
  reg [15:0] buffers_1_8_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_297;
  reg [15:0] buffers_1_8_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_298;
  reg [15:0] buffers_1_8_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_299;
  reg [15:0] buffers_1_9_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_300;
  reg [15:0] buffers_1_9_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_301;
  reg [15:0] buffers_1_9_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_302;
  reg [15:0] buffers_1_9_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_303;
  reg [15:0] buffers_1_10_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_304;
  reg [15:0] buffers_1_10_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_305;
  reg [15:0] buffers_1_10_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_306;
  reg [15:0] buffers_1_10_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_307;
  reg [15:0] buffers_1_11_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_308;
  reg [15:0] buffers_1_11_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_309;
  reg [15:0] buffers_1_11_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_310;
  reg [15:0] buffers_1_11_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_311;
  reg [15:0] buffers_1_12_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_312;
  reg [15:0] buffers_1_12_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_313;
  reg [15:0] buffers_1_12_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_314;
  reg [15:0] buffers_1_12_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_315;
  reg [15:0] buffers_1_13_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_316;
  reg [15:0] buffers_1_13_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_317;
  reg [15:0] buffers_1_13_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_318;
  reg [15:0] buffers_1_13_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_319;
  reg [15:0] buffers_1_14_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_320;
  reg [15:0] buffers_1_14_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_321;
  reg [15:0] buffers_1_14_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_322;
  reg [15:0] buffers_1_14_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_323;
  reg [15:0] buffers_1_15_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_324;
  reg [15:0] buffers_1_15_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_325;
  reg [15:0] buffers_1_15_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_326;
  reg [15:0] buffers_1_15_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_327;
  reg [15:0] buffers_2_0_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_328;
  reg [15:0] buffers_2_0_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_329;
  reg [15:0] buffers_2_0_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_330;
  reg [15:0] buffers_2_0_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_331;
  reg [15:0] buffers_2_1_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_332;
  reg [15:0] buffers_2_1_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_333;
  reg [15:0] buffers_2_1_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_334;
  reg [15:0] buffers_2_1_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_335;
  reg [15:0] buffers_2_2_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_336;
  reg [15:0] buffers_2_2_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_337;
  reg [15:0] buffers_2_2_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_338;
  reg [15:0] buffers_2_2_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_339;
  reg [15:0] buffers_2_3_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_340;
  reg [15:0] buffers_2_3_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_341;
  reg [15:0] buffers_2_3_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_342;
  reg [15:0] buffers_2_3_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_343;
  reg [15:0] buffers_3_0_0; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_344;
  reg [15:0] buffers_3_0_1; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_345;
  reg [15:0] buffers_3_0_2; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_346;
  reg [15:0] buffers_3_0_3; // @[MuxLayer.scala 59:14]
  reg [31:0] _RAND_347;
  reg  _T_1988; // @[Reg.scala 19:20]
  reg [31:0] _RAND_348;
  reg  _T_1990; // @[Reg.scala 19:20]
  reg [31:0] _RAND_349;
  reg  vld; // @[Reg.scala 19:20]
  reg [31:0] _RAND_350;
  reg  lastVld; // @[MuxLayer.scala 66:24]
  reg [31:0] _RAND_351;
  wire  _T_1052; // @[MuxLayer.scala 19:15]
  wire [6:0] _T_1054; // @[MuxLayer.scala 20:18]
  wire [5:0] _T_1055; // @[MuxLayer.scala 20:18]
  wire [5:0] _GEN_0; // @[MuxLayer.scala 19:23]
  wire  _T_1057; // @[MuxLayer.scala 22:34]
  wire  _T_1058; // @[MuxLayer.scala 22:26]
  wire [5:0] _GEN_1; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_2; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_3; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_4; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_5; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_6; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_7; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_8; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_9; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_10; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_11; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_12; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_13; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_14; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_15; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_16; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_17; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_18; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_19; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_20; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_21; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_22; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_23; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_24; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_25; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_26; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_27; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_28; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_29; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_30; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_31; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_32; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_33; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_34; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_35; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_36; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_37; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_38; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_39; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_40; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_41; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_42; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_43; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_44; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_45; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_46; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_47; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_48; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_49; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_50; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_51; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_52; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_53; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_54; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_55; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_56; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_57; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_58; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_59; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_60; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_61; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_62; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_63; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_64; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_65; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_66; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_67; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_68; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_69; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_70; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_71; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_72; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_73; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_74; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_75; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_76; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_77; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_78; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_79; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_80; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_81; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_82; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_83; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_84; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_85; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_86; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_87; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_88; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_89; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_90; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_91; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_92; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_93; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_94; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_95; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_96; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_97; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_98; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_99; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_100; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_101; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_102; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_103; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_104; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_105; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_106; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_107; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_108; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_109; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_110; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_111; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_112; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_113; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_114; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_115; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_116; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_117; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_118; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_119; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_120; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_121; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_122; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_123; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_124; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_125; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_126; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_127; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_128; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_129; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_130; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_131; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_132; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_133; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_134; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_135; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_136; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_137; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_138; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_139; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_140; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_141; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_142; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_143; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_144; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_145; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_146; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_147; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_148; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_149; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_150; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_151; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_152; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_153; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_154; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_155; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_156; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_157; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_158; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_159; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_160; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_161; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_162; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_163; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_164; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_165; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_166; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_167; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_168; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_169; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_170; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_171; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_172; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_173; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_174; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_175; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_176; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_177; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_178; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_179; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_180; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_181; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_182; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_183; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_184; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_185; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_186; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_187; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_188; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_189; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_190; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_191; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_192; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_193; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_194; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_195; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_196; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_197; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_198; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_199; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_200; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_201; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_202; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_203; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_204; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_205; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_206; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_207; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_208; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_209; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_210; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_211; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_212; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_213; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_214; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_215; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_216; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_217; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_218; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_219; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_220; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_221; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_222; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_223; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_224; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_225; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_226; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_227; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_228; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_229; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_230; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_231; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_232; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_233; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_234; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_235; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_236; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_237; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_238; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_239; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_240; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_241; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_242; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_243; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_244; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_245; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_246; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_247; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_248; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_249; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_250; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_251; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_252; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_253; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_254; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_255; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_256; // @[MuxLayer.scala 22:44]
  wire [15:0] _GEN_257; // @[MuxLayer.scala 22:44]
  wire  _T_1061; // @[MuxLayer.scala 29:15]
  wire  _GEN_258; // @[MuxLayer.scala 29:36]
  wire  _T_1063; // @[MuxLayer.scala 32:26]
  wire  _GEN_259; // @[MuxLayer.scala 32:38]
  wire [1:0] _T_1065; // @[MuxLayer.scala 45:19]
  wire [1:0] _T_1068; // @[MuxLayer.scala 45:19]
  wire [1:0] _T_1073; // @[MuxLayer.scala 45:19]
  wire  _T_1090; // @[MuxLayer.scala 55:25]
  wire [15:0] _GEN_266; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_267; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_268; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_269; // @[MuxLayer.scala 55:35]
  wire  _T_1092; // @[MuxLayer.scala 55:25]
  wire [15:0] _GEN_270; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_271; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_272; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_273; // @[MuxLayer.scala 55:35]
  wire  _T_1094; // @[MuxLayer.scala 55:25]
  wire [15:0] _GEN_274; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_275; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_276; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_277; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_278; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_279; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_280; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_281; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_282; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_283; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_284; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_285; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_286; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_287; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_288; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_289; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_290; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_291; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_292; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_293; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_294; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_295; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_296; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_297; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_298; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_299; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_300; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_301; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_302; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_303; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_304; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_305; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_306; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_307; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_308; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_309; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_310; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_311; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_312; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_313; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_314; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_315; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_316; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_317; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_318; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_319; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_320; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_321; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_322; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_323; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_324; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_325; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_326; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_327; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_328; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_329; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_330; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_331; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_332; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_333; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_334; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_335; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_336; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_337; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_338; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_339; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_340; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_341; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_342; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_343; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_344; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_345; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_346; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_347; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_348; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_349; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_350; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_351; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_352; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_353; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_354; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_355; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_356; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_357; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_358; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_359; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_360; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_361; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_362; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_363; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_364; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_365; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_366; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_367; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_368; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_369; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_370; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_371; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_372; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_373; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_374; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_375; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_376; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_377; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_378; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_379; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_380; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_381; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_382; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_383; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_384; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_385; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_386; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_387; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_388; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_389; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_390; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_391; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_392; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_393; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_394; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_395; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_396; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_397; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_398; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_399; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_400; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_401; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_402; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_403; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_404; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_405; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_406; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_407; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_408; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_409; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_410; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_411; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_412; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_413; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_414; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_415; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_416; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_417; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_418; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_419; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_420; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_421; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_422; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_423; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_424; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_425; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_426; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_427; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_428; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_429; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_430; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_431; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_432; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_433; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_434; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_435; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_436; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_437; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_438; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_439; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_440; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_441; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_442; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_443; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_444; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_445; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_446; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_447; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_448; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_449; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_450; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_451; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_452; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_453; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_454; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_455; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_456; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_457; // @[MuxLayer.scala 55:35]
  wire  _T_1778; // @[MuxLayer.scala 55:25]
  wire [15:0] _GEN_458; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_459; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_460; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_461; // @[MuxLayer.scala 55:35]
  wire  _T_1780; // @[MuxLayer.scala 55:25]
  wire [15:0] _GEN_462; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_463; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_464; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_465; // @[MuxLayer.scala 55:35]
  wire  _T_1782; // @[MuxLayer.scala 55:25]
  wire [15:0] _GEN_466; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_467; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_468; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_469; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_470; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_471; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_472; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_473; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_474; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_475; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_476; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_477; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_478; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_479; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_480; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_481; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_482; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_483; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_484; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_485; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_486; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_487; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_488; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_489; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_490; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_491; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_492; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_493; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_494; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_495; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_496; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_497; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_498; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_499; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_500; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_501; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_502; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_503; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_504; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_505; // @[MuxLayer.scala 55:35]
  wire  _T_1950; // @[MuxLayer.scala 55:25]
  wire [15:0] _GEN_506; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_507; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_508; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_509; // @[MuxLayer.scala 55:35]
  wire  _T_1952; // @[MuxLayer.scala 55:25]
  wire [15:0] _GEN_510; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_511; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_512; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_513; // @[MuxLayer.scala 55:35]
  wire  _T_1954; // @[MuxLayer.scala 55:25]
  wire [15:0] _GEN_514; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_515; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_516; // @[MuxLayer.scala 55:35]
  wire [15:0] _GEN_517; // @[MuxLayer.scala 55:35]
  wire  _T_1994; // @[MuxLayer.scala 68:27]
  assign _T_1052 = cntr > 6'h0; // @[MuxLayer.scala 19:15]
  assign _T_1054 = cntr + 6'h1; // @[MuxLayer.scala 20:18]
  assign _T_1055 = _T_1054[5:0]; // @[MuxLayer.scala 20:18]
  assign _GEN_0 = _T_1052 ? _T_1055 : cntr; // @[MuxLayer.scala 19:23]
  assign _T_1057 = cntr == 6'h0; // @[MuxLayer.scala 22:34]
  assign _T_1058 = io_dataIn_valid & _T_1057; // @[MuxLayer.scala 22:26]
  assign _GEN_1 = _T_1058 ? 6'h1 : _GEN_0; // @[MuxLayer.scala 22:44]
  assign _GEN_2 = _T_1058 ? $signed(io_dataIn_bits_0) : $signed(buffers_0_0_0); // @[MuxLayer.scala 22:44]
  assign _GEN_3 = _T_1058 ? $signed(io_dataIn_bits_1) : $signed(buffers_0_0_1); // @[MuxLayer.scala 22:44]
  assign _GEN_4 = _T_1058 ? $signed(io_dataIn_bits_2) : $signed(buffers_0_0_2); // @[MuxLayer.scala 22:44]
  assign _GEN_5 = _T_1058 ? $signed(io_dataIn_bits_3) : $signed(buffers_0_0_3); // @[MuxLayer.scala 22:44]
  assign _GEN_6 = _T_1058 ? $signed(io_dataIn_bits_4) : $signed(buffers_0_1_0); // @[MuxLayer.scala 22:44]
  assign _GEN_7 = _T_1058 ? $signed(io_dataIn_bits_5) : $signed(buffers_0_1_1); // @[MuxLayer.scala 22:44]
  assign _GEN_8 = _T_1058 ? $signed(io_dataIn_bits_6) : $signed(buffers_0_1_2); // @[MuxLayer.scala 22:44]
  assign _GEN_9 = _T_1058 ? $signed(io_dataIn_bits_7) : $signed(buffers_0_1_3); // @[MuxLayer.scala 22:44]
  assign _GEN_10 = _T_1058 ? $signed(io_dataIn_bits_8) : $signed(buffers_0_2_0); // @[MuxLayer.scala 22:44]
  assign _GEN_11 = _T_1058 ? $signed(io_dataIn_bits_9) : $signed(buffers_0_2_1); // @[MuxLayer.scala 22:44]
  assign _GEN_12 = _T_1058 ? $signed(io_dataIn_bits_10) : $signed(buffers_0_2_2); // @[MuxLayer.scala 22:44]
  assign _GEN_13 = _T_1058 ? $signed(io_dataIn_bits_11) : $signed(buffers_0_2_3); // @[MuxLayer.scala 22:44]
  assign _GEN_14 = _T_1058 ? $signed(io_dataIn_bits_12) : $signed(buffers_0_3_0); // @[MuxLayer.scala 22:44]
  assign _GEN_15 = _T_1058 ? $signed(io_dataIn_bits_13) : $signed(buffers_0_3_1); // @[MuxLayer.scala 22:44]
  assign _GEN_16 = _T_1058 ? $signed(io_dataIn_bits_14) : $signed(buffers_0_3_2); // @[MuxLayer.scala 22:44]
  assign _GEN_17 = _T_1058 ? $signed(io_dataIn_bits_15) : $signed(buffers_0_3_3); // @[MuxLayer.scala 22:44]
  assign _GEN_18 = _T_1058 ? $signed(io_dataIn_bits_16) : $signed(buffers_0_4_0); // @[MuxLayer.scala 22:44]
  assign _GEN_19 = _T_1058 ? $signed(io_dataIn_bits_17) : $signed(buffers_0_4_1); // @[MuxLayer.scala 22:44]
  assign _GEN_20 = _T_1058 ? $signed(io_dataIn_bits_18) : $signed(buffers_0_4_2); // @[MuxLayer.scala 22:44]
  assign _GEN_21 = _T_1058 ? $signed(io_dataIn_bits_19) : $signed(buffers_0_4_3); // @[MuxLayer.scala 22:44]
  assign _GEN_22 = _T_1058 ? $signed(io_dataIn_bits_20) : $signed(buffers_0_5_0); // @[MuxLayer.scala 22:44]
  assign _GEN_23 = _T_1058 ? $signed(io_dataIn_bits_21) : $signed(buffers_0_5_1); // @[MuxLayer.scala 22:44]
  assign _GEN_24 = _T_1058 ? $signed(io_dataIn_bits_22) : $signed(buffers_0_5_2); // @[MuxLayer.scala 22:44]
  assign _GEN_25 = _T_1058 ? $signed(io_dataIn_bits_23) : $signed(buffers_0_5_3); // @[MuxLayer.scala 22:44]
  assign _GEN_26 = _T_1058 ? $signed(io_dataIn_bits_24) : $signed(buffers_0_6_0); // @[MuxLayer.scala 22:44]
  assign _GEN_27 = _T_1058 ? $signed(io_dataIn_bits_25) : $signed(buffers_0_6_1); // @[MuxLayer.scala 22:44]
  assign _GEN_28 = _T_1058 ? $signed(io_dataIn_bits_26) : $signed(buffers_0_6_2); // @[MuxLayer.scala 22:44]
  assign _GEN_29 = _T_1058 ? $signed(io_dataIn_bits_27) : $signed(buffers_0_6_3); // @[MuxLayer.scala 22:44]
  assign _GEN_30 = _T_1058 ? $signed(io_dataIn_bits_28) : $signed(buffers_0_7_0); // @[MuxLayer.scala 22:44]
  assign _GEN_31 = _T_1058 ? $signed(io_dataIn_bits_29) : $signed(buffers_0_7_1); // @[MuxLayer.scala 22:44]
  assign _GEN_32 = _T_1058 ? $signed(io_dataIn_bits_30) : $signed(buffers_0_7_2); // @[MuxLayer.scala 22:44]
  assign _GEN_33 = _T_1058 ? $signed(io_dataIn_bits_31) : $signed(buffers_0_7_3); // @[MuxLayer.scala 22:44]
  assign _GEN_34 = _T_1058 ? $signed(io_dataIn_bits_32) : $signed(buffers_0_8_0); // @[MuxLayer.scala 22:44]
  assign _GEN_35 = _T_1058 ? $signed(io_dataIn_bits_33) : $signed(buffers_0_8_1); // @[MuxLayer.scala 22:44]
  assign _GEN_36 = _T_1058 ? $signed(io_dataIn_bits_34) : $signed(buffers_0_8_2); // @[MuxLayer.scala 22:44]
  assign _GEN_37 = _T_1058 ? $signed(io_dataIn_bits_35) : $signed(buffers_0_8_3); // @[MuxLayer.scala 22:44]
  assign _GEN_38 = _T_1058 ? $signed(io_dataIn_bits_36) : $signed(buffers_0_9_0); // @[MuxLayer.scala 22:44]
  assign _GEN_39 = _T_1058 ? $signed(io_dataIn_bits_37) : $signed(buffers_0_9_1); // @[MuxLayer.scala 22:44]
  assign _GEN_40 = _T_1058 ? $signed(io_dataIn_bits_38) : $signed(buffers_0_9_2); // @[MuxLayer.scala 22:44]
  assign _GEN_41 = _T_1058 ? $signed(io_dataIn_bits_39) : $signed(buffers_0_9_3); // @[MuxLayer.scala 22:44]
  assign _GEN_42 = _T_1058 ? $signed(io_dataIn_bits_40) : $signed(buffers_0_10_0); // @[MuxLayer.scala 22:44]
  assign _GEN_43 = _T_1058 ? $signed(io_dataIn_bits_41) : $signed(buffers_0_10_1); // @[MuxLayer.scala 22:44]
  assign _GEN_44 = _T_1058 ? $signed(io_dataIn_bits_42) : $signed(buffers_0_10_2); // @[MuxLayer.scala 22:44]
  assign _GEN_45 = _T_1058 ? $signed(io_dataIn_bits_43) : $signed(buffers_0_10_3); // @[MuxLayer.scala 22:44]
  assign _GEN_46 = _T_1058 ? $signed(io_dataIn_bits_44) : $signed(buffers_0_11_0); // @[MuxLayer.scala 22:44]
  assign _GEN_47 = _T_1058 ? $signed(io_dataIn_bits_45) : $signed(buffers_0_11_1); // @[MuxLayer.scala 22:44]
  assign _GEN_48 = _T_1058 ? $signed(io_dataIn_bits_46) : $signed(buffers_0_11_2); // @[MuxLayer.scala 22:44]
  assign _GEN_49 = _T_1058 ? $signed(io_dataIn_bits_47) : $signed(buffers_0_11_3); // @[MuxLayer.scala 22:44]
  assign _GEN_50 = _T_1058 ? $signed(io_dataIn_bits_48) : $signed(buffers_0_12_0); // @[MuxLayer.scala 22:44]
  assign _GEN_51 = _T_1058 ? $signed(io_dataIn_bits_49) : $signed(buffers_0_12_1); // @[MuxLayer.scala 22:44]
  assign _GEN_52 = _T_1058 ? $signed(io_dataIn_bits_50) : $signed(buffers_0_12_2); // @[MuxLayer.scala 22:44]
  assign _GEN_53 = _T_1058 ? $signed(io_dataIn_bits_51) : $signed(buffers_0_12_3); // @[MuxLayer.scala 22:44]
  assign _GEN_54 = _T_1058 ? $signed(io_dataIn_bits_52) : $signed(buffers_0_13_0); // @[MuxLayer.scala 22:44]
  assign _GEN_55 = _T_1058 ? $signed(io_dataIn_bits_53) : $signed(buffers_0_13_1); // @[MuxLayer.scala 22:44]
  assign _GEN_56 = _T_1058 ? $signed(io_dataIn_bits_54) : $signed(buffers_0_13_2); // @[MuxLayer.scala 22:44]
  assign _GEN_57 = _T_1058 ? $signed(io_dataIn_bits_55) : $signed(buffers_0_13_3); // @[MuxLayer.scala 22:44]
  assign _GEN_58 = _T_1058 ? $signed(io_dataIn_bits_56) : $signed(buffers_0_14_0); // @[MuxLayer.scala 22:44]
  assign _GEN_59 = _T_1058 ? $signed(io_dataIn_bits_57) : $signed(buffers_0_14_1); // @[MuxLayer.scala 22:44]
  assign _GEN_60 = _T_1058 ? $signed(io_dataIn_bits_58) : $signed(buffers_0_14_2); // @[MuxLayer.scala 22:44]
  assign _GEN_61 = _T_1058 ? $signed(io_dataIn_bits_59) : $signed(buffers_0_14_3); // @[MuxLayer.scala 22:44]
  assign _GEN_62 = _T_1058 ? $signed(io_dataIn_bits_60) : $signed(buffers_0_15_0); // @[MuxLayer.scala 22:44]
  assign _GEN_63 = _T_1058 ? $signed(io_dataIn_bits_61) : $signed(buffers_0_15_1); // @[MuxLayer.scala 22:44]
  assign _GEN_64 = _T_1058 ? $signed(io_dataIn_bits_62) : $signed(buffers_0_15_2); // @[MuxLayer.scala 22:44]
  assign _GEN_65 = _T_1058 ? $signed(io_dataIn_bits_63) : $signed(buffers_0_15_3); // @[MuxLayer.scala 22:44]
  assign _GEN_66 = _T_1058 ? $signed(io_dataIn_bits_64) : $signed(buffers_0_16_0); // @[MuxLayer.scala 22:44]
  assign _GEN_67 = _T_1058 ? $signed(io_dataIn_bits_65) : $signed(buffers_0_16_1); // @[MuxLayer.scala 22:44]
  assign _GEN_68 = _T_1058 ? $signed(io_dataIn_bits_66) : $signed(buffers_0_16_2); // @[MuxLayer.scala 22:44]
  assign _GEN_69 = _T_1058 ? $signed(io_dataIn_bits_67) : $signed(buffers_0_16_3); // @[MuxLayer.scala 22:44]
  assign _GEN_70 = _T_1058 ? $signed(io_dataIn_bits_68) : $signed(buffers_0_17_0); // @[MuxLayer.scala 22:44]
  assign _GEN_71 = _T_1058 ? $signed(io_dataIn_bits_69) : $signed(buffers_0_17_1); // @[MuxLayer.scala 22:44]
  assign _GEN_72 = _T_1058 ? $signed(io_dataIn_bits_70) : $signed(buffers_0_17_2); // @[MuxLayer.scala 22:44]
  assign _GEN_73 = _T_1058 ? $signed(io_dataIn_bits_71) : $signed(buffers_0_17_3); // @[MuxLayer.scala 22:44]
  assign _GEN_74 = _T_1058 ? $signed(io_dataIn_bits_72) : $signed(buffers_0_18_0); // @[MuxLayer.scala 22:44]
  assign _GEN_75 = _T_1058 ? $signed(io_dataIn_bits_73) : $signed(buffers_0_18_1); // @[MuxLayer.scala 22:44]
  assign _GEN_76 = _T_1058 ? $signed(io_dataIn_bits_74) : $signed(buffers_0_18_2); // @[MuxLayer.scala 22:44]
  assign _GEN_77 = _T_1058 ? $signed(io_dataIn_bits_75) : $signed(buffers_0_18_3); // @[MuxLayer.scala 22:44]
  assign _GEN_78 = _T_1058 ? $signed(io_dataIn_bits_76) : $signed(buffers_0_19_0); // @[MuxLayer.scala 22:44]
  assign _GEN_79 = _T_1058 ? $signed(io_dataIn_bits_77) : $signed(buffers_0_19_1); // @[MuxLayer.scala 22:44]
  assign _GEN_80 = _T_1058 ? $signed(io_dataIn_bits_78) : $signed(buffers_0_19_2); // @[MuxLayer.scala 22:44]
  assign _GEN_81 = _T_1058 ? $signed(io_dataIn_bits_79) : $signed(buffers_0_19_3); // @[MuxLayer.scala 22:44]
  assign _GEN_82 = _T_1058 ? $signed(io_dataIn_bits_80) : $signed(buffers_0_20_0); // @[MuxLayer.scala 22:44]
  assign _GEN_83 = _T_1058 ? $signed(io_dataIn_bits_81) : $signed(buffers_0_20_1); // @[MuxLayer.scala 22:44]
  assign _GEN_84 = _T_1058 ? $signed(io_dataIn_bits_82) : $signed(buffers_0_20_2); // @[MuxLayer.scala 22:44]
  assign _GEN_85 = _T_1058 ? $signed(io_dataIn_bits_83) : $signed(buffers_0_20_3); // @[MuxLayer.scala 22:44]
  assign _GEN_86 = _T_1058 ? $signed(io_dataIn_bits_84) : $signed(buffers_0_21_0); // @[MuxLayer.scala 22:44]
  assign _GEN_87 = _T_1058 ? $signed(io_dataIn_bits_85) : $signed(buffers_0_21_1); // @[MuxLayer.scala 22:44]
  assign _GEN_88 = _T_1058 ? $signed(io_dataIn_bits_86) : $signed(buffers_0_21_2); // @[MuxLayer.scala 22:44]
  assign _GEN_89 = _T_1058 ? $signed(io_dataIn_bits_87) : $signed(buffers_0_21_3); // @[MuxLayer.scala 22:44]
  assign _GEN_90 = _T_1058 ? $signed(io_dataIn_bits_88) : $signed(buffers_0_22_0); // @[MuxLayer.scala 22:44]
  assign _GEN_91 = _T_1058 ? $signed(io_dataIn_bits_89) : $signed(buffers_0_22_1); // @[MuxLayer.scala 22:44]
  assign _GEN_92 = _T_1058 ? $signed(io_dataIn_bits_90) : $signed(buffers_0_22_2); // @[MuxLayer.scala 22:44]
  assign _GEN_93 = _T_1058 ? $signed(io_dataIn_bits_91) : $signed(buffers_0_22_3); // @[MuxLayer.scala 22:44]
  assign _GEN_94 = _T_1058 ? $signed(io_dataIn_bits_92) : $signed(buffers_0_23_0); // @[MuxLayer.scala 22:44]
  assign _GEN_95 = _T_1058 ? $signed(io_dataIn_bits_93) : $signed(buffers_0_23_1); // @[MuxLayer.scala 22:44]
  assign _GEN_96 = _T_1058 ? $signed(io_dataIn_bits_94) : $signed(buffers_0_23_2); // @[MuxLayer.scala 22:44]
  assign _GEN_97 = _T_1058 ? $signed(io_dataIn_bits_95) : $signed(buffers_0_23_3); // @[MuxLayer.scala 22:44]
  assign _GEN_98 = _T_1058 ? $signed(io_dataIn_bits_96) : $signed(buffers_0_24_0); // @[MuxLayer.scala 22:44]
  assign _GEN_99 = _T_1058 ? $signed(io_dataIn_bits_97) : $signed(buffers_0_24_1); // @[MuxLayer.scala 22:44]
  assign _GEN_100 = _T_1058 ? $signed(io_dataIn_bits_98) : $signed(buffers_0_24_2); // @[MuxLayer.scala 22:44]
  assign _GEN_101 = _T_1058 ? $signed(io_dataIn_bits_99) : $signed(buffers_0_24_3); // @[MuxLayer.scala 22:44]
  assign _GEN_102 = _T_1058 ? $signed(io_dataIn_bits_100) : $signed(buffers_0_25_0); // @[MuxLayer.scala 22:44]
  assign _GEN_103 = _T_1058 ? $signed(io_dataIn_bits_101) : $signed(buffers_0_25_1); // @[MuxLayer.scala 22:44]
  assign _GEN_104 = _T_1058 ? $signed(io_dataIn_bits_102) : $signed(buffers_0_25_2); // @[MuxLayer.scala 22:44]
  assign _GEN_105 = _T_1058 ? $signed(io_dataIn_bits_103) : $signed(buffers_0_25_3); // @[MuxLayer.scala 22:44]
  assign _GEN_106 = _T_1058 ? $signed(io_dataIn_bits_104) : $signed(buffers_0_26_0); // @[MuxLayer.scala 22:44]
  assign _GEN_107 = _T_1058 ? $signed(io_dataIn_bits_105) : $signed(buffers_0_26_1); // @[MuxLayer.scala 22:44]
  assign _GEN_108 = _T_1058 ? $signed(io_dataIn_bits_106) : $signed(buffers_0_26_2); // @[MuxLayer.scala 22:44]
  assign _GEN_109 = _T_1058 ? $signed(io_dataIn_bits_107) : $signed(buffers_0_26_3); // @[MuxLayer.scala 22:44]
  assign _GEN_110 = _T_1058 ? $signed(io_dataIn_bits_108) : $signed(buffers_0_27_0); // @[MuxLayer.scala 22:44]
  assign _GEN_111 = _T_1058 ? $signed(io_dataIn_bits_109) : $signed(buffers_0_27_1); // @[MuxLayer.scala 22:44]
  assign _GEN_112 = _T_1058 ? $signed(io_dataIn_bits_110) : $signed(buffers_0_27_2); // @[MuxLayer.scala 22:44]
  assign _GEN_113 = _T_1058 ? $signed(io_dataIn_bits_111) : $signed(buffers_0_27_3); // @[MuxLayer.scala 22:44]
  assign _GEN_114 = _T_1058 ? $signed(io_dataIn_bits_112) : $signed(buffers_0_28_0); // @[MuxLayer.scala 22:44]
  assign _GEN_115 = _T_1058 ? $signed(io_dataIn_bits_113) : $signed(buffers_0_28_1); // @[MuxLayer.scala 22:44]
  assign _GEN_116 = _T_1058 ? $signed(io_dataIn_bits_114) : $signed(buffers_0_28_2); // @[MuxLayer.scala 22:44]
  assign _GEN_117 = _T_1058 ? $signed(io_dataIn_bits_115) : $signed(buffers_0_28_3); // @[MuxLayer.scala 22:44]
  assign _GEN_118 = _T_1058 ? $signed(io_dataIn_bits_116) : $signed(buffers_0_29_0); // @[MuxLayer.scala 22:44]
  assign _GEN_119 = _T_1058 ? $signed(io_dataIn_bits_117) : $signed(buffers_0_29_1); // @[MuxLayer.scala 22:44]
  assign _GEN_120 = _T_1058 ? $signed(io_dataIn_bits_118) : $signed(buffers_0_29_2); // @[MuxLayer.scala 22:44]
  assign _GEN_121 = _T_1058 ? $signed(io_dataIn_bits_119) : $signed(buffers_0_29_3); // @[MuxLayer.scala 22:44]
  assign _GEN_122 = _T_1058 ? $signed(io_dataIn_bits_120) : $signed(buffers_0_30_0); // @[MuxLayer.scala 22:44]
  assign _GEN_123 = _T_1058 ? $signed(io_dataIn_bits_121) : $signed(buffers_0_30_1); // @[MuxLayer.scala 22:44]
  assign _GEN_124 = _T_1058 ? $signed(io_dataIn_bits_122) : $signed(buffers_0_30_2); // @[MuxLayer.scala 22:44]
  assign _GEN_125 = _T_1058 ? $signed(io_dataIn_bits_123) : $signed(buffers_0_30_3); // @[MuxLayer.scala 22:44]
  assign _GEN_126 = _T_1058 ? $signed(io_dataIn_bits_124) : $signed(buffers_0_31_0); // @[MuxLayer.scala 22:44]
  assign _GEN_127 = _T_1058 ? $signed(io_dataIn_bits_125) : $signed(buffers_0_31_1); // @[MuxLayer.scala 22:44]
  assign _GEN_128 = _T_1058 ? $signed(io_dataIn_bits_126) : $signed(buffers_0_31_2); // @[MuxLayer.scala 22:44]
  assign _GEN_129 = _T_1058 ? $signed(io_dataIn_bits_127) : $signed(buffers_0_31_3); // @[MuxLayer.scala 22:44]
  assign _GEN_130 = _T_1058 ? $signed(io_dataIn_bits_128) : $signed(buffers_0_32_0); // @[MuxLayer.scala 22:44]
  assign _GEN_131 = _T_1058 ? $signed(io_dataIn_bits_129) : $signed(buffers_0_32_1); // @[MuxLayer.scala 22:44]
  assign _GEN_132 = _T_1058 ? $signed(io_dataIn_bits_130) : $signed(buffers_0_32_2); // @[MuxLayer.scala 22:44]
  assign _GEN_133 = _T_1058 ? $signed(io_dataIn_bits_131) : $signed(buffers_0_32_3); // @[MuxLayer.scala 22:44]
  assign _GEN_134 = _T_1058 ? $signed(io_dataIn_bits_132) : $signed(buffers_0_33_0); // @[MuxLayer.scala 22:44]
  assign _GEN_135 = _T_1058 ? $signed(io_dataIn_bits_133) : $signed(buffers_0_33_1); // @[MuxLayer.scala 22:44]
  assign _GEN_136 = _T_1058 ? $signed(io_dataIn_bits_134) : $signed(buffers_0_33_2); // @[MuxLayer.scala 22:44]
  assign _GEN_137 = _T_1058 ? $signed(io_dataIn_bits_135) : $signed(buffers_0_33_3); // @[MuxLayer.scala 22:44]
  assign _GEN_138 = _T_1058 ? $signed(io_dataIn_bits_136) : $signed(buffers_0_34_0); // @[MuxLayer.scala 22:44]
  assign _GEN_139 = _T_1058 ? $signed(io_dataIn_bits_137) : $signed(buffers_0_34_1); // @[MuxLayer.scala 22:44]
  assign _GEN_140 = _T_1058 ? $signed(io_dataIn_bits_138) : $signed(buffers_0_34_2); // @[MuxLayer.scala 22:44]
  assign _GEN_141 = _T_1058 ? $signed(io_dataIn_bits_139) : $signed(buffers_0_34_3); // @[MuxLayer.scala 22:44]
  assign _GEN_142 = _T_1058 ? $signed(io_dataIn_bits_140) : $signed(buffers_0_35_0); // @[MuxLayer.scala 22:44]
  assign _GEN_143 = _T_1058 ? $signed(io_dataIn_bits_141) : $signed(buffers_0_35_1); // @[MuxLayer.scala 22:44]
  assign _GEN_144 = _T_1058 ? $signed(io_dataIn_bits_142) : $signed(buffers_0_35_2); // @[MuxLayer.scala 22:44]
  assign _GEN_145 = _T_1058 ? $signed(io_dataIn_bits_143) : $signed(buffers_0_35_3); // @[MuxLayer.scala 22:44]
  assign _GEN_146 = _T_1058 ? $signed(io_dataIn_bits_144) : $signed(buffers_0_36_0); // @[MuxLayer.scala 22:44]
  assign _GEN_147 = _T_1058 ? $signed(io_dataIn_bits_145) : $signed(buffers_0_36_1); // @[MuxLayer.scala 22:44]
  assign _GEN_148 = _T_1058 ? $signed(io_dataIn_bits_146) : $signed(buffers_0_36_2); // @[MuxLayer.scala 22:44]
  assign _GEN_149 = _T_1058 ? $signed(io_dataIn_bits_147) : $signed(buffers_0_36_3); // @[MuxLayer.scala 22:44]
  assign _GEN_150 = _T_1058 ? $signed(io_dataIn_bits_148) : $signed(buffers_0_37_0); // @[MuxLayer.scala 22:44]
  assign _GEN_151 = _T_1058 ? $signed(io_dataIn_bits_149) : $signed(buffers_0_37_1); // @[MuxLayer.scala 22:44]
  assign _GEN_152 = _T_1058 ? $signed(io_dataIn_bits_150) : $signed(buffers_0_37_2); // @[MuxLayer.scala 22:44]
  assign _GEN_153 = _T_1058 ? $signed(io_dataIn_bits_151) : $signed(buffers_0_37_3); // @[MuxLayer.scala 22:44]
  assign _GEN_154 = _T_1058 ? $signed(io_dataIn_bits_152) : $signed(buffers_0_38_0); // @[MuxLayer.scala 22:44]
  assign _GEN_155 = _T_1058 ? $signed(io_dataIn_bits_153) : $signed(buffers_0_38_1); // @[MuxLayer.scala 22:44]
  assign _GEN_156 = _T_1058 ? $signed(io_dataIn_bits_154) : $signed(buffers_0_38_2); // @[MuxLayer.scala 22:44]
  assign _GEN_157 = _T_1058 ? $signed(io_dataIn_bits_155) : $signed(buffers_0_38_3); // @[MuxLayer.scala 22:44]
  assign _GEN_158 = _T_1058 ? $signed(io_dataIn_bits_156) : $signed(buffers_0_39_0); // @[MuxLayer.scala 22:44]
  assign _GEN_159 = _T_1058 ? $signed(io_dataIn_bits_157) : $signed(buffers_0_39_1); // @[MuxLayer.scala 22:44]
  assign _GEN_160 = _T_1058 ? $signed(io_dataIn_bits_158) : $signed(buffers_0_39_2); // @[MuxLayer.scala 22:44]
  assign _GEN_161 = _T_1058 ? $signed(io_dataIn_bits_159) : $signed(buffers_0_39_3); // @[MuxLayer.scala 22:44]
  assign _GEN_162 = _T_1058 ? $signed(io_dataIn_bits_160) : $signed(buffers_0_40_0); // @[MuxLayer.scala 22:44]
  assign _GEN_163 = _T_1058 ? $signed(io_dataIn_bits_161) : $signed(buffers_0_40_1); // @[MuxLayer.scala 22:44]
  assign _GEN_164 = _T_1058 ? $signed(io_dataIn_bits_162) : $signed(buffers_0_40_2); // @[MuxLayer.scala 22:44]
  assign _GEN_165 = _T_1058 ? $signed(io_dataIn_bits_163) : $signed(buffers_0_40_3); // @[MuxLayer.scala 22:44]
  assign _GEN_166 = _T_1058 ? $signed(io_dataIn_bits_164) : $signed(buffers_0_41_0); // @[MuxLayer.scala 22:44]
  assign _GEN_167 = _T_1058 ? $signed(io_dataIn_bits_165) : $signed(buffers_0_41_1); // @[MuxLayer.scala 22:44]
  assign _GEN_168 = _T_1058 ? $signed(io_dataIn_bits_166) : $signed(buffers_0_41_2); // @[MuxLayer.scala 22:44]
  assign _GEN_169 = _T_1058 ? $signed(io_dataIn_bits_167) : $signed(buffers_0_41_3); // @[MuxLayer.scala 22:44]
  assign _GEN_170 = _T_1058 ? $signed(io_dataIn_bits_168) : $signed(buffers_0_42_0); // @[MuxLayer.scala 22:44]
  assign _GEN_171 = _T_1058 ? $signed(io_dataIn_bits_169) : $signed(buffers_0_42_1); // @[MuxLayer.scala 22:44]
  assign _GEN_172 = _T_1058 ? $signed(io_dataIn_bits_170) : $signed(buffers_0_42_2); // @[MuxLayer.scala 22:44]
  assign _GEN_173 = _T_1058 ? $signed(io_dataIn_bits_171) : $signed(buffers_0_42_3); // @[MuxLayer.scala 22:44]
  assign _GEN_174 = _T_1058 ? $signed(io_dataIn_bits_172) : $signed(buffers_0_43_0); // @[MuxLayer.scala 22:44]
  assign _GEN_175 = _T_1058 ? $signed(io_dataIn_bits_173) : $signed(buffers_0_43_1); // @[MuxLayer.scala 22:44]
  assign _GEN_176 = _T_1058 ? $signed(io_dataIn_bits_174) : $signed(buffers_0_43_2); // @[MuxLayer.scala 22:44]
  assign _GEN_177 = _T_1058 ? $signed(io_dataIn_bits_175) : $signed(buffers_0_43_3); // @[MuxLayer.scala 22:44]
  assign _GEN_178 = _T_1058 ? $signed(io_dataIn_bits_176) : $signed(buffers_0_44_0); // @[MuxLayer.scala 22:44]
  assign _GEN_179 = _T_1058 ? $signed(io_dataIn_bits_177) : $signed(buffers_0_44_1); // @[MuxLayer.scala 22:44]
  assign _GEN_180 = _T_1058 ? $signed(io_dataIn_bits_178) : $signed(buffers_0_44_2); // @[MuxLayer.scala 22:44]
  assign _GEN_181 = _T_1058 ? $signed(io_dataIn_bits_179) : $signed(buffers_0_44_3); // @[MuxLayer.scala 22:44]
  assign _GEN_182 = _T_1058 ? $signed(io_dataIn_bits_180) : $signed(buffers_0_45_0); // @[MuxLayer.scala 22:44]
  assign _GEN_183 = _T_1058 ? $signed(io_dataIn_bits_181) : $signed(buffers_0_45_1); // @[MuxLayer.scala 22:44]
  assign _GEN_184 = _T_1058 ? $signed(io_dataIn_bits_182) : $signed(buffers_0_45_2); // @[MuxLayer.scala 22:44]
  assign _GEN_185 = _T_1058 ? $signed(io_dataIn_bits_183) : $signed(buffers_0_45_3); // @[MuxLayer.scala 22:44]
  assign _GEN_186 = _T_1058 ? $signed(io_dataIn_bits_184) : $signed(buffers_0_46_0); // @[MuxLayer.scala 22:44]
  assign _GEN_187 = _T_1058 ? $signed(io_dataIn_bits_185) : $signed(buffers_0_46_1); // @[MuxLayer.scala 22:44]
  assign _GEN_188 = _T_1058 ? $signed(io_dataIn_bits_186) : $signed(buffers_0_46_2); // @[MuxLayer.scala 22:44]
  assign _GEN_189 = _T_1058 ? $signed(io_dataIn_bits_187) : $signed(buffers_0_46_3); // @[MuxLayer.scala 22:44]
  assign _GEN_190 = _T_1058 ? $signed(io_dataIn_bits_188) : $signed(buffers_0_47_0); // @[MuxLayer.scala 22:44]
  assign _GEN_191 = _T_1058 ? $signed(io_dataIn_bits_189) : $signed(buffers_0_47_1); // @[MuxLayer.scala 22:44]
  assign _GEN_192 = _T_1058 ? $signed(io_dataIn_bits_190) : $signed(buffers_0_47_2); // @[MuxLayer.scala 22:44]
  assign _GEN_193 = _T_1058 ? $signed(io_dataIn_bits_191) : $signed(buffers_0_47_3); // @[MuxLayer.scala 22:44]
  assign _GEN_194 = _T_1058 ? $signed(io_dataIn_bits_192) : $signed(buffers_0_48_0); // @[MuxLayer.scala 22:44]
  assign _GEN_195 = _T_1058 ? $signed(io_dataIn_bits_193) : $signed(buffers_0_48_1); // @[MuxLayer.scala 22:44]
  assign _GEN_196 = _T_1058 ? $signed(io_dataIn_bits_194) : $signed(buffers_0_48_2); // @[MuxLayer.scala 22:44]
  assign _GEN_197 = _T_1058 ? $signed(io_dataIn_bits_195) : $signed(buffers_0_48_3); // @[MuxLayer.scala 22:44]
  assign _GEN_198 = _T_1058 ? $signed(io_dataIn_bits_196) : $signed(buffers_0_49_0); // @[MuxLayer.scala 22:44]
  assign _GEN_199 = _T_1058 ? $signed(io_dataIn_bits_197) : $signed(buffers_0_49_1); // @[MuxLayer.scala 22:44]
  assign _GEN_200 = _T_1058 ? $signed(io_dataIn_bits_198) : $signed(buffers_0_49_2); // @[MuxLayer.scala 22:44]
  assign _GEN_201 = _T_1058 ? $signed(io_dataIn_bits_199) : $signed(buffers_0_49_3); // @[MuxLayer.scala 22:44]
  assign _GEN_202 = _T_1058 ? $signed(io_dataIn_bits_200) : $signed(buffers_0_50_0); // @[MuxLayer.scala 22:44]
  assign _GEN_203 = _T_1058 ? $signed(io_dataIn_bits_201) : $signed(buffers_0_50_1); // @[MuxLayer.scala 22:44]
  assign _GEN_204 = _T_1058 ? $signed(io_dataIn_bits_202) : $signed(buffers_0_50_2); // @[MuxLayer.scala 22:44]
  assign _GEN_205 = _T_1058 ? $signed(io_dataIn_bits_203) : $signed(buffers_0_50_3); // @[MuxLayer.scala 22:44]
  assign _GEN_206 = _T_1058 ? $signed(io_dataIn_bits_204) : $signed(buffers_0_51_0); // @[MuxLayer.scala 22:44]
  assign _GEN_207 = _T_1058 ? $signed(io_dataIn_bits_205) : $signed(buffers_0_51_1); // @[MuxLayer.scala 22:44]
  assign _GEN_208 = _T_1058 ? $signed(io_dataIn_bits_206) : $signed(buffers_0_51_2); // @[MuxLayer.scala 22:44]
  assign _GEN_209 = _T_1058 ? $signed(io_dataIn_bits_207) : $signed(buffers_0_51_3); // @[MuxLayer.scala 22:44]
  assign _GEN_210 = _T_1058 ? $signed(io_dataIn_bits_208) : $signed(buffers_0_52_0); // @[MuxLayer.scala 22:44]
  assign _GEN_211 = _T_1058 ? $signed(io_dataIn_bits_209) : $signed(buffers_0_52_1); // @[MuxLayer.scala 22:44]
  assign _GEN_212 = _T_1058 ? $signed(io_dataIn_bits_210) : $signed(buffers_0_52_2); // @[MuxLayer.scala 22:44]
  assign _GEN_213 = _T_1058 ? $signed(io_dataIn_bits_211) : $signed(buffers_0_52_3); // @[MuxLayer.scala 22:44]
  assign _GEN_214 = _T_1058 ? $signed(io_dataIn_bits_212) : $signed(buffers_0_53_0); // @[MuxLayer.scala 22:44]
  assign _GEN_215 = _T_1058 ? $signed(io_dataIn_bits_213) : $signed(buffers_0_53_1); // @[MuxLayer.scala 22:44]
  assign _GEN_216 = _T_1058 ? $signed(io_dataIn_bits_214) : $signed(buffers_0_53_2); // @[MuxLayer.scala 22:44]
  assign _GEN_217 = _T_1058 ? $signed(io_dataIn_bits_215) : $signed(buffers_0_53_3); // @[MuxLayer.scala 22:44]
  assign _GEN_218 = _T_1058 ? $signed(io_dataIn_bits_216) : $signed(buffers_0_54_0); // @[MuxLayer.scala 22:44]
  assign _GEN_219 = _T_1058 ? $signed(io_dataIn_bits_217) : $signed(buffers_0_54_1); // @[MuxLayer.scala 22:44]
  assign _GEN_220 = _T_1058 ? $signed(io_dataIn_bits_218) : $signed(buffers_0_54_2); // @[MuxLayer.scala 22:44]
  assign _GEN_221 = _T_1058 ? $signed(io_dataIn_bits_219) : $signed(buffers_0_54_3); // @[MuxLayer.scala 22:44]
  assign _GEN_222 = _T_1058 ? $signed(io_dataIn_bits_220) : $signed(buffers_0_55_0); // @[MuxLayer.scala 22:44]
  assign _GEN_223 = _T_1058 ? $signed(io_dataIn_bits_221) : $signed(buffers_0_55_1); // @[MuxLayer.scala 22:44]
  assign _GEN_224 = _T_1058 ? $signed(io_dataIn_bits_222) : $signed(buffers_0_55_2); // @[MuxLayer.scala 22:44]
  assign _GEN_225 = _T_1058 ? $signed(io_dataIn_bits_223) : $signed(buffers_0_55_3); // @[MuxLayer.scala 22:44]
  assign _GEN_226 = _T_1058 ? $signed(io_dataIn_bits_224) : $signed(buffers_0_56_0); // @[MuxLayer.scala 22:44]
  assign _GEN_227 = _T_1058 ? $signed(io_dataIn_bits_225) : $signed(buffers_0_56_1); // @[MuxLayer.scala 22:44]
  assign _GEN_228 = _T_1058 ? $signed(io_dataIn_bits_226) : $signed(buffers_0_56_2); // @[MuxLayer.scala 22:44]
  assign _GEN_229 = _T_1058 ? $signed(io_dataIn_bits_227) : $signed(buffers_0_56_3); // @[MuxLayer.scala 22:44]
  assign _GEN_230 = _T_1058 ? $signed(io_dataIn_bits_228) : $signed(buffers_0_57_0); // @[MuxLayer.scala 22:44]
  assign _GEN_231 = _T_1058 ? $signed(io_dataIn_bits_229) : $signed(buffers_0_57_1); // @[MuxLayer.scala 22:44]
  assign _GEN_232 = _T_1058 ? $signed(io_dataIn_bits_230) : $signed(buffers_0_57_2); // @[MuxLayer.scala 22:44]
  assign _GEN_233 = _T_1058 ? $signed(io_dataIn_bits_231) : $signed(buffers_0_57_3); // @[MuxLayer.scala 22:44]
  assign _GEN_234 = _T_1058 ? $signed(io_dataIn_bits_232) : $signed(buffers_0_58_0); // @[MuxLayer.scala 22:44]
  assign _GEN_235 = _T_1058 ? $signed(io_dataIn_bits_233) : $signed(buffers_0_58_1); // @[MuxLayer.scala 22:44]
  assign _GEN_236 = _T_1058 ? $signed(io_dataIn_bits_234) : $signed(buffers_0_58_2); // @[MuxLayer.scala 22:44]
  assign _GEN_237 = _T_1058 ? $signed(io_dataIn_bits_235) : $signed(buffers_0_58_3); // @[MuxLayer.scala 22:44]
  assign _GEN_238 = _T_1058 ? $signed(io_dataIn_bits_236) : $signed(buffers_0_59_0); // @[MuxLayer.scala 22:44]
  assign _GEN_239 = _T_1058 ? $signed(io_dataIn_bits_237) : $signed(buffers_0_59_1); // @[MuxLayer.scala 22:44]
  assign _GEN_240 = _T_1058 ? $signed(io_dataIn_bits_238) : $signed(buffers_0_59_2); // @[MuxLayer.scala 22:44]
  assign _GEN_241 = _T_1058 ? $signed(io_dataIn_bits_239) : $signed(buffers_0_59_3); // @[MuxLayer.scala 22:44]
  assign _GEN_242 = _T_1058 ? $signed(io_dataIn_bits_240) : $signed(buffers_0_60_0); // @[MuxLayer.scala 22:44]
  assign _GEN_243 = _T_1058 ? $signed(io_dataIn_bits_241) : $signed(buffers_0_60_1); // @[MuxLayer.scala 22:44]
  assign _GEN_244 = _T_1058 ? $signed(io_dataIn_bits_242) : $signed(buffers_0_60_2); // @[MuxLayer.scala 22:44]
  assign _GEN_245 = _T_1058 ? $signed(io_dataIn_bits_243) : $signed(buffers_0_60_3); // @[MuxLayer.scala 22:44]
  assign _GEN_246 = _T_1058 ? $signed(io_dataIn_bits_244) : $signed(buffers_0_61_0); // @[MuxLayer.scala 22:44]
  assign _GEN_247 = _T_1058 ? $signed(io_dataIn_bits_245) : $signed(buffers_0_61_1); // @[MuxLayer.scala 22:44]
  assign _GEN_248 = _T_1058 ? $signed(io_dataIn_bits_246) : $signed(buffers_0_61_2); // @[MuxLayer.scala 22:44]
  assign _GEN_249 = _T_1058 ? $signed(io_dataIn_bits_247) : $signed(buffers_0_61_3); // @[MuxLayer.scala 22:44]
  assign _GEN_250 = _T_1058 ? $signed(io_dataIn_bits_248) : $signed(buffers_0_62_0); // @[MuxLayer.scala 22:44]
  assign _GEN_251 = _T_1058 ? $signed(io_dataIn_bits_249) : $signed(buffers_0_62_1); // @[MuxLayer.scala 22:44]
  assign _GEN_252 = _T_1058 ? $signed(io_dataIn_bits_250) : $signed(buffers_0_62_2); // @[MuxLayer.scala 22:44]
  assign _GEN_253 = _T_1058 ? $signed(io_dataIn_bits_251) : $signed(buffers_0_62_3); // @[MuxLayer.scala 22:44]
  assign _GEN_254 = _T_1058 ? $signed(io_dataIn_bits_252) : $signed(buffers_0_63_0); // @[MuxLayer.scala 22:44]
  assign _GEN_255 = _T_1058 ? $signed(io_dataIn_bits_253) : $signed(buffers_0_63_1); // @[MuxLayer.scala 22:44]
  assign _GEN_256 = _T_1058 ? $signed(io_dataIn_bits_254) : $signed(buffers_0_63_2); // @[MuxLayer.scala 22:44]
  assign _GEN_257 = _T_1058 ? $signed(io_dataIn_bits_255) : $signed(buffers_0_63_3); // @[MuxLayer.scala 22:44]
  assign _T_1061 = cntr == 6'h3f; // @[MuxLayer.scala 29:15]
  assign _GEN_258 = _T_1061 ? 1'h1 : rdyReg; // @[MuxLayer.scala 29:36]
  assign _T_1063 = io_dataIn_valid & rdyReg; // @[MuxLayer.scala 32:26]
  assign _GEN_259 = _T_1063 ? 1'h0 : _GEN_258; // @[MuxLayer.scala 32:38]
  assign _T_1065 = cntr[1:0]; // @[MuxLayer.scala 45:19]
  assign _T_1068 = cntr[3:2]; // @[MuxLayer.scala 45:19]
  assign _T_1073 = cntr[5:4]; // @[MuxLayer.scala 45:19]
  assign _T_1090 = cntrs_0 == 2'h1; // @[MuxLayer.scala 55:25]
  assign _GEN_266 = _T_1090 ? $signed(buffers_0_1_0) : $signed(buffers_0_0_0); // @[MuxLayer.scala 55:35]
  assign _GEN_267 = _T_1090 ? $signed(buffers_0_1_1) : $signed(buffers_0_0_1); // @[MuxLayer.scala 55:35]
  assign _GEN_268 = _T_1090 ? $signed(buffers_0_1_2) : $signed(buffers_0_0_2); // @[MuxLayer.scala 55:35]
  assign _GEN_269 = _T_1090 ? $signed(buffers_0_1_3) : $signed(buffers_0_0_3); // @[MuxLayer.scala 55:35]
  assign _T_1092 = cntrs_0 == 2'h2; // @[MuxLayer.scala 55:25]
  assign _GEN_270 = _T_1092 ? $signed(buffers_0_2_0) : $signed(_GEN_266); // @[MuxLayer.scala 55:35]
  assign _GEN_271 = _T_1092 ? $signed(buffers_0_2_1) : $signed(_GEN_267); // @[MuxLayer.scala 55:35]
  assign _GEN_272 = _T_1092 ? $signed(buffers_0_2_2) : $signed(_GEN_268); // @[MuxLayer.scala 55:35]
  assign _GEN_273 = _T_1092 ? $signed(buffers_0_2_3) : $signed(_GEN_269); // @[MuxLayer.scala 55:35]
  assign _T_1094 = cntrs_0 == 2'h3; // @[MuxLayer.scala 55:25]
  assign _GEN_274 = _T_1094 ? $signed(buffers_0_3_0) : $signed(_GEN_270); // @[MuxLayer.scala 55:35]
  assign _GEN_275 = _T_1094 ? $signed(buffers_0_3_1) : $signed(_GEN_271); // @[MuxLayer.scala 55:35]
  assign _GEN_276 = _T_1094 ? $signed(buffers_0_3_2) : $signed(_GEN_272); // @[MuxLayer.scala 55:35]
  assign _GEN_277 = _T_1094 ? $signed(buffers_0_3_3) : $signed(_GEN_273); // @[MuxLayer.scala 55:35]
  assign _GEN_278 = _T_1090 ? $signed(buffers_0_5_0) : $signed(buffers_0_4_0); // @[MuxLayer.scala 55:35]
  assign _GEN_279 = _T_1090 ? $signed(buffers_0_5_1) : $signed(buffers_0_4_1); // @[MuxLayer.scala 55:35]
  assign _GEN_280 = _T_1090 ? $signed(buffers_0_5_2) : $signed(buffers_0_4_2); // @[MuxLayer.scala 55:35]
  assign _GEN_281 = _T_1090 ? $signed(buffers_0_5_3) : $signed(buffers_0_4_3); // @[MuxLayer.scala 55:35]
  assign _GEN_282 = _T_1092 ? $signed(buffers_0_6_0) : $signed(_GEN_278); // @[MuxLayer.scala 55:35]
  assign _GEN_283 = _T_1092 ? $signed(buffers_0_6_1) : $signed(_GEN_279); // @[MuxLayer.scala 55:35]
  assign _GEN_284 = _T_1092 ? $signed(buffers_0_6_2) : $signed(_GEN_280); // @[MuxLayer.scala 55:35]
  assign _GEN_285 = _T_1092 ? $signed(buffers_0_6_3) : $signed(_GEN_281); // @[MuxLayer.scala 55:35]
  assign _GEN_286 = _T_1094 ? $signed(buffers_0_7_0) : $signed(_GEN_282); // @[MuxLayer.scala 55:35]
  assign _GEN_287 = _T_1094 ? $signed(buffers_0_7_1) : $signed(_GEN_283); // @[MuxLayer.scala 55:35]
  assign _GEN_288 = _T_1094 ? $signed(buffers_0_7_2) : $signed(_GEN_284); // @[MuxLayer.scala 55:35]
  assign _GEN_289 = _T_1094 ? $signed(buffers_0_7_3) : $signed(_GEN_285); // @[MuxLayer.scala 55:35]
  assign _GEN_290 = _T_1090 ? $signed(buffers_0_9_0) : $signed(buffers_0_8_0); // @[MuxLayer.scala 55:35]
  assign _GEN_291 = _T_1090 ? $signed(buffers_0_9_1) : $signed(buffers_0_8_1); // @[MuxLayer.scala 55:35]
  assign _GEN_292 = _T_1090 ? $signed(buffers_0_9_2) : $signed(buffers_0_8_2); // @[MuxLayer.scala 55:35]
  assign _GEN_293 = _T_1090 ? $signed(buffers_0_9_3) : $signed(buffers_0_8_3); // @[MuxLayer.scala 55:35]
  assign _GEN_294 = _T_1092 ? $signed(buffers_0_10_0) : $signed(_GEN_290); // @[MuxLayer.scala 55:35]
  assign _GEN_295 = _T_1092 ? $signed(buffers_0_10_1) : $signed(_GEN_291); // @[MuxLayer.scala 55:35]
  assign _GEN_296 = _T_1092 ? $signed(buffers_0_10_2) : $signed(_GEN_292); // @[MuxLayer.scala 55:35]
  assign _GEN_297 = _T_1092 ? $signed(buffers_0_10_3) : $signed(_GEN_293); // @[MuxLayer.scala 55:35]
  assign _GEN_298 = _T_1094 ? $signed(buffers_0_11_0) : $signed(_GEN_294); // @[MuxLayer.scala 55:35]
  assign _GEN_299 = _T_1094 ? $signed(buffers_0_11_1) : $signed(_GEN_295); // @[MuxLayer.scala 55:35]
  assign _GEN_300 = _T_1094 ? $signed(buffers_0_11_2) : $signed(_GEN_296); // @[MuxLayer.scala 55:35]
  assign _GEN_301 = _T_1094 ? $signed(buffers_0_11_3) : $signed(_GEN_297); // @[MuxLayer.scala 55:35]
  assign _GEN_302 = _T_1090 ? $signed(buffers_0_13_0) : $signed(buffers_0_12_0); // @[MuxLayer.scala 55:35]
  assign _GEN_303 = _T_1090 ? $signed(buffers_0_13_1) : $signed(buffers_0_12_1); // @[MuxLayer.scala 55:35]
  assign _GEN_304 = _T_1090 ? $signed(buffers_0_13_2) : $signed(buffers_0_12_2); // @[MuxLayer.scala 55:35]
  assign _GEN_305 = _T_1090 ? $signed(buffers_0_13_3) : $signed(buffers_0_12_3); // @[MuxLayer.scala 55:35]
  assign _GEN_306 = _T_1092 ? $signed(buffers_0_14_0) : $signed(_GEN_302); // @[MuxLayer.scala 55:35]
  assign _GEN_307 = _T_1092 ? $signed(buffers_0_14_1) : $signed(_GEN_303); // @[MuxLayer.scala 55:35]
  assign _GEN_308 = _T_1092 ? $signed(buffers_0_14_2) : $signed(_GEN_304); // @[MuxLayer.scala 55:35]
  assign _GEN_309 = _T_1092 ? $signed(buffers_0_14_3) : $signed(_GEN_305); // @[MuxLayer.scala 55:35]
  assign _GEN_310 = _T_1094 ? $signed(buffers_0_15_0) : $signed(_GEN_306); // @[MuxLayer.scala 55:35]
  assign _GEN_311 = _T_1094 ? $signed(buffers_0_15_1) : $signed(_GEN_307); // @[MuxLayer.scala 55:35]
  assign _GEN_312 = _T_1094 ? $signed(buffers_0_15_2) : $signed(_GEN_308); // @[MuxLayer.scala 55:35]
  assign _GEN_313 = _T_1094 ? $signed(buffers_0_15_3) : $signed(_GEN_309); // @[MuxLayer.scala 55:35]
  assign _GEN_314 = _T_1090 ? $signed(buffers_0_17_0) : $signed(buffers_0_16_0); // @[MuxLayer.scala 55:35]
  assign _GEN_315 = _T_1090 ? $signed(buffers_0_17_1) : $signed(buffers_0_16_1); // @[MuxLayer.scala 55:35]
  assign _GEN_316 = _T_1090 ? $signed(buffers_0_17_2) : $signed(buffers_0_16_2); // @[MuxLayer.scala 55:35]
  assign _GEN_317 = _T_1090 ? $signed(buffers_0_17_3) : $signed(buffers_0_16_3); // @[MuxLayer.scala 55:35]
  assign _GEN_318 = _T_1092 ? $signed(buffers_0_18_0) : $signed(_GEN_314); // @[MuxLayer.scala 55:35]
  assign _GEN_319 = _T_1092 ? $signed(buffers_0_18_1) : $signed(_GEN_315); // @[MuxLayer.scala 55:35]
  assign _GEN_320 = _T_1092 ? $signed(buffers_0_18_2) : $signed(_GEN_316); // @[MuxLayer.scala 55:35]
  assign _GEN_321 = _T_1092 ? $signed(buffers_0_18_3) : $signed(_GEN_317); // @[MuxLayer.scala 55:35]
  assign _GEN_322 = _T_1094 ? $signed(buffers_0_19_0) : $signed(_GEN_318); // @[MuxLayer.scala 55:35]
  assign _GEN_323 = _T_1094 ? $signed(buffers_0_19_1) : $signed(_GEN_319); // @[MuxLayer.scala 55:35]
  assign _GEN_324 = _T_1094 ? $signed(buffers_0_19_2) : $signed(_GEN_320); // @[MuxLayer.scala 55:35]
  assign _GEN_325 = _T_1094 ? $signed(buffers_0_19_3) : $signed(_GEN_321); // @[MuxLayer.scala 55:35]
  assign _GEN_326 = _T_1090 ? $signed(buffers_0_21_0) : $signed(buffers_0_20_0); // @[MuxLayer.scala 55:35]
  assign _GEN_327 = _T_1090 ? $signed(buffers_0_21_1) : $signed(buffers_0_20_1); // @[MuxLayer.scala 55:35]
  assign _GEN_328 = _T_1090 ? $signed(buffers_0_21_2) : $signed(buffers_0_20_2); // @[MuxLayer.scala 55:35]
  assign _GEN_329 = _T_1090 ? $signed(buffers_0_21_3) : $signed(buffers_0_20_3); // @[MuxLayer.scala 55:35]
  assign _GEN_330 = _T_1092 ? $signed(buffers_0_22_0) : $signed(_GEN_326); // @[MuxLayer.scala 55:35]
  assign _GEN_331 = _T_1092 ? $signed(buffers_0_22_1) : $signed(_GEN_327); // @[MuxLayer.scala 55:35]
  assign _GEN_332 = _T_1092 ? $signed(buffers_0_22_2) : $signed(_GEN_328); // @[MuxLayer.scala 55:35]
  assign _GEN_333 = _T_1092 ? $signed(buffers_0_22_3) : $signed(_GEN_329); // @[MuxLayer.scala 55:35]
  assign _GEN_334 = _T_1094 ? $signed(buffers_0_23_0) : $signed(_GEN_330); // @[MuxLayer.scala 55:35]
  assign _GEN_335 = _T_1094 ? $signed(buffers_0_23_1) : $signed(_GEN_331); // @[MuxLayer.scala 55:35]
  assign _GEN_336 = _T_1094 ? $signed(buffers_0_23_2) : $signed(_GEN_332); // @[MuxLayer.scala 55:35]
  assign _GEN_337 = _T_1094 ? $signed(buffers_0_23_3) : $signed(_GEN_333); // @[MuxLayer.scala 55:35]
  assign _GEN_338 = _T_1090 ? $signed(buffers_0_25_0) : $signed(buffers_0_24_0); // @[MuxLayer.scala 55:35]
  assign _GEN_339 = _T_1090 ? $signed(buffers_0_25_1) : $signed(buffers_0_24_1); // @[MuxLayer.scala 55:35]
  assign _GEN_340 = _T_1090 ? $signed(buffers_0_25_2) : $signed(buffers_0_24_2); // @[MuxLayer.scala 55:35]
  assign _GEN_341 = _T_1090 ? $signed(buffers_0_25_3) : $signed(buffers_0_24_3); // @[MuxLayer.scala 55:35]
  assign _GEN_342 = _T_1092 ? $signed(buffers_0_26_0) : $signed(_GEN_338); // @[MuxLayer.scala 55:35]
  assign _GEN_343 = _T_1092 ? $signed(buffers_0_26_1) : $signed(_GEN_339); // @[MuxLayer.scala 55:35]
  assign _GEN_344 = _T_1092 ? $signed(buffers_0_26_2) : $signed(_GEN_340); // @[MuxLayer.scala 55:35]
  assign _GEN_345 = _T_1092 ? $signed(buffers_0_26_3) : $signed(_GEN_341); // @[MuxLayer.scala 55:35]
  assign _GEN_346 = _T_1094 ? $signed(buffers_0_27_0) : $signed(_GEN_342); // @[MuxLayer.scala 55:35]
  assign _GEN_347 = _T_1094 ? $signed(buffers_0_27_1) : $signed(_GEN_343); // @[MuxLayer.scala 55:35]
  assign _GEN_348 = _T_1094 ? $signed(buffers_0_27_2) : $signed(_GEN_344); // @[MuxLayer.scala 55:35]
  assign _GEN_349 = _T_1094 ? $signed(buffers_0_27_3) : $signed(_GEN_345); // @[MuxLayer.scala 55:35]
  assign _GEN_350 = _T_1090 ? $signed(buffers_0_29_0) : $signed(buffers_0_28_0); // @[MuxLayer.scala 55:35]
  assign _GEN_351 = _T_1090 ? $signed(buffers_0_29_1) : $signed(buffers_0_28_1); // @[MuxLayer.scala 55:35]
  assign _GEN_352 = _T_1090 ? $signed(buffers_0_29_2) : $signed(buffers_0_28_2); // @[MuxLayer.scala 55:35]
  assign _GEN_353 = _T_1090 ? $signed(buffers_0_29_3) : $signed(buffers_0_28_3); // @[MuxLayer.scala 55:35]
  assign _GEN_354 = _T_1092 ? $signed(buffers_0_30_0) : $signed(_GEN_350); // @[MuxLayer.scala 55:35]
  assign _GEN_355 = _T_1092 ? $signed(buffers_0_30_1) : $signed(_GEN_351); // @[MuxLayer.scala 55:35]
  assign _GEN_356 = _T_1092 ? $signed(buffers_0_30_2) : $signed(_GEN_352); // @[MuxLayer.scala 55:35]
  assign _GEN_357 = _T_1092 ? $signed(buffers_0_30_3) : $signed(_GEN_353); // @[MuxLayer.scala 55:35]
  assign _GEN_358 = _T_1094 ? $signed(buffers_0_31_0) : $signed(_GEN_354); // @[MuxLayer.scala 55:35]
  assign _GEN_359 = _T_1094 ? $signed(buffers_0_31_1) : $signed(_GEN_355); // @[MuxLayer.scala 55:35]
  assign _GEN_360 = _T_1094 ? $signed(buffers_0_31_2) : $signed(_GEN_356); // @[MuxLayer.scala 55:35]
  assign _GEN_361 = _T_1094 ? $signed(buffers_0_31_3) : $signed(_GEN_357); // @[MuxLayer.scala 55:35]
  assign _GEN_362 = _T_1090 ? $signed(buffers_0_33_0) : $signed(buffers_0_32_0); // @[MuxLayer.scala 55:35]
  assign _GEN_363 = _T_1090 ? $signed(buffers_0_33_1) : $signed(buffers_0_32_1); // @[MuxLayer.scala 55:35]
  assign _GEN_364 = _T_1090 ? $signed(buffers_0_33_2) : $signed(buffers_0_32_2); // @[MuxLayer.scala 55:35]
  assign _GEN_365 = _T_1090 ? $signed(buffers_0_33_3) : $signed(buffers_0_32_3); // @[MuxLayer.scala 55:35]
  assign _GEN_366 = _T_1092 ? $signed(buffers_0_34_0) : $signed(_GEN_362); // @[MuxLayer.scala 55:35]
  assign _GEN_367 = _T_1092 ? $signed(buffers_0_34_1) : $signed(_GEN_363); // @[MuxLayer.scala 55:35]
  assign _GEN_368 = _T_1092 ? $signed(buffers_0_34_2) : $signed(_GEN_364); // @[MuxLayer.scala 55:35]
  assign _GEN_369 = _T_1092 ? $signed(buffers_0_34_3) : $signed(_GEN_365); // @[MuxLayer.scala 55:35]
  assign _GEN_370 = _T_1094 ? $signed(buffers_0_35_0) : $signed(_GEN_366); // @[MuxLayer.scala 55:35]
  assign _GEN_371 = _T_1094 ? $signed(buffers_0_35_1) : $signed(_GEN_367); // @[MuxLayer.scala 55:35]
  assign _GEN_372 = _T_1094 ? $signed(buffers_0_35_2) : $signed(_GEN_368); // @[MuxLayer.scala 55:35]
  assign _GEN_373 = _T_1094 ? $signed(buffers_0_35_3) : $signed(_GEN_369); // @[MuxLayer.scala 55:35]
  assign _GEN_374 = _T_1090 ? $signed(buffers_0_37_0) : $signed(buffers_0_36_0); // @[MuxLayer.scala 55:35]
  assign _GEN_375 = _T_1090 ? $signed(buffers_0_37_1) : $signed(buffers_0_36_1); // @[MuxLayer.scala 55:35]
  assign _GEN_376 = _T_1090 ? $signed(buffers_0_37_2) : $signed(buffers_0_36_2); // @[MuxLayer.scala 55:35]
  assign _GEN_377 = _T_1090 ? $signed(buffers_0_37_3) : $signed(buffers_0_36_3); // @[MuxLayer.scala 55:35]
  assign _GEN_378 = _T_1092 ? $signed(buffers_0_38_0) : $signed(_GEN_374); // @[MuxLayer.scala 55:35]
  assign _GEN_379 = _T_1092 ? $signed(buffers_0_38_1) : $signed(_GEN_375); // @[MuxLayer.scala 55:35]
  assign _GEN_380 = _T_1092 ? $signed(buffers_0_38_2) : $signed(_GEN_376); // @[MuxLayer.scala 55:35]
  assign _GEN_381 = _T_1092 ? $signed(buffers_0_38_3) : $signed(_GEN_377); // @[MuxLayer.scala 55:35]
  assign _GEN_382 = _T_1094 ? $signed(buffers_0_39_0) : $signed(_GEN_378); // @[MuxLayer.scala 55:35]
  assign _GEN_383 = _T_1094 ? $signed(buffers_0_39_1) : $signed(_GEN_379); // @[MuxLayer.scala 55:35]
  assign _GEN_384 = _T_1094 ? $signed(buffers_0_39_2) : $signed(_GEN_380); // @[MuxLayer.scala 55:35]
  assign _GEN_385 = _T_1094 ? $signed(buffers_0_39_3) : $signed(_GEN_381); // @[MuxLayer.scala 55:35]
  assign _GEN_386 = _T_1090 ? $signed(buffers_0_41_0) : $signed(buffers_0_40_0); // @[MuxLayer.scala 55:35]
  assign _GEN_387 = _T_1090 ? $signed(buffers_0_41_1) : $signed(buffers_0_40_1); // @[MuxLayer.scala 55:35]
  assign _GEN_388 = _T_1090 ? $signed(buffers_0_41_2) : $signed(buffers_0_40_2); // @[MuxLayer.scala 55:35]
  assign _GEN_389 = _T_1090 ? $signed(buffers_0_41_3) : $signed(buffers_0_40_3); // @[MuxLayer.scala 55:35]
  assign _GEN_390 = _T_1092 ? $signed(buffers_0_42_0) : $signed(_GEN_386); // @[MuxLayer.scala 55:35]
  assign _GEN_391 = _T_1092 ? $signed(buffers_0_42_1) : $signed(_GEN_387); // @[MuxLayer.scala 55:35]
  assign _GEN_392 = _T_1092 ? $signed(buffers_0_42_2) : $signed(_GEN_388); // @[MuxLayer.scala 55:35]
  assign _GEN_393 = _T_1092 ? $signed(buffers_0_42_3) : $signed(_GEN_389); // @[MuxLayer.scala 55:35]
  assign _GEN_394 = _T_1094 ? $signed(buffers_0_43_0) : $signed(_GEN_390); // @[MuxLayer.scala 55:35]
  assign _GEN_395 = _T_1094 ? $signed(buffers_0_43_1) : $signed(_GEN_391); // @[MuxLayer.scala 55:35]
  assign _GEN_396 = _T_1094 ? $signed(buffers_0_43_2) : $signed(_GEN_392); // @[MuxLayer.scala 55:35]
  assign _GEN_397 = _T_1094 ? $signed(buffers_0_43_3) : $signed(_GEN_393); // @[MuxLayer.scala 55:35]
  assign _GEN_398 = _T_1090 ? $signed(buffers_0_45_0) : $signed(buffers_0_44_0); // @[MuxLayer.scala 55:35]
  assign _GEN_399 = _T_1090 ? $signed(buffers_0_45_1) : $signed(buffers_0_44_1); // @[MuxLayer.scala 55:35]
  assign _GEN_400 = _T_1090 ? $signed(buffers_0_45_2) : $signed(buffers_0_44_2); // @[MuxLayer.scala 55:35]
  assign _GEN_401 = _T_1090 ? $signed(buffers_0_45_3) : $signed(buffers_0_44_3); // @[MuxLayer.scala 55:35]
  assign _GEN_402 = _T_1092 ? $signed(buffers_0_46_0) : $signed(_GEN_398); // @[MuxLayer.scala 55:35]
  assign _GEN_403 = _T_1092 ? $signed(buffers_0_46_1) : $signed(_GEN_399); // @[MuxLayer.scala 55:35]
  assign _GEN_404 = _T_1092 ? $signed(buffers_0_46_2) : $signed(_GEN_400); // @[MuxLayer.scala 55:35]
  assign _GEN_405 = _T_1092 ? $signed(buffers_0_46_3) : $signed(_GEN_401); // @[MuxLayer.scala 55:35]
  assign _GEN_406 = _T_1094 ? $signed(buffers_0_47_0) : $signed(_GEN_402); // @[MuxLayer.scala 55:35]
  assign _GEN_407 = _T_1094 ? $signed(buffers_0_47_1) : $signed(_GEN_403); // @[MuxLayer.scala 55:35]
  assign _GEN_408 = _T_1094 ? $signed(buffers_0_47_2) : $signed(_GEN_404); // @[MuxLayer.scala 55:35]
  assign _GEN_409 = _T_1094 ? $signed(buffers_0_47_3) : $signed(_GEN_405); // @[MuxLayer.scala 55:35]
  assign _GEN_410 = _T_1090 ? $signed(buffers_0_49_0) : $signed(buffers_0_48_0); // @[MuxLayer.scala 55:35]
  assign _GEN_411 = _T_1090 ? $signed(buffers_0_49_1) : $signed(buffers_0_48_1); // @[MuxLayer.scala 55:35]
  assign _GEN_412 = _T_1090 ? $signed(buffers_0_49_2) : $signed(buffers_0_48_2); // @[MuxLayer.scala 55:35]
  assign _GEN_413 = _T_1090 ? $signed(buffers_0_49_3) : $signed(buffers_0_48_3); // @[MuxLayer.scala 55:35]
  assign _GEN_414 = _T_1092 ? $signed(buffers_0_50_0) : $signed(_GEN_410); // @[MuxLayer.scala 55:35]
  assign _GEN_415 = _T_1092 ? $signed(buffers_0_50_1) : $signed(_GEN_411); // @[MuxLayer.scala 55:35]
  assign _GEN_416 = _T_1092 ? $signed(buffers_0_50_2) : $signed(_GEN_412); // @[MuxLayer.scala 55:35]
  assign _GEN_417 = _T_1092 ? $signed(buffers_0_50_3) : $signed(_GEN_413); // @[MuxLayer.scala 55:35]
  assign _GEN_418 = _T_1094 ? $signed(buffers_0_51_0) : $signed(_GEN_414); // @[MuxLayer.scala 55:35]
  assign _GEN_419 = _T_1094 ? $signed(buffers_0_51_1) : $signed(_GEN_415); // @[MuxLayer.scala 55:35]
  assign _GEN_420 = _T_1094 ? $signed(buffers_0_51_2) : $signed(_GEN_416); // @[MuxLayer.scala 55:35]
  assign _GEN_421 = _T_1094 ? $signed(buffers_0_51_3) : $signed(_GEN_417); // @[MuxLayer.scala 55:35]
  assign _GEN_422 = _T_1090 ? $signed(buffers_0_53_0) : $signed(buffers_0_52_0); // @[MuxLayer.scala 55:35]
  assign _GEN_423 = _T_1090 ? $signed(buffers_0_53_1) : $signed(buffers_0_52_1); // @[MuxLayer.scala 55:35]
  assign _GEN_424 = _T_1090 ? $signed(buffers_0_53_2) : $signed(buffers_0_52_2); // @[MuxLayer.scala 55:35]
  assign _GEN_425 = _T_1090 ? $signed(buffers_0_53_3) : $signed(buffers_0_52_3); // @[MuxLayer.scala 55:35]
  assign _GEN_426 = _T_1092 ? $signed(buffers_0_54_0) : $signed(_GEN_422); // @[MuxLayer.scala 55:35]
  assign _GEN_427 = _T_1092 ? $signed(buffers_0_54_1) : $signed(_GEN_423); // @[MuxLayer.scala 55:35]
  assign _GEN_428 = _T_1092 ? $signed(buffers_0_54_2) : $signed(_GEN_424); // @[MuxLayer.scala 55:35]
  assign _GEN_429 = _T_1092 ? $signed(buffers_0_54_3) : $signed(_GEN_425); // @[MuxLayer.scala 55:35]
  assign _GEN_430 = _T_1094 ? $signed(buffers_0_55_0) : $signed(_GEN_426); // @[MuxLayer.scala 55:35]
  assign _GEN_431 = _T_1094 ? $signed(buffers_0_55_1) : $signed(_GEN_427); // @[MuxLayer.scala 55:35]
  assign _GEN_432 = _T_1094 ? $signed(buffers_0_55_2) : $signed(_GEN_428); // @[MuxLayer.scala 55:35]
  assign _GEN_433 = _T_1094 ? $signed(buffers_0_55_3) : $signed(_GEN_429); // @[MuxLayer.scala 55:35]
  assign _GEN_434 = _T_1090 ? $signed(buffers_0_57_0) : $signed(buffers_0_56_0); // @[MuxLayer.scala 55:35]
  assign _GEN_435 = _T_1090 ? $signed(buffers_0_57_1) : $signed(buffers_0_56_1); // @[MuxLayer.scala 55:35]
  assign _GEN_436 = _T_1090 ? $signed(buffers_0_57_2) : $signed(buffers_0_56_2); // @[MuxLayer.scala 55:35]
  assign _GEN_437 = _T_1090 ? $signed(buffers_0_57_3) : $signed(buffers_0_56_3); // @[MuxLayer.scala 55:35]
  assign _GEN_438 = _T_1092 ? $signed(buffers_0_58_0) : $signed(_GEN_434); // @[MuxLayer.scala 55:35]
  assign _GEN_439 = _T_1092 ? $signed(buffers_0_58_1) : $signed(_GEN_435); // @[MuxLayer.scala 55:35]
  assign _GEN_440 = _T_1092 ? $signed(buffers_0_58_2) : $signed(_GEN_436); // @[MuxLayer.scala 55:35]
  assign _GEN_441 = _T_1092 ? $signed(buffers_0_58_3) : $signed(_GEN_437); // @[MuxLayer.scala 55:35]
  assign _GEN_442 = _T_1094 ? $signed(buffers_0_59_0) : $signed(_GEN_438); // @[MuxLayer.scala 55:35]
  assign _GEN_443 = _T_1094 ? $signed(buffers_0_59_1) : $signed(_GEN_439); // @[MuxLayer.scala 55:35]
  assign _GEN_444 = _T_1094 ? $signed(buffers_0_59_2) : $signed(_GEN_440); // @[MuxLayer.scala 55:35]
  assign _GEN_445 = _T_1094 ? $signed(buffers_0_59_3) : $signed(_GEN_441); // @[MuxLayer.scala 55:35]
  assign _GEN_446 = _T_1090 ? $signed(buffers_0_61_0) : $signed(buffers_0_60_0); // @[MuxLayer.scala 55:35]
  assign _GEN_447 = _T_1090 ? $signed(buffers_0_61_1) : $signed(buffers_0_60_1); // @[MuxLayer.scala 55:35]
  assign _GEN_448 = _T_1090 ? $signed(buffers_0_61_2) : $signed(buffers_0_60_2); // @[MuxLayer.scala 55:35]
  assign _GEN_449 = _T_1090 ? $signed(buffers_0_61_3) : $signed(buffers_0_60_3); // @[MuxLayer.scala 55:35]
  assign _GEN_450 = _T_1092 ? $signed(buffers_0_62_0) : $signed(_GEN_446); // @[MuxLayer.scala 55:35]
  assign _GEN_451 = _T_1092 ? $signed(buffers_0_62_1) : $signed(_GEN_447); // @[MuxLayer.scala 55:35]
  assign _GEN_452 = _T_1092 ? $signed(buffers_0_62_2) : $signed(_GEN_448); // @[MuxLayer.scala 55:35]
  assign _GEN_453 = _T_1092 ? $signed(buffers_0_62_3) : $signed(_GEN_449); // @[MuxLayer.scala 55:35]
  assign _GEN_454 = _T_1094 ? $signed(buffers_0_63_0) : $signed(_GEN_450); // @[MuxLayer.scala 55:35]
  assign _GEN_455 = _T_1094 ? $signed(buffers_0_63_1) : $signed(_GEN_451); // @[MuxLayer.scala 55:35]
  assign _GEN_456 = _T_1094 ? $signed(buffers_0_63_2) : $signed(_GEN_452); // @[MuxLayer.scala 55:35]
  assign _GEN_457 = _T_1094 ? $signed(buffers_0_63_3) : $signed(_GEN_453); // @[MuxLayer.scala 55:35]
  assign _T_1778 = cntrs_1 == 2'h1; // @[MuxLayer.scala 55:25]
  assign _GEN_458 = _T_1778 ? $signed(buffers_1_1_0) : $signed(buffers_1_0_0); // @[MuxLayer.scala 55:35]
  assign _GEN_459 = _T_1778 ? $signed(buffers_1_1_1) : $signed(buffers_1_0_1); // @[MuxLayer.scala 55:35]
  assign _GEN_460 = _T_1778 ? $signed(buffers_1_1_2) : $signed(buffers_1_0_2); // @[MuxLayer.scala 55:35]
  assign _GEN_461 = _T_1778 ? $signed(buffers_1_1_3) : $signed(buffers_1_0_3); // @[MuxLayer.scala 55:35]
  assign _T_1780 = cntrs_1 == 2'h2; // @[MuxLayer.scala 55:25]
  assign _GEN_462 = _T_1780 ? $signed(buffers_1_2_0) : $signed(_GEN_458); // @[MuxLayer.scala 55:35]
  assign _GEN_463 = _T_1780 ? $signed(buffers_1_2_1) : $signed(_GEN_459); // @[MuxLayer.scala 55:35]
  assign _GEN_464 = _T_1780 ? $signed(buffers_1_2_2) : $signed(_GEN_460); // @[MuxLayer.scala 55:35]
  assign _GEN_465 = _T_1780 ? $signed(buffers_1_2_3) : $signed(_GEN_461); // @[MuxLayer.scala 55:35]
  assign _T_1782 = cntrs_1 == 2'h3; // @[MuxLayer.scala 55:25]
  assign _GEN_466 = _T_1782 ? $signed(buffers_1_3_0) : $signed(_GEN_462); // @[MuxLayer.scala 55:35]
  assign _GEN_467 = _T_1782 ? $signed(buffers_1_3_1) : $signed(_GEN_463); // @[MuxLayer.scala 55:35]
  assign _GEN_468 = _T_1782 ? $signed(buffers_1_3_2) : $signed(_GEN_464); // @[MuxLayer.scala 55:35]
  assign _GEN_469 = _T_1782 ? $signed(buffers_1_3_3) : $signed(_GEN_465); // @[MuxLayer.scala 55:35]
  assign _GEN_470 = _T_1778 ? $signed(buffers_1_5_0) : $signed(buffers_1_4_0); // @[MuxLayer.scala 55:35]
  assign _GEN_471 = _T_1778 ? $signed(buffers_1_5_1) : $signed(buffers_1_4_1); // @[MuxLayer.scala 55:35]
  assign _GEN_472 = _T_1778 ? $signed(buffers_1_5_2) : $signed(buffers_1_4_2); // @[MuxLayer.scala 55:35]
  assign _GEN_473 = _T_1778 ? $signed(buffers_1_5_3) : $signed(buffers_1_4_3); // @[MuxLayer.scala 55:35]
  assign _GEN_474 = _T_1780 ? $signed(buffers_1_6_0) : $signed(_GEN_470); // @[MuxLayer.scala 55:35]
  assign _GEN_475 = _T_1780 ? $signed(buffers_1_6_1) : $signed(_GEN_471); // @[MuxLayer.scala 55:35]
  assign _GEN_476 = _T_1780 ? $signed(buffers_1_6_2) : $signed(_GEN_472); // @[MuxLayer.scala 55:35]
  assign _GEN_477 = _T_1780 ? $signed(buffers_1_6_3) : $signed(_GEN_473); // @[MuxLayer.scala 55:35]
  assign _GEN_478 = _T_1782 ? $signed(buffers_1_7_0) : $signed(_GEN_474); // @[MuxLayer.scala 55:35]
  assign _GEN_479 = _T_1782 ? $signed(buffers_1_7_1) : $signed(_GEN_475); // @[MuxLayer.scala 55:35]
  assign _GEN_480 = _T_1782 ? $signed(buffers_1_7_2) : $signed(_GEN_476); // @[MuxLayer.scala 55:35]
  assign _GEN_481 = _T_1782 ? $signed(buffers_1_7_3) : $signed(_GEN_477); // @[MuxLayer.scala 55:35]
  assign _GEN_482 = _T_1778 ? $signed(buffers_1_9_0) : $signed(buffers_1_8_0); // @[MuxLayer.scala 55:35]
  assign _GEN_483 = _T_1778 ? $signed(buffers_1_9_1) : $signed(buffers_1_8_1); // @[MuxLayer.scala 55:35]
  assign _GEN_484 = _T_1778 ? $signed(buffers_1_9_2) : $signed(buffers_1_8_2); // @[MuxLayer.scala 55:35]
  assign _GEN_485 = _T_1778 ? $signed(buffers_1_9_3) : $signed(buffers_1_8_3); // @[MuxLayer.scala 55:35]
  assign _GEN_486 = _T_1780 ? $signed(buffers_1_10_0) : $signed(_GEN_482); // @[MuxLayer.scala 55:35]
  assign _GEN_487 = _T_1780 ? $signed(buffers_1_10_1) : $signed(_GEN_483); // @[MuxLayer.scala 55:35]
  assign _GEN_488 = _T_1780 ? $signed(buffers_1_10_2) : $signed(_GEN_484); // @[MuxLayer.scala 55:35]
  assign _GEN_489 = _T_1780 ? $signed(buffers_1_10_3) : $signed(_GEN_485); // @[MuxLayer.scala 55:35]
  assign _GEN_490 = _T_1782 ? $signed(buffers_1_11_0) : $signed(_GEN_486); // @[MuxLayer.scala 55:35]
  assign _GEN_491 = _T_1782 ? $signed(buffers_1_11_1) : $signed(_GEN_487); // @[MuxLayer.scala 55:35]
  assign _GEN_492 = _T_1782 ? $signed(buffers_1_11_2) : $signed(_GEN_488); // @[MuxLayer.scala 55:35]
  assign _GEN_493 = _T_1782 ? $signed(buffers_1_11_3) : $signed(_GEN_489); // @[MuxLayer.scala 55:35]
  assign _GEN_494 = _T_1778 ? $signed(buffers_1_13_0) : $signed(buffers_1_12_0); // @[MuxLayer.scala 55:35]
  assign _GEN_495 = _T_1778 ? $signed(buffers_1_13_1) : $signed(buffers_1_12_1); // @[MuxLayer.scala 55:35]
  assign _GEN_496 = _T_1778 ? $signed(buffers_1_13_2) : $signed(buffers_1_12_2); // @[MuxLayer.scala 55:35]
  assign _GEN_497 = _T_1778 ? $signed(buffers_1_13_3) : $signed(buffers_1_12_3); // @[MuxLayer.scala 55:35]
  assign _GEN_498 = _T_1780 ? $signed(buffers_1_14_0) : $signed(_GEN_494); // @[MuxLayer.scala 55:35]
  assign _GEN_499 = _T_1780 ? $signed(buffers_1_14_1) : $signed(_GEN_495); // @[MuxLayer.scala 55:35]
  assign _GEN_500 = _T_1780 ? $signed(buffers_1_14_2) : $signed(_GEN_496); // @[MuxLayer.scala 55:35]
  assign _GEN_501 = _T_1780 ? $signed(buffers_1_14_3) : $signed(_GEN_497); // @[MuxLayer.scala 55:35]
  assign _GEN_502 = _T_1782 ? $signed(buffers_1_15_0) : $signed(_GEN_498); // @[MuxLayer.scala 55:35]
  assign _GEN_503 = _T_1782 ? $signed(buffers_1_15_1) : $signed(_GEN_499); // @[MuxLayer.scala 55:35]
  assign _GEN_504 = _T_1782 ? $signed(buffers_1_15_2) : $signed(_GEN_500); // @[MuxLayer.scala 55:35]
  assign _GEN_505 = _T_1782 ? $signed(buffers_1_15_3) : $signed(_GEN_501); // @[MuxLayer.scala 55:35]
  assign _T_1950 = cntrs_2 == 2'h1; // @[MuxLayer.scala 55:25]
  assign _GEN_506 = _T_1950 ? $signed(buffers_2_1_0) : $signed(buffers_2_0_0); // @[MuxLayer.scala 55:35]
  assign _GEN_507 = _T_1950 ? $signed(buffers_2_1_1) : $signed(buffers_2_0_1); // @[MuxLayer.scala 55:35]
  assign _GEN_508 = _T_1950 ? $signed(buffers_2_1_2) : $signed(buffers_2_0_2); // @[MuxLayer.scala 55:35]
  assign _GEN_509 = _T_1950 ? $signed(buffers_2_1_3) : $signed(buffers_2_0_3); // @[MuxLayer.scala 55:35]
  assign _T_1952 = cntrs_2 == 2'h2; // @[MuxLayer.scala 55:25]
  assign _GEN_510 = _T_1952 ? $signed(buffers_2_2_0) : $signed(_GEN_506); // @[MuxLayer.scala 55:35]
  assign _GEN_511 = _T_1952 ? $signed(buffers_2_2_1) : $signed(_GEN_507); // @[MuxLayer.scala 55:35]
  assign _GEN_512 = _T_1952 ? $signed(buffers_2_2_2) : $signed(_GEN_508); // @[MuxLayer.scala 55:35]
  assign _GEN_513 = _T_1952 ? $signed(buffers_2_2_3) : $signed(_GEN_509); // @[MuxLayer.scala 55:35]
  assign _T_1954 = cntrs_2 == 2'h3; // @[MuxLayer.scala 55:25]
  assign _GEN_514 = _T_1954 ? $signed(buffers_2_3_0) : $signed(_GEN_510); // @[MuxLayer.scala 55:35]
  assign _GEN_515 = _T_1954 ? $signed(buffers_2_3_1) : $signed(_GEN_511); // @[MuxLayer.scala 55:35]
  assign _GEN_516 = _T_1954 ? $signed(buffers_2_3_2) : $signed(_GEN_512); // @[MuxLayer.scala 55:35]
  assign _GEN_517 = _T_1954 ? $signed(buffers_2_3_3) : $signed(_GEN_513); // @[MuxLayer.scala 55:35]
  assign _T_1994 = vld | lastVld; // @[MuxLayer.scala 68:27]
  assign io_dataIn_ready = rdyReg;
  assign io_dataOut_valid = _T_1994;
  assign io_dataOut_bits_0 = buffers_3_0_0;
  assign io_dataOut_bits_1 = buffers_3_0_1;
  assign io_dataOut_bits_2 = buffers_3_0_2;
  assign io_dataOut_bits_3 = buffers_3_0_3;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  rdyReg = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  cntr = _RAND_1[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  buffers_0_0_0 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  buffers_0_0_1 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  buffers_0_0_2 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  buffers_0_0_3 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  buffers_0_1_0 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  buffers_0_1_1 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  buffers_0_1_2 = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  buffers_0_1_3 = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  buffers_0_2_0 = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  buffers_0_2_1 = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  buffers_0_2_2 = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  buffers_0_2_3 = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  buffers_0_3_0 = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  buffers_0_3_1 = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  buffers_0_3_2 = _RAND_16[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  buffers_0_3_3 = _RAND_17[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  buffers_0_4_0 = _RAND_18[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  buffers_0_4_1 = _RAND_19[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  buffers_0_4_2 = _RAND_20[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  buffers_0_4_3 = _RAND_21[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  buffers_0_5_0 = _RAND_22[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  buffers_0_5_1 = _RAND_23[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  buffers_0_5_2 = _RAND_24[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  buffers_0_5_3 = _RAND_25[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  buffers_0_6_0 = _RAND_26[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  buffers_0_6_1 = _RAND_27[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  buffers_0_6_2 = _RAND_28[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  buffers_0_6_3 = _RAND_29[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  buffers_0_7_0 = _RAND_30[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  buffers_0_7_1 = _RAND_31[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  buffers_0_7_2 = _RAND_32[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{$random}};
  buffers_0_7_3 = _RAND_33[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{$random}};
  buffers_0_8_0 = _RAND_34[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{$random}};
  buffers_0_8_1 = _RAND_35[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{$random}};
  buffers_0_8_2 = _RAND_36[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{$random}};
  buffers_0_8_3 = _RAND_37[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{$random}};
  buffers_0_9_0 = _RAND_38[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{$random}};
  buffers_0_9_1 = _RAND_39[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{$random}};
  buffers_0_9_2 = _RAND_40[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{$random}};
  buffers_0_9_3 = _RAND_41[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{$random}};
  buffers_0_10_0 = _RAND_42[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{$random}};
  buffers_0_10_1 = _RAND_43[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{$random}};
  buffers_0_10_2 = _RAND_44[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{$random}};
  buffers_0_10_3 = _RAND_45[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{$random}};
  buffers_0_11_0 = _RAND_46[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{$random}};
  buffers_0_11_1 = _RAND_47[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{$random}};
  buffers_0_11_2 = _RAND_48[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{$random}};
  buffers_0_11_3 = _RAND_49[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{$random}};
  buffers_0_12_0 = _RAND_50[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{$random}};
  buffers_0_12_1 = _RAND_51[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{$random}};
  buffers_0_12_2 = _RAND_52[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{$random}};
  buffers_0_12_3 = _RAND_53[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{$random}};
  buffers_0_13_0 = _RAND_54[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{$random}};
  buffers_0_13_1 = _RAND_55[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{$random}};
  buffers_0_13_2 = _RAND_56[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{$random}};
  buffers_0_13_3 = _RAND_57[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{$random}};
  buffers_0_14_0 = _RAND_58[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{$random}};
  buffers_0_14_1 = _RAND_59[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{$random}};
  buffers_0_14_2 = _RAND_60[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{$random}};
  buffers_0_14_3 = _RAND_61[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{$random}};
  buffers_0_15_0 = _RAND_62[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{$random}};
  buffers_0_15_1 = _RAND_63[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{$random}};
  buffers_0_15_2 = _RAND_64[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{$random}};
  buffers_0_15_3 = _RAND_65[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{$random}};
  buffers_0_16_0 = _RAND_66[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{$random}};
  buffers_0_16_1 = _RAND_67[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{$random}};
  buffers_0_16_2 = _RAND_68[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{$random}};
  buffers_0_16_3 = _RAND_69[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{$random}};
  buffers_0_17_0 = _RAND_70[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{$random}};
  buffers_0_17_1 = _RAND_71[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{$random}};
  buffers_0_17_2 = _RAND_72[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{$random}};
  buffers_0_17_3 = _RAND_73[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{$random}};
  buffers_0_18_0 = _RAND_74[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{$random}};
  buffers_0_18_1 = _RAND_75[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{$random}};
  buffers_0_18_2 = _RAND_76[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{$random}};
  buffers_0_18_3 = _RAND_77[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{$random}};
  buffers_0_19_0 = _RAND_78[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{$random}};
  buffers_0_19_1 = _RAND_79[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{$random}};
  buffers_0_19_2 = _RAND_80[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{$random}};
  buffers_0_19_3 = _RAND_81[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{$random}};
  buffers_0_20_0 = _RAND_82[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{$random}};
  buffers_0_20_1 = _RAND_83[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{$random}};
  buffers_0_20_2 = _RAND_84[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{$random}};
  buffers_0_20_3 = _RAND_85[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{$random}};
  buffers_0_21_0 = _RAND_86[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{$random}};
  buffers_0_21_1 = _RAND_87[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{$random}};
  buffers_0_21_2 = _RAND_88[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{$random}};
  buffers_0_21_3 = _RAND_89[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{$random}};
  buffers_0_22_0 = _RAND_90[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{$random}};
  buffers_0_22_1 = _RAND_91[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{$random}};
  buffers_0_22_2 = _RAND_92[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{$random}};
  buffers_0_22_3 = _RAND_93[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{$random}};
  buffers_0_23_0 = _RAND_94[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{$random}};
  buffers_0_23_1 = _RAND_95[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{$random}};
  buffers_0_23_2 = _RAND_96[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{$random}};
  buffers_0_23_3 = _RAND_97[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{$random}};
  buffers_0_24_0 = _RAND_98[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{$random}};
  buffers_0_24_1 = _RAND_99[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{$random}};
  buffers_0_24_2 = _RAND_100[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{$random}};
  buffers_0_24_3 = _RAND_101[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{$random}};
  buffers_0_25_0 = _RAND_102[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{$random}};
  buffers_0_25_1 = _RAND_103[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{$random}};
  buffers_0_25_2 = _RAND_104[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{$random}};
  buffers_0_25_3 = _RAND_105[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{$random}};
  buffers_0_26_0 = _RAND_106[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{$random}};
  buffers_0_26_1 = _RAND_107[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{$random}};
  buffers_0_26_2 = _RAND_108[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{$random}};
  buffers_0_26_3 = _RAND_109[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{$random}};
  buffers_0_27_0 = _RAND_110[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{$random}};
  buffers_0_27_1 = _RAND_111[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{$random}};
  buffers_0_27_2 = _RAND_112[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{$random}};
  buffers_0_27_3 = _RAND_113[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{$random}};
  buffers_0_28_0 = _RAND_114[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{$random}};
  buffers_0_28_1 = _RAND_115[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{$random}};
  buffers_0_28_2 = _RAND_116[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{$random}};
  buffers_0_28_3 = _RAND_117[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{$random}};
  buffers_0_29_0 = _RAND_118[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{$random}};
  buffers_0_29_1 = _RAND_119[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{$random}};
  buffers_0_29_2 = _RAND_120[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{$random}};
  buffers_0_29_3 = _RAND_121[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{$random}};
  buffers_0_30_0 = _RAND_122[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{$random}};
  buffers_0_30_1 = _RAND_123[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{$random}};
  buffers_0_30_2 = _RAND_124[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{$random}};
  buffers_0_30_3 = _RAND_125[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{$random}};
  buffers_0_31_0 = _RAND_126[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{$random}};
  buffers_0_31_1 = _RAND_127[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{$random}};
  buffers_0_31_2 = _RAND_128[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{$random}};
  buffers_0_31_3 = _RAND_129[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{$random}};
  buffers_0_32_0 = _RAND_130[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{$random}};
  buffers_0_32_1 = _RAND_131[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{$random}};
  buffers_0_32_2 = _RAND_132[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{$random}};
  buffers_0_32_3 = _RAND_133[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{$random}};
  buffers_0_33_0 = _RAND_134[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{$random}};
  buffers_0_33_1 = _RAND_135[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{$random}};
  buffers_0_33_2 = _RAND_136[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{$random}};
  buffers_0_33_3 = _RAND_137[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{$random}};
  buffers_0_34_0 = _RAND_138[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{$random}};
  buffers_0_34_1 = _RAND_139[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{$random}};
  buffers_0_34_2 = _RAND_140[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{$random}};
  buffers_0_34_3 = _RAND_141[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{$random}};
  buffers_0_35_0 = _RAND_142[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{$random}};
  buffers_0_35_1 = _RAND_143[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{$random}};
  buffers_0_35_2 = _RAND_144[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{$random}};
  buffers_0_35_3 = _RAND_145[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{$random}};
  buffers_0_36_0 = _RAND_146[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{$random}};
  buffers_0_36_1 = _RAND_147[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{$random}};
  buffers_0_36_2 = _RAND_148[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{$random}};
  buffers_0_36_3 = _RAND_149[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{$random}};
  buffers_0_37_0 = _RAND_150[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{$random}};
  buffers_0_37_1 = _RAND_151[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{$random}};
  buffers_0_37_2 = _RAND_152[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{$random}};
  buffers_0_37_3 = _RAND_153[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{$random}};
  buffers_0_38_0 = _RAND_154[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{$random}};
  buffers_0_38_1 = _RAND_155[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{$random}};
  buffers_0_38_2 = _RAND_156[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{$random}};
  buffers_0_38_3 = _RAND_157[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{$random}};
  buffers_0_39_0 = _RAND_158[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{$random}};
  buffers_0_39_1 = _RAND_159[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{$random}};
  buffers_0_39_2 = _RAND_160[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{$random}};
  buffers_0_39_3 = _RAND_161[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{$random}};
  buffers_0_40_0 = _RAND_162[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{$random}};
  buffers_0_40_1 = _RAND_163[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{$random}};
  buffers_0_40_2 = _RAND_164[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{$random}};
  buffers_0_40_3 = _RAND_165[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{$random}};
  buffers_0_41_0 = _RAND_166[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{$random}};
  buffers_0_41_1 = _RAND_167[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{$random}};
  buffers_0_41_2 = _RAND_168[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{$random}};
  buffers_0_41_3 = _RAND_169[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{$random}};
  buffers_0_42_0 = _RAND_170[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{$random}};
  buffers_0_42_1 = _RAND_171[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{$random}};
  buffers_0_42_2 = _RAND_172[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{$random}};
  buffers_0_42_3 = _RAND_173[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{$random}};
  buffers_0_43_0 = _RAND_174[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{$random}};
  buffers_0_43_1 = _RAND_175[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{$random}};
  buffers_0_43_2 = _RAND_176[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{$random}};
  buffers_0_43_3 = _RAND_177[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{$random}};
  buffers_0_44_0 = _RAND_178[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{$random}};
  buffers_0_44_1 = _RAND_179[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{$random}};
  buffers_0_44_2 = _RAND_180[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{$random}};
  buffers_0_44_3 = _RAND_181[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{$random}};
  buffers_0_45_0 = _RAND_182[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{$random}};
  buffers_0_45_1 = _RAND_183[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{$random}};
  buffers_0_45_2 = _RAND_184[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{$random}};
  buffers_0_45_3 = _RAND_185[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{$random}};
  buffers_0_46_0 = _RAND_186[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{$random}};
  buffers_0_46_1 = _RAND_187[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{$random}};
  buffers_0_46_2 = _RAND_188[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{$random}};
  buffers_0_46_3 = _RAND_189[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{$random}};
  buffers_0_47_0 = _RAND_190[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{$random}};
  buffers_0_47_1 = _RAND_191[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{$random}};
  buffers_0_47_2 = _RAND_192[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{$random}};
  buffers_0_47_3 = _RAND_193[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{$random}};
  buffers_0_48_0 = _RAND_194[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{$random}};
  buffers_0_48_1 = _RAND_195[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{$random}};
  buffers_0_48_2 = _RAND_196[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{$random}};
  buffers_0_48_3 = _RAND_197[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{$random}};
  buffers_0_49_0 = _RAND_198[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{$random}};
  buffers_0_49_1 = _RAND_199[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{$random}};
  buffers_0_49_2 = _RAND_200[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{$random}};
  buffers_0_49_3 = _RAND_201[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{$random}};
  buffers_0_50_0 = _RAND_202[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{$random}};
  buffers_0_50_1 = _RAND_203[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{$random}};
  buffers_0_50_2 = _RAND_204[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{$random}};
  buffers_0_50_3 = _RAND_205[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{$random}};
  buffers_0_51_0 = _RAND_206[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{$random}};
  buffers_0_51_1 = _RAND_207[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{$random}};
  buffers_0_51_2 = _RAND_208[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{$random}};
  buffers_0_51_3 = _RAND_209[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{$random}};
  buffers_0_52_0 = _RAND_210[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{$random}};
  buffers_0_52_1 = _RAND_211[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{$random}};
  buffers_0_52_2 = _RAND_212[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{$random}};
  buffers_0_52_3 = _RAND_213[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{$random}};
  buffers_0_53_0 = _RAND_214[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{$random}};
  buffers_0_53_1 = _RAND_215[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{$random}};
  buffers_0_53_2 = _RAND_216[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{$random}};
  buffers_0_53_3 = _RAND_217[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{$random}};
  buffers_0_54_0 = _RAND_218[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{$random}};
  buffers_0_54_1 = _RAND_219[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{$random}};
  buffers_0_54_2 = _RAND_220[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{$random}};
  buffers_0_54_3 = _RAND_221[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{$random}};
  buffers_0_55_0 = _RAND_222[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{$random}};
  buffers_0_55_1 = _RAND_223[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{$random}};
  buffers_0_55_2 = _RAND_224[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{$random}};
  buffers_0_55_3 = _RAND_225[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{$random}};
  buffers_0_56_0 = _RAND_226[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{$random}};
  buffers_0_56_1 = _RAND_227[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{$random}};
  buffers_0_56_2 = _RAND_228[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{$random}};
  buffers_0_56_3 = _RAND_229[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{$random}};
  buffers_0_57_0 = _RAND_230[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{$random}};
  buffers_0_57_1 = _RAND_231[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{$random}};
  buffers_0_57_2 = _RAND_232[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{$random}};
  buffers_0_57_3 = _RAND_233[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{$random}};
  buffers_0_58_0 = _RAND_234[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{$random}};
  buffers_0_58_1 = _RAND_235[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{$random}};
  buffers_0_58_2 = _RAND_236[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{$random}};
  buffers_0_58_3 = _RAND_237[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{$random}};
  buffers_0_59_0 = _RAND_238[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{$random}};
  buffers_0_59_1 = _RAND_239[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{$random}};
  buffers_0_59_2 = _RAND_240[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{$random}};
  buffers_0_59_3 = _RAND_241[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{$random}};
  buffers_0_60_0 = _RAND_242[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{$random}};
  buffers_0_60_1 = _RAND_243[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{$random}};
  buffers_0_60_2 = _RAND_244[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{$random}};
  buffers_0_60_3 = _RAND_245[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{$random}};
  buffers_0_61_0 = _RAND_246[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{$random}};
  buffers_0_61_1 = _RAND_247[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{$random}};
  buffers_0_61_2 = _RAND_248[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{$random}};
  buffers_0_61_3 = _RAND_249[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{$random}};
  buffers_0_62_0 = _RAND_250[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{$random}};
  buffers_0_62_1 = _RAND_251[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{$random}};
  buffers_0_62_2 = _RAND_252[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{$random}};
  buffers_0_62_3 = _RAND_253[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{$random}};
  buffers_0_63_0 = _RAND_254[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{$random}};
  buffers_0_63_1 = _RAND_255[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{$random}};
  buffers_0_63_2 = _RAND_256[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{$random}};
  buffers_0_63_3 = _RAND_257[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{$random}};
  cntrs_0 = _RAND_258[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{$random}};
  _T_1071 = _RAND_259[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{$random}};
  cntrs_1 = _RAND_260[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{$random}};
  _T_1076 = _RAND_261[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{$random}};
  _T_1078 = _RAND_262[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{$random}};
  cntrs_2 = _RAND_263[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{$random}};
  buffers_1_0_0 = _RAND_264[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{$random}};
  buffers_1_0_1 = _RAND_265[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{$random}};
  buffers_1_0_2 = _RAND_266[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{$random}};
  buffers_1_0_3 = _RAND_267[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{$random}};
  buffers_1_1_0 = _RAND_268[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{$random}};
  buffers_1_1_1 = _RAND_269[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{$random}};
  buffers_1_1_2 = _RAND_270[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{$random}};
  buffers_1_1_3 = _RAND_271[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{$random}};
  buffers_1_2_0 = _RAND_272[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{$random}};
  buffers_1_2_1 = _RAND_273[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{$random}};
  buffers_1_2_2 = _RAND_274[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{$random}};
  buffers_1_2_3 = _RAND_275[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{$random}};
  buffers_1_3_0 = _RAND_276[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{$random}};
  buffers_1_3_1 = _RAND_277[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{$random}};
  buffers_1_3_2 = _RAND_278[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{$random}};
  buffers_1_3_3 = _RAND_279[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{$random}};
  buffers_1_4_0 = _RAND_280[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{$random}};
  buffers_1_4_1 = _RAND_281[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{$random}};
  buffers_1_4_2 = _RAND_282[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{$random}};
  buffers_1_4_3 = _RAND_283[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{$random}};
  buffers_1_5_0 = _RAND_284[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{$random}};
  buffers_1_5_1 = _RAND_285[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{$random}};
  buffers_1_5_2 = _RAND_286[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{$random}};
  buffers_1_5_3 = _RAND_287[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{$random}};
  buffers_1_6_0 = _RAND_288[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{$random}};
  buffers_1_6_1 = _RAND_289[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{$random}};
  buffers_1_6_2 = _RAND_290[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{$random}};
  buffers_1_6_3 = _RAND_291[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{$random}};
  buffers_1_7_0 = _RAND_292[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{$random}};
  buffers_1_7_1 = _RAND_293[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{$random}};
  buffers_1_7_2 = _RAND_294[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{$random}};
  buffers_1_7_3 = _RAND_295[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{$random}};
  buffers_1_8_0 = _RAND_296[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{$random}};
  buffers_1_8_1 = _RAND_297[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{$random}};
  buffers_1_8_2 = _RAND_298[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{$random}};
  buffers_1_8_3 = _RAND_299[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{$random}};
  buffers_1_9_0 = _RAND_300[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{$random}};
  buffers_1_9_1 = _RAND_301[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{$random}};
  buffers_1_9_2 = _RAND_302[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{$random}};
  buffers_1_9_3 = _RAND_303[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{$random}};
  buffers_1_10_0 = _RAND_304[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{$random}};
  buffers_1_10_1 = _RAND_305[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{$random}};
  buffers_1_10_2 = _RAND_306[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{$random}};
  buffers_1_10_3 = _RAND_307[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{$random}};
  buffers_1_11_0 = _RAND_308[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{$random}};
  buffers_1_11_1 = _RAND_309[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{$random}};
  buffers_1_11_2 = _RAND_310[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{$random}};
  buffers_1_11_3 = _RAND_311[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{$random}};
  buffers_1_12_0 = _RAND_312[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{$random}};
  buffers_1_12_1 = _RAND_313[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{$random}};
  buffers_1_12_2 = _RAND_314[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{$random}};
  buffers_1_12_3 = _RAND_315[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{$random}};
  buffers_1_13_0 = _RAND_316[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{$random}};
  buffers_1_13_1 = _RAND_317[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{$random}};
  buffers_1_13_2 = _RAND_318[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{$random}};
  buffers_1_13_3 = _RAND_319[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{$random}};
  buffers_1_14_0 = _RAND_320[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{$random}};
  buffers_1_14_1 = _RAND_321[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{$random}};
  buffers_1_14_2 = _RAND_322[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{$random}};
  buffers_1_14_3 = _RAND_323[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{$random}};
  buffers_1_15_0 = _RAND_324[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{$random}};
  buffers_1_15_1 = _RAND_325[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{$random}};
  buffers_1_15_2 = _RAND_326[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{$random}};
  buffers_1_15_3 = _RAND_327[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{$random}};
  buffers_2_0_0 = _RAND_328[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{$random}};
  buffers_2_0_1 = _RAND_329[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{$random}};
  buffers_2_0_2 = _RAND_330[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{$random}};
  buffers_2_0_3 = _RAND_331[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{$random}};
  buffers_2_1_0 = _RAND_332[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{$random}};
  buffers_2_1_1 = _RAND_333[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{$random}};
  buffers_2_1_2 = _RAND_334[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{$random}};
  buffers_2_1_3 = _RAND_335[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{$random}};
  buffers_2_2_0 = _RAND_336[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{$random}};
  buffers_2_2_1 = _RAND_337[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{$random}};
  buffers_2_2_2 = _RAND_338[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{$random}};
  buffers_2_2_3 = _RAND_339[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{$random}};
  buffers_2_3_0 = _RAND_340[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{$random}};
  buffers_2_3_1 = _RAND_341[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{$random}};
  buffers_2_3_2 = _RAND_342[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{$random}};
  buffers_2_3_3 = _RAND_343[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{$random}};
  buffers_3_0_0 = _RAND_344[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{$random}};
  buffers_3_0_1 = _RAND_345[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{$random}};
  buffers_3_0_2 = _RAND_346[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{$random}};
  buffers_3_0_3 = _RAND_347[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{$random}};
  _T_1988 = _RAND_348[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{$random}};
  _T_1990 = _RAND_349[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{$random}};
  vld = _RAND_350[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{$random}};
  lastVld = _RAND_351[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      rdyReg <= 1'h1;
    end else begin
      if (_T_1063) begin
        rdyReg <= 1'h0;
      end else begin
        if (_T_1061) begin
          rdyReg <= 1'h1;
        end
      end
    end
    if (reset) begin
      cntr <= 6'h0;
    end else begin
      if (_T_1058) begin
        cntr <= 6'h1;
      end else begin
        if (_T_1052) begin
          cntr <= _T_1055;
        end
      end
    end
    if (_T_1058) begin
      buffers_0_0_0 <= io_dataIn_bits_0;
    end
    if (_T_1058) begin
      buffers_0_0_1 <= io_dataIn_bits_1;
    end
    if (_T_1058) begin
      buffers_0_0_2 <= io_dataIn_bits_2;
    end
    if (_T_1058) begin
      buffers_0_0_3 <= io_dataIn_bits_3;
    end
    if (_T_1058) begin
      buffers_0_1_0 <= io_dataIn_bits_4;
    end
    if (_T_1058) begin
      buffers_0_1_1 <= io_dataIn_bits_5;
    end
    if (_T_1058) begin
      buffers_0_1_2 <= io_dataIn_bits_6;
    end
    if (_T_1058) begin
      buffers_0_1_3 <= io_dataIn_bits_7;
    end
    if (_T_1058) begin
      buffers_0_2_0 <= io_dataIn_bits_8;
    end
    if (_T_1058) begin
      buffers_0_2_1 <= io_dataIn_bits_9;
    end
    if (_T_1058) begin
      buffers_0_2_2 <= io_dataIn_bits_10;
    end
    if (_T_1058) begin
      buffers_0_2_3 <= io_dataIn_bits_11;
    end
    if (_T_1058) begin
      buffers_0_3_0 <= io_dataIn_bits_12;
    end
    if (_T_1058) begin
      buffers_0_3_1 <= io_dataIn_bits_13;
    end
    if (_T_1058) begin
      buffers_0_3_2 <= io_dataIn_bits_14;
    end
    if (_T_1058) begin
      buffers_0_3_3 <= io_dataIn_bits_15;
    end
    if (_T_1058) begin
      buffers_0_4_0 <= io_dataIn_bits_16;
    end
    if (_T_1058) begin
      buffers_0_4_1 <= io_dataIn_bits_17;
    end
    if (_T_1058) begin
      buffers_0_4_2 <= io_dataIn_bits_18;
    end
    if (_T_1058) begin
      buffers_0_4_3 <= io_dataIn_bits_19;
    end
    if (_T_1058) begin
      buffers_0_5_0 <= io_dataIn_bits_20;
    end
    if (_T_1058) begin
      buffers_0_5_1 <= io_dataIn_bits_21;
    end
    if (_T_1058) begin
      buffers_0_5_2 <= io_dataIn_bits_22;
    end
    if (_T_1058) begin
      buffers_0_5_3 <= io_dataIn_bits_23;
    end
    if (_T_1058) begin
      buffers_0_6_0 <= io_dataIn_bits_24;
    end
    if (_T_1058) begin
      buffers_0_6_1 <= io_dataIn_bits_25;
    end
    if (_T_1058) begin
      buffers_0_6_2 <= io_dataIn_bits_26;
    end
    if (_T_1058) begin
      buffers_0_6_3 <= io_dataIn_bits_27;
    end
    if (_T_1058) begin
      buffers_0_7_0 <= io_dataIn_bits_28;
    end
    if (_T_1058) begin
      buffers_0_7_1 <= io_dataIn_bits_29;
    end
    if (_T_1058) begin
      buffers_0_7_2 <= io_dataIn_bits_30;
    end
    if (_T_1058) begin
      buffers_0_7_3 <= io_dataIn_bits_31;
    end
    if (_T_1058) begin
      buffers_0_8_0 <= io_dataIn_bits_32;
    end
    if (_T_1058) begin
      buffers_0_8_1 <= io_dataIn_bits_33;
    end
    if (_T_1058) begin
      buffers_0_8_2 <= io_dataIn_bits_34;
    end
    if (_T_1058) begin
      buffers_0_8_3 <= io_dataIn_bits_35;
    end
    if (_T_1058) begin
      buffers_0_9_0 <= io_dataIn_bits_36;
    end
    if (_T_1058) begin
      buffers_0_9_1 <= io_dataIn_bits_37;
    end
    if (_T_1058) begin
      buffers_0_9_2 <= io_dataIn_bits_38;
    end
    if (_T_1058) begin
      buffers_0_9_3 <= io_dataIn_bits_39;
    end
    if (_T_1058) begin
      buffers_0_10_0 <= io_dataIn_bits_40;
    end
    if (_T_1058) begin
      buffers_0_10_1 <= io_dataIn_bits_41;
    end
    if (_T_1058) begin
      buffers_0_10_2 <= io_dataIn_bits_42;
    end
    if (_T_1058) begin
      buffers_0_10_3 <= io_dataIn_bits_43;
    end
    if (_T_1058) begin
      buffers_0_11_0 <= io_dataIn_bits_44;
    end
    if (_T_1058) begin
      buffers_0_11_1 <= io_dataIn_bits_45;
    end
    if (_T_1058) begin
      buffers_0_11_2 <= io_dataIn_bits_46;
    end
    if (_T_1058) begin
      buffers_0_11_3 <= io_dataIn_bits_47;
    end
    if (_T_1058) begin
      buffers_0_12_0 <= io_dataIn_bits_48;
    end
    if (_T_1058) begin
      buffers_0_12_1 <= io_dataIn_bits_49;
    end
    if (_T_1058) begin
      buffers_0_12_2 <= io_dataIn_bits_50;
    end
    if (_T_1058) begin
      buffers_0_12_3 <= io_dataIn_bits_51;
    end
    if (_T_1058) begin
      buffers_0_13_0 <= io_dataIn_bits_52;
    end
    if (_T_1058) begin
      buffers_0_13_1 <= io_dataIn_bits_53;
    end
    if (_T_1058) begin
      buffers_0_13_2 <= io_dataIn_bits_54;
    end
    if (_T_1058) begin
      buffers_0_13_3 <= io_dataIn_bits_55;
    end
    if (_T_1058) begin
      buffers_0_14_0 <= io_dataIn_bits_56;
    end
    if (_T_1058) begin
      buffers_0_14_1 <= io_dataIn_bits_57;
    end
    if (_T_1058) begin
      buffers_0_14_2 <= io_dataIn_bits_58;
    end
    if (_T_1058) begin
      buffers_0_14_3 <= io_dataIn_bits_59;
    end
    if (_T_1058) begin
      buffers_0_15_0 <= io_dataIn_bits_60;
    end
    if (_T_1058) begin
      buffers_0_15_1 <= io_dataIn_bits_61;
    end
    if (_T_1058) begin
      buffers_0_15_2 <= io_dataIn_bits_62;
    end
    if (_T_1058) begin
      buffers_0_15_3 <= io_dataIn_bits_63;
    end
    if (_T_1058) begin
      buffers_0_16_0 <= io_dataIn_bits_64;
    end
    if (_T_1058) begin
      buffers_0_16_1 <= io_dataIn_bits_65;
    end
    if (_T_1058) begin
      buffers_0_16_2 <= io_dataIn_bits_66;
    end
    if (_T_1058) begin
      buffers_0_16_3 <= io_dataIn_bits_67;
    end
    if (_T_1058) begin
      buffers_0_17_0 <= io_dataIn_bits_68;
    end
    if (_T_1058) begin
      buffers_0_17_1 <= io_dataIn_bits_69;
    end
    if (_T_1058) begin
      buffers_0_17_2 <= io_dataIn_bits_70;
    end
    if (_T_1058) begin
      buffers_0_17_3 <= io_dataIn_bits_71;
    end
    if (_T_1058) begin
      buffers_0_18_0 <= io_dataIn_bits_72;
    end
    if (_T_1058) begin
      buffers_0_18_1 <= io_dataIn_bits_73;
    end
    if (_T_1058) begin
      buffers_0_18_2 <= io_dataIn_bits_74;
    end
    if (_T_1058) begin
      buffers_0_18_3 <= io_dataIn_bits_75;
    end
    if (_T_1058) begin
      buffers_0_19_0 <= io_dataIn_bits_76;
    end
    if (_T_1058) begin
      buffers_0_19_1 <= io_dataIn_bits_77;
    end
    if (_T_1058) begin
      buffers_0_19_2 <= io_dataIn_bits_78;
    end
    if (_T_1058) begin
      buffers_0_19_3 <= io_dataIn_bits_79;
    end
    if (_T_1058) begin
      buffers_0_20_0 <= io_dataIn_bits_80;
    end
    if (_T_1058) begin
      buffers_0_20_1 <= io_dataIn_bits_81;
    end
    if (_T_1058) begin
      buffers_0_20_2 <= io_dataIn_bits_82;
    end
    if (_T_1058) begin
      buffers_0_20_3 <= io_dataIn_bits_83;
    end
    if (_T_1058) begin
      buffers_0_21_0 <= io_dataIn_bits_84;
    end
    if (_T_1058) begin
      buffers_0_21_1 <= io_dataIn_bits_85;
    end
    if (_T_1058) begin
      buffers_0_21_2 <= io_dataIn_bits_86;
    end
    if (_T_1058) begin
      buffers_0_21_3 <= io_dataIn_bits_87;
    end
    if (_T_1058) begin
      buffers_0_22_0 <= io_dataIn_bits_88;
    end
    if (_T_1058) begin
      buffers_0_22_1 <= io_dataIn_bits_89;
    end
    if (_T_1058) begin
      buffers_0_22_2 <= io_dataIn_bits_90;
    end
    if (_T_1058) begin
      buffers_0_22_3 <= io_dataIn_bits_91;
    end
    if (_T_1058) begin
      buffers_0_23_0 <= io_dataIn_bits_92;
    end
    if (_T_1058) begin
      buffers_0_23_1 <= io_dataIn_bits_93;
    end
    if (_T_1058) begin
      buffers_0_23_2 <= io_dataIn_bits_94;
    end
    if (_T_1058) begin
      buffers_0_23_3 <= io_dataIn_bits_95;
    end
    if (_T_1058) begin
      buffers_0_24_0 <= io_dataIn_bits_96;
    end
    if (_T_1058) begin
      buffers_0_24_1 <= io_dataIn_bits_97;
    end
    if (_T_1058) begin
      buffers_0_24_2 <= io_dataIn_bits_98;
    end
    if (_T_1058) begin
      buffers_0_24_3 <= io_dataIn_bits_99;
    end
    if (_T_1058) begin
      buffers_0_25_0 <= io_dataIn_bits_100;
    end
    if (_T_1058) begin
      buffers_0_25_1 <= io_dataIn_bits_101;
    end
    if (_T_1058) begin
      buffers_0_25_2 <= io_dataIn_bits_102;
    end
    if (_T_1058) begin
      buffers_0_25_3 <= io_dataIn_bits_103;
    end
    if (_T_1058) begin
      buffers_0_26_0 <= io_dataIn_bits_104;
    end
    if (_T_1058) begin
      buffers_0_26_1 <= io_dataIn_bits_105;
    end
    if (_T_1058) begin
      buffers_0_26_2 <= io_dataIn_bits_106;
    end
    if (_T_1058) begin
      buffers_0_26_3 <= io_dataIn_bits_107;
    end
    if (_T_1058) begin
      buffers_0_27_0 <= io_dataIn_bits_108;
    end
    if (_T_1058) begin
      buffers_0_27_1 <= io_dataIn_bits_109;
    end
    if (_T_1058) begin
      buffers_0_27_2 <= io_dataIn_bits_110;
    end
    if (_T_1058) begin
      buffers_0_27_3 <= io_dataIn_bits_111;
    end
    if (_T_1058) begin
      buffers_0_28_0 <= io_dataIn_bits_112;
    end
    if (_T_1058) begin
      buffers_0_28_1 <= io_dataIn_bits_113;
    end
    if (_T_1058) begin
      buffers_0_28_2 <= io_dataIn_bits_114;
    end
    if (_T_1058) begin
      buffers_0_28_3 <= io_dataIn_bits_115;
    end
    if (_T_1058) begin
      buffers_0_29_0 <= io_dataIn_bits_116;
    end
    if (_T_1058) begin
      buffers_0_29_1 <= io_dataIn_bits_117;
    end
    if (_T_1058) begin
      buffers_0_29_2 <= io_dataIn_bits_118;
    end
    if (_T_1058) begin
      buffers_0_29_3 <= io_dataIn_bits_119;
    end
    if (_T_1058) begin
      buffers_0_30_0 <= io_dataIn_bits_120;
    end
    if (_T_1058) begin
      buffers_0_30_1 <= io_dataIn_bits_121;
    end
    if (_T_1058) begin
      buffers_0_30_2 <= io_dataIn_bits_122;
    end
    if (_T_1058) begin
      buffers_0_30_3 <= io_dataIn_bits_123;
    end
    if (_T_1058) begin
      buffers_0_31_0 <= io_dataIn_bits_124;
    end
    if (_T_1058) begin
      buffers_0_31_1 <= io_dataIn_bits_125;
    end
    if (_T_1058) begin
      buffers_0_31_2 <= io_dataIn_bits_126;
    end
    if (_T_1058) begin
      buffers_0_31_3 <= io_dataIn_bits_127;
    end
    if (_T_1058) begin
      buffers_0_32_0 <= io_dataIn_bits_128;
    end
    if (_T_1058) begin
      buffers_0_32_1 <= io_dataIn_bits_129;
    end
    if (_T_1058) begin
      buffers_0_32_2 <= io_dataIn_bits_130;
    end
    if (_T_1058) begin
      buffers_0_32_3 <= io_dataIn_bits_131;
    end
    if (_T_1058) begin
      buffers_0_33_0 <= io_dataIn_bits_132;
    end
    if (_T_1058) begin
      buffers_0_33_1 <= io_dataIn_bits_133;
    end
    if (_T_1058) begin
      buffers_0_33_2 <= io_dataIn_bits_134;
    end
    if (_T_1058) begin
      buffers_0_33_3 <= io_dataIn_bits_135;
    end
    if (_T_1058) begin
      buffers_0_34_0 <= io_dataIn_bits_136;
    end
    if (_T_1058) begin
      buffers_0_34_1 <= io_dataIn_bits_137;
    end
    if (_T_1058) begin
      buffers_0_34_2 <= io_dataIn_bits_138;
    end
    if (_T_1058) begin
      buffers_0_34_3 <= io_dataIn_bits_139;
    end
    if (_T_1058) begin
      buffers_0_35_0 <= io_dataIn_bits_140;
    end
    if (_T_1058) begin
      buffers_0_35_1 <= io_dataIn_bits_141;
    end
    if (_T_1058) begin
      buffers_0_35_2 <= io_dataIn_bits_142;
    end
    if (_T_1058) begin
      buffers_0_35_3 <= io_dataIn_bits_143;
    end
    if (_T_1058) begin
      buffers_0_36_0 <= io_dataIn_bits_144;
    end
    if (_T_1058) begin
      buffers_0_36_1 <= io_dataIn_bits_145;
    end
    if (_T_1058) begin
      buffers_0_36_2 <= io_dataIn_bits_146;
    end
    if (_T_1058) begin
      buffers_0_36_3 <= io_dataIn_bits_147;
    end
    if (_T_1058) begin
      buffers_0_37_0 <= io_dataIn_bits_148;
    end
    if (_T_1058) begin
      buffers_0_37_1 <= io_dataIn_bits_149;
    end
    if (_T_1058) begin
      buffers_0_37_2 <= io_dataIn_bits_150;
    end
    if (_T_1058) begin
      buffers_0_37_3 <= io_dataIn_bits_151;
    end
    if (_T_1058) begin
      buffers_0_38_0 <= io_dataIn_bits_152;
    end
    if (_T_1058) begin
      buffers_0_38_1 <= io_dataIn_bits_153;
    end
    if (_T_1058) begin
      buffers_0_38_2 <= io_dataIn_bits_154;
    end
    if (_T_1058) begin
      buffers_0_38_3 <= io_dataIn_bits_155;
    end
    if (_T_1058) begin
      buffers_0_39_0 <= io_dataIn_bits_156;
    end
    if (_T_1058) begin
      buffers_0_39_1 <= io_dataIn_bits_157;
    end
    if (_T_1058) begin
      buffers_0_39_2 <= io_dataIn_bits_158;
    end
    if (_T_1058) begin
      buffers_0_39_3 <= io_dataIn_bits_159;
    end
    if (_T_1058) begin
      buffers_0_40_0 <= io_dataIn_bits_160;
    end
    if (_T_1058) begin
      buffers_0_40_1 <= io_dataIn_bits_161;
    end
    if (_T_1058) begin
      buffers_0_40_2 <= io_dataIn_bits_162;
    end
    if (_T_1058) begin
      buffers_0_40_3 <= io_dataIn_bits_163;
    end
    if (_T_1058) begin
      buffers_0_41_0 <= io_dataIn_bits_164;
    end
    if (_T_1058) begin
      buffers_0_41_1 <= io_dataIn_bits_165;
    end
    if (_T_1058) begin
      buffers_0_41_2 <= io_dataIn_bits_166;
    end
    if (_T_1058) begin
      buffers_0_41_3 <= io_dataIn_bits_167;
    end
    if (_T_1058) begin
      buffers_0_42_0 <= io_dataIn_bits_168;
    end
    if (_T_1058) begin
      buffers_0_42_1 <= io_dataIn_bits_169;
    end
    if (_T_1058) begin
      buffers_0_42_2 <= io_dataIn_bits_170;
    end
    if (_T_1058) begin
      buffers_0_42_3 <= io_dataIn_bits_171;
    end
    if (_T_1058) begin
      buffers_0_43_0 <= io_dataIn_bits_172;
    end
    if (_T_1058) begin
      buffers_0_43_1 <= io_dataIn_bits_173;
    end
    if (_T_1058) begin
      buffers_0_43_2 <= io_dataIn_bits_174;
    end
    if (_T_1058) begin
      buffers_0_43_3 <= io_dataIn_bits_175;
    end
    if (_T_1058) begin
      buffers_0_44_0 <= io_dataIn_bits_176;
    end
    if (_T_1058) begin
      buffers_0_44_1 <= io_dataIn_bits_177;
    end
    if (_T_1058) begin
      buffers_0_44_2 <= io_dataIn_bits_178;
    end
    if (_T_1058) begin
      buffers_0_44_3 <= io_dataIn_bits_179;
    end
    if (_T_1058) begin
      buffers_0_45_0 <= io_dataIn_bits_180;
    end
    if (_T_1058) begin
      buffers_0_45_1 <= io_dataIn_bits_181;
    end
    if (_T_1058) begin
      buffers_0_45_2 <= io_dataIn_bits_182;
    end
    if (_T_1058) begin
      buffers_0_45_3 <= io_dataIn_bits_183;
    end
    if (_T_1058) begin
      buffers_0_46_0 <= io_dataIn_bits_184;
    end
    if (_T_1058) begin
      buffers_0_46_1 <= io_dataIn_bits_185;
    end
    if (_T_1058) begin
      buffers_0_46_2 <= io_dataIn_bits_186;
    end
    if (_T_1058) begin
      buffers_0_46_3 <= io_dataIn_bits_187;
    end
    if (_T_1058) begin
      buffers_0_47_0 <= io_dataIn_bits_188;
    end
    if (_T_1058) begin
      buffers_0_47_1 <= io_dataIn_bits_189;
    end
    if (_T_1058) begin
      buffers_0_47_2 <= io_dataIn_bits_190;
    end
    if (_T_1058) begin
      buffers_0_47_3 <= io_dataIn_bits_191;
    end
    if (_T_1058) begin
      buffers_0_48_0 <= io_dataIn_bits_192;
    end
    if (_T_1058) begin
      buffers_0_48_1 <= io_dataIn_bits_193;
    end
    if (_T_1058) begin
      buffers_0_48_2 <= io_dataIn_bits_194;
    end
    if (_T_1058) begin
      buffers_0_48_3 <= io_dataIn_bits_195;
    end
    if (_T_1058) begin
      buffers_0_49_0 <= io_dataIn_bits_196;
    end
    if (_T_1058) begin
      buffers_0_49_1 <= io_dataIn_bits_197;
    end
    if (_T_1058) begin
      buffers_0_49_2 <= io_dataIn_bits_198;
    end
    if (_T_1058) begin
      buffers_0_49_3 <= io_dataIn_bits_199;
    end
    if (_T_1058) begin
      buffers_0_50_0 <= io_dataIn_bits_200;
    end
    if (_T_1058) begin
      buffers_0_50_1 <= io_dataIn_bits_201;
    end
    if (_T_1058) begin
      buffers_0_50_2 <= io_dataIn_bits_202;
    end
    if (_T_1058) begin
      buffers_0_50_3 <= io_dataIn_bits_203;
    end
    if (_T_1058) begin
      buffers_0_51_0 <= io_dataIn_bits_204;
    end
    if (_T_1058) begin
      buffers_0_51_1 <= io_dataIn_bits_205;
    end
    if (_T_1058) begin
      buffers_0_51_2 <= io_dataIn_bits_206;
    end
    if (_T_1058) begin
      buffers_0_51_3 <= io_dataIn_bits_207;
    end
    if (_T_1058) begin
      buffers_0_52_0 <= io_dataIn_bits_208;
    end
    if (_T_1058) begin
      buffers_0_52_1 <= io_dataIn_bits_209;
    end
    if (_T_1058) begin
      buffers_0_52_2 <= io_dataIn_bits_210;
    end
    if (_T_1058) begin
      buffers_0_52_3 <= io_dataIn_bits_211;
    end
    if (_T_1058) begin
      buffers_0_53_0 <= io_dataIn_bits_212;
    end
    if (_T_1058) begin
      buffers_0_53_1 <= io_dataIn_bits_213;
    end
    if (_T_1058) begin
      buffers_0_53_2 <= io_dataIn_bits_214;
    end
    if (_T_1058) begin
      buffers_0_53_3 <= io_dataIn_bits_215;
    end
    if (_T_1058) begin
      buffers_0_54_0 <= io_dataIn_bits_216;
    end
    if (_T_1058) begin
      buffers_0_54_1 <= io_dataIn_bits_217;
    end
    if (_T_1058) begin
      buffers_0_54_2 <= io_dataIn_bits_218;
    end
    if (_T_1058) begin
      buffers_0_54_3 <= io_dataIn_bits_219;
    end
    if (_T_1058) begin
      buffers_0_55_0 <= io_dataIn_bits_220;
    end
    if (_T_1058) begin
      buffers_0_55_1 <= io_dataIn_bits_221;
    end
    if (_T_1058) begin
      buffers_0_55_2 <= io_dataIn_bits_222;
    end
    if (_T_1058) begin
      buffers_0_55_3 <= io_dataIn_bits_223;
    end
    if (_T_1058) begin
      buffers_0_56_0 <= io_dataIn_bits_224;
    end
    if (_T_1058) begin
      buffers_0_56_1 <= io_dataIn_bits_225;
    end
    if (_T_1058) begin
      buffers_0_56_2 <= io_dataIn_bits_226;
    end
    if (_T_1058) begin
      buffers_0_56_3 <= io_dataIn_bits_227;
    end
    if (_T_1058) begin
      buffers_0_57_0 <= io_dataIn_bits_228;
    end
    if (_T_1058) begin
      buffers_0_57_1 <= io_dataIn_bits_229;
    end
    if (_T_1058) begin
      buffers_0_57_2 <= io_dataIn_bits_230;
    end
    if (_T_1058) begin
      buffers_0_57_3 <= io_dataIn_bits_231;
    end
    if (_T_1058) begin
      buffers_0_58_0 <= io_dataIn_bits_232;
    end
    if (_T_1058) begin
      buffers_0_58_1 <= io_dataIn_bits_233;
    end
    if (_T_1058) begin
      buffers_0_58_2 <= io_dataIn_bits_234;
    end
    if (_T_1058) begin
      buffers_0_58_3 <= io_dataIn_bits_235;
    end
    if (_T_1058) begin
      buffers_0_59_0 <= io_dataIn_bits_236;
    end
    if (_T_1058) begin
      buffers_0_59_1 <= io_dataIn_bits_237;
    end
    if (_T_1058) begin
      buffers_0_59_2 <= io_dataIn_bits_238;
    end
    if (_T_1058) begin
      buffers_0_59_3 <= io_dataIn_bits_239;
    end
    if (_T_1058) begin
      buffers_0_60_0 <= io_dataIn_bits_240;
    end
    if (_T_1058) begin
      buffers_0_60_1 <= io_dataIn_bits_241;
    end
    if (_T_1058) begin
      buffers_0_60_2 <= io_dataIn_bits_242;
    end
    if (_T_1058) begin
      buffers_0_60_3 <= io_dataIn_bits_243;
    end
    if (_T_1058) begin
      buffers_0_61_0 <= io_dataIn_bits_244;
    end
    if (_T_1058) begin
      buffers_0_61_1 <= io_dataIn_bits_245;
    end
    if (_T_1058) begin
      buffers_0_61_2 <= io_dataIn_bits_246;
    end
    if (_T_1058) begin
      buffers_0_61_3 <= io_dataIn_bits_247;
    end
    if (_T_1058) begin
      buffers_0_62_0 <= io_dataIn_bits_248;
    end
    if (_T_1058) begin
      buffers_0_62_1 <= io_dataIn_bits_249;
    end
    if (_T_1058) begin
      buffers_0_62_2 <= io_dataIn_bits_250;
    end
    if (_T_1058) begin
      buffers_0_62_3 <= io_dataIn_bits_251;
    end
    if (_T_1058) begin
      buffers_0_63_0 <= io_dataIn_bits_252;
    end
    if (_T_1058) begin
      buffers_0_63_1 <= io_dataIn_bits_253;
    end
    if (_T_1058) begin
      buffers_0_63_2 <= io_dataIn_bits_254;
    end
    if (_T_1058) begin
      buffers_0_63_3 <= io_dataIn_bits_255;
    end
    cntrs_0 <= _T_1065;
    _T_1071 <= _T_1068;
    cntrs_1 <= _T_1071;
    _T_1076 <= _T_1073;
    _T_1078 <= _T_1076;
    cntrs_2 <= _T_1078;
    if (_T_1094) begin
      buffers_1_0_0 <= buffers_0_3_0;
    end else begin
      if (_T_1092) begin
        buffers_1_0_0 <= buffers_0_2_0;
      end else begin
        if (_T_1090) begin
          buffers_1_0_0 <= buffers_0_1_0;
        end else begin
          buffers_1_0_0 <= buffers_0_0_0;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_0_1 <= buffers_0_3_1;
    end else begin
      if (_T_1092) begin
        buffers_1_0_1 <= buffers_0_2_1;
      end else begin
        if (_T_1090) begin
          buffers_1_0_1 <= buffers_0_1_1;
        end else begin
          buffers_1_0_1 <= buffers_0_0_1;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_0_2 <= buffers_0_3_2;
    end else begin
      if (_T_1092) begin
        buffers_1_0_2 <= buffers_0_2_2;
      end else begin
        if (_T_1090) begin
          buffers_1_0_2 <= buffers_0_1_2;
        end else begin
          buffers_1_0_2 <= buffers_0_0_2;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_0_3 <= buffers_0_3_3;
    end else begin
      if (_T_1092) begin
        buffers_1_0_3 <= buffers_0_2_3;
      end else begin
        if (_T_1090) begin
          buffers_1_0_3 <= buffers_0_1_3;
        end else begin
          buffers_1_0_3 <= buffers_0_0_3;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_1_0 <= buffers_0_7_0;
    end else begin
      if (_T_1092) begin
        buffers_1_1_0 <= buffers_0_6_0;
      end else begin
        if (_T_1090) begin
          buffers_1_1_0 <= buffers_0_5_0;
        end else begin
          buffers_1_1_0 <= buffers_0_4_0;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_1_1 <= buffers_0_7_1;
    end else begin
      if (_T_1092) begin
        buffers_1_1_1 <= buffers_0_6_1;
      end else begin
        if (_T_1090) begin
          buffers_1_1_1 <= buffers_0_5_1;
        end else begin
          buffers_1_1_1 <= buffers_0_4_1;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_1_2 <= buffers_0_7_2;
    end else begin
      if (_T_1092) begin
        buffers_1_1_2 <= buffers_0_6_2;
      end else begin
        if (_T_1090) begin
          buffers_1_1_2 <= buffers_0_5_2;
        end else begin
          buffers_1_1_2 <= buffers_0_4_2;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_1_3 <= buffers_0_7_3;
    end else begin
      if (_T_1092) begin
        buffers_1_1_3 <= buffers_0_6_3;
      end else begin
        if (_T_1090) begin
          buffers_1_1_3 <= buffers_0_5_3;
        end else begin
          buffers_1_1_3 <= buffers_0_4_3;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_2_0 <= buffers_0_11_0;
    end else begin
      if (_T_1092) begin
        buffers_1_2_0 <= buffers_0_10_0;
      end else begin
        if (_T_1090) begin
          buffers_1_2_0 <= buffers_0_9_0;
        end else begin
          buffers_1_2_0 <= buffers_0_8_0;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_2_1 <= buffers_0_11_1;
    end else begin
      if (_T_1092) begin
        buffers_1_2_1 <= buffers_0_10_1;
      end else begin
        if (_T_1090) begin
          buffers_1_2_1 <= buffers_0_9_1;
        end else begin
          buffers_1_2_1 <= buffers_0_8_1;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_2_2 <= buffers_0_11_2;
    end else begin
      if (_T_1092) begin
        buffers_1_2_2 <= buffers_0_10_2;
      end else begin
        if (_T_1090) begin
          buffers_1_2_2 <= buffers_0_9_2;
        end else begin
          buffers_1_2_2 <= buffers_0_8_2;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_2_3 <= buffers_0_11_3;
    end else begin
      if (_T_1092) begin
        buffers_1_2_3 <= buffers_0_10_3;
      end else begin
        if (_T_1090) begin
          buffers_1_2_3 <= buffers_0_9_3;
        end else begin
          buffers_1_2_3 <= buffers_0_8_3;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_3_0 <= buffers_0_15_0;
    end else begin
      if (_T_1092) begin
        buffers_1_3_0 <= buffers_0_14_0;
      end else begin
        if (_T_1090) begin
          buffers_1_3_0 <= buffers_0_13_0;
        end else begin
          buffers_1_3_0 <= buffers_0_12_0;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_3_1 <= buffers_0_15_1;
    end else begin
      if (_T_1092) begin
        buffers_1_3_1 <= buffers_0_14_1;
      end else begin
        if (_T_1090) begin
          buffers_1_3_1 <= buffers_0_13_1;
        end else begin
          buffers_1_3_1 <= buffers_0_12_1;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_3_2 <= buffers_0_15_2;
    end else begin
      if (_T_1092) begin
        buffers_1_3_2 <= buffers_0_14_2;
      end else begin
        if (_T_1090) begin
          buffers_1_3_2 <= buffers_0_13_2;
        end else begin
          buffers_1_3_2 <= buffers_0_12_2;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_3_3 <= buffers_0_15_3;
    end else begin
      if (_T_1092) begin
        buffers_1_3_3 <= buffers_0_14_3;
      end else begin
        if (_T_1090) begin
          buffers_1_3_3 <= buffers_0_13_3;
        end else begin
          buffers_1_3_3 <= buffers_0_12_3;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_4_0 <= buffers_0_19_0;
    end else begin
      if (_T_1092) begin
        buffers_1_4_0 <= buffers_0_18_0;
      end else begin
        if (_T_1090) begin
          buffers_1_4_0 <= buffers_0_17_0;
        end else begin
          buffers_1_4_0 <= buffers_0_16_0;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_4_1 <= buffers_0_19_1;
    end else begin
      if (_T_1092) begin
        buffers_1_4_1 <= buffers_0_18_1;
      end else begin
        if (_T_1090) begin
          buffers_1_4_1 <= buffers_0_17_1;
        end else begin
          buffers_1_4_1 <= buffers_0_16_1;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_4_2 <= buffers_0_19_2;
    end else begin
      if (_T_1092) begin
        buffers_1_4_2 <= buffers_0_18_2;
      end else begin
        if (_T_1090) begin
          buffers_1_4_2 <= buffers_0_17_2;
        end else begin
          buffers_1_4_2 <= buffers_0_16_2;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_4_3 <= buffers_0_19_3;
    end else begin
      if (_T_1092) begin
        buffers_1_4_3 <= buffers_0_18_3;
      end else begin
        if (_T_1090) begin
          buffers_1_4_3 <= buffers_0_17_3;
        end else begin
          buffers_1_4_3 <= buffers_0_16_3;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_5_0 <= buffers_0_23_0;
    end else begin
      if (_T_1092) begin
        buffers_1_5_0 <= buffers_0_22_0;
      end else begin
        if (_T_1090) begin
          buffers_1_5_0 <= buffers_0_21_0;
        end else begin
          buffers_1_5_0 <= buffers_0_20_0;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_5_1 <= buffers_0_23_1;
    end else begin
      if (_T_1092) begin
        buffers_1_5_1 <= buffers_0_22_1;
      end else begin
        if (_T_1090) begin
          buffers_1_5_1 <= buffers_0_21_1;
        end else begin
          buffers_1_5_1 <= buffers_0_20_1;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_5_2 <= buffers_0_23_2;
    end else begin
      if (_T_1092) begin
        buffers_1_5_2 <= buffers_0_22_2;
      end else begin
        if (_T_1090) begin
          buffers_1_5_2 <= buffers_0_21_2;
        end else begin
          buffers_1_5_2 <= buffers_0_20_2;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_5_3 <= buffers_0_23_3;
    end else begin
      if (_T_1092) begin
        buffers_1_5_3 <= buffers_0_22_3;
      end else begin
        if (_T_1090) begin
          buffers_1_5_3 <= buffers_0_21_3;
        end else begin
          buffers_1_5_3 <= buffers_0_20_3;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_6_0 <= buffers_0_27_0;
    end else begin
      if (_T_1092) begin
        buffers_1_6_0 <= buffers_0_26_0;
      end else begin
        if (_T_1090) begin
          buffers_1_6_0 <= buffers_0_25_0;
        end else begin
          buffers_1_6_0 <= buffers_0_24_0;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_6_1 <= buffers_0_27_1;
    end else begin
      if (_T_1092) begin
        buffers_1_6_1 <= buffers_0_26_1;
      end else begin
        if (_T_1090) begin
          buffers_1_6_1 <= buffers_0_25_1;
        end else begin
          buffers_1_6_1 <= buffers_0_24_1;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_6_2 <= buffers_0_27_2;
    end else begin
      if (_T_1092) begin
        buffers_1_6_2 <= buffers_0_26_2;
      end else begin
        if (_T_1090) begin
          buffers_1_6_2 <= buffers_0_25_2;
        end else begin
          buffers_1_6_2 <= buffers_0_24_2;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_6_3 <= buffers_0_27_3;
    end else begin
      if (_T_1092) begin
        buffers_1_6_3 <= buffers_0_26_3;
      end else begin
        if (_T_1090) begin
          buffers_1_6_3 <= buffers_0_25_3;
        end else begin
          buffers_1_6_3 <= buffers_0_24_3;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_7_0 <= buffers_0_31_0;
    end else begin
      if (_T_1092) begin
        buffers_1_7_0 <= buffers_0_30_0;
      end else begin
        if (_T_1090) begin
          buffers_1_7_0 <= buffers_0_29_0;
        end else begin
          buffers_1_7_0 <= buffers_0_28_0;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_7_1 <= buffers_0_31_1;
    end else begin
      if (_T_1092) begin
        buffers_1_7_1 <= buffers_0_30_1;
      end else begin
        if (_T_1090) begin
          buffers_1_7_1 <= buffers_0_29_1;
        end else begin
          buffers_1_7_1 <= buffers_0_28_1;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_7_2 <= buffers_0_31_2;
    end else begin
      if (_T_1092) begin
        buffers_1_7_2 <= buffers_0_30_2;
      end else begin
        if (_T_1090) begin
          buffers_1_7_2 <= buffers_0_29_2;
        end else begin
          buffers_1_7_2 <= buffers_0_28_2;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_7_3 <= buffers_0_31_3;
    end else begin
      if (_T_1092) begin
        buffers_1_7_3 <= buffers_0_30_3;
      end else begin
        if (_T_1090) begin
          buffers_1_7_3 <= buffers_0_29_3;
        end else begin
          buffers_1_7_3 <= buffers_0_28_3;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_8_0 <= buffers_0_35_0;
    end else begin
      if (_T_1092) begin
        buffers_1_8_0 <= buffers_0_34_0;
      end else begin
        if (_T_1090) begin
          buffers_1_8_0 <= buffers_0_33_0;
        end else begin
          buffers_1_8_0 <= buffers_0_32_0;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_8_1 <= buffers_0_35_1;
    end else begin
      if (_T_1092) begin
        buffers_1_8_1 <= buffers_0_34_1;
      end else begin
        if (_T_1090) begin
          buffers_1_8_1 <= buffers_0_33_1;
        end else begin
          buffers_1_8_1 <= buffers_0_32_1;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_8_2 <= buffers_0_35_2;
    end else begin
      if (_T_1092) begin
        buffers_1_8_2 <= buffers_0_34_2;
      end else begin
        if (_T_1090) begin
          buffers_1_8_2 <= buffers_0_33_2;
        end else begin
          buffers_1_8_2 <= buffers_0_32_2;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_8_3 <= buffers_0_35_3;
    end else begin
      if (_T_1092) begin
        buffers_1_8_3 <= buffers_0_34_3;
      end else begin
        if (_T_1090) begin
          buffers_1_8_3 <= buffers_0_33_3;
        end else begin
          buffers_1_8_3 <= buffers_0_32_3;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_9_0 <= buffers_0_39_0;
    end else begin
      if (_T_1092) begin
        buffers_1_9_0 <= buffers_0_38_0;
      end else begin
        if (_T_1090) begin
          buffers_1_9_0 <= buffers_0_37_0;
        end else begin
          buffers_1_9_0 <= buffers_0_36_0;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_9_1 <= buffers_0_39_1;
    end else begin
      if (_T_1092) begin
        buffers_1_9_1 <= buffers_0_38_1;
      end else begin
        if (_T_1090) begin
          buffers_1_9_1 <= buffers_0_37_1;
        end else begin
          buffers_1_9_1 <= buffers_0_36_1;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_9_2 <= buffers_0_39_2;
    end else begin
      if (_T_1092) begin
        buffers_1_9_2 <= buffers_0_38_2;
      end else begin
        if (_T_1090) begin
          buffers_1_9_2 <= buffers_0_37_2;
        end else begin
          buffers_1_9_2 <= buffers_0_36_2;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_9_3 <= buffers_0_39_3;
    end else begin
      if (_T_1092) begin
        buffers_1_9_3 <= buffers_0_38_3;
      end else begin
        if (_T_1090) begin
          buffers_1_9_3 <= buffers_0_37_3;
        end else begin
          buffers_1_9_3 <= buffers_0_36_3;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_10_0 <= buffers_0_43_0;
    end else begin
      if (_T_1092) begin
        buffers_1_10_0 <= buffers_0_42_0;
      end else begin
        if (_T_1090) begin
          buffers_1_10_0 <= buffers_0_41_0;
        end else begin
          buffers_1_10_0 <= buffers_0_40_0;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_10_1 <= buffers_0_43_1;
    end else begin
      if (_T_1092) begin
        buffers_1_10_1 <= buffers_0_42_1;
      end else begin
        if (_T_1090) begin
          buffers_1_10_1 <= buffers_0_41_1;
        end else begin
          buffers_1_10_1 <= buffers_0_40_1;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_10_2 <= buffers_0_43_2;
    end else begin
      if (_T_1092) begin
        buffers_1_10_2 <= buffers_0_42_2;
      end else begin
        if (_T_1090) begin
          buffers_1_10_2 <= buffers_0_41_2;
        end else begin
          buffers_1_10_2 <= buffers_0_40_2;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_10_3 <= buffers_0_43_3;
    end else begin
      if (_T_1092) begin
        buffers_1_10_3 <= buffers_0_42_3;
      end else begin
        if (_T_1090) begin
          buffers_1_10_3 <= buffers_0_41_3;
        end else begin
          buffers_1_10_3 <= buffers_0_40_3;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_11_0 <= buffers_0_47_0;
    end else begin
      if (_T_1092) begin
        buffers_1_11_0 <= buffers_0_46_0;
      end else begin
        if (_T_1090) begin
          buffers_1_11_0 <= buffers_0_45_0;
        end else begin
          buffers_1_11_0 <= buffers_0_44_0;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_11_1 <= buffers_0_47_1;
    end else begin
      if (_T_1092) begin
        buffers_1_11_1 <= buffers_0_46_1;
      end else begin
        if (_T_1090) begin
          buffers_1_11_1 <= buffers_0_45_1;
        end else begin
          buffers_1_11_1 <= buffers_0_44_1;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_11_2 <= buffers_0_47_2;
    end else begin
      if (_T_1092) begin
        buffers_1_11_2 <= buffers_0_46_2;
      end else begin
        if (_T_1090) begin
          buffers_1_11_2 <= buffers_0_45_2;
        end else begin
          buffers_1_11_2 <= buffers_0_44_2;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_11_3 <= buffers_0_47_3;
    end else begin
      if (_T_1092) begin
        buffers_1_11_3 <= buffers_0_46_3;
      end else begin
        if (_T_1090) begin
          buffers_1_11_3 <= buffers_0_45_3;
        end else begin
          buffers_1_11_3 <= buffers_0_44_3;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_12_0 <= buffers_0_51_0;
    end else begin
      if (_T_1092) begin
        buffers_1_12_0 <= buffers_0_50_0;
      end else begin
        if (_T_1090) begin
          buffers_1_12_0 <= buffers_0_49_0;
        end else begin
          buffers_1_12_0 <= buffers_0_48_0;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_12_1 <= buffers_0_51_1;
    end else begin
      if (_T_1092) begin
        buffers_1_12_1 <= buffers_0_50_1;
      end else begin
        if (_T_1090) begin
          buffers_1_12_1 <= buffers_0_49_1;
        end else begin
          buffers_1_12_1 <= buffers_0_48_1;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_12_2 <= buffers_0_51_2;
    end else begin
      if (_T_1092) begin
        buffers_1_12_2 <= buffers_0_50_2;
      end else begin
        if (_T_1090) begin
          buffers_1_12_2 <= buffers_0_49_2;
        end else begin
          buffers_1_12_2 <= buffers_0_48_2;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_12_3 <= buffers_0_51_3;
    end else begin
      if (_T_1092) begin
        buffers_1_12_3 <= buffers_0_50_3;
      end else begin
        if (_T_1090) begin
          buffers_1_12_3 <= buffers_0_49_3;
        end else begin
          buffers_1_12_3 <= buffers_0_48_3;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_13_0 <= buffers_0_55_0;
    end else begin
      if (_T_1092) begin
        buffers_1_13_0 <= buffers_0_54_0;
      end else begin
        if (_T_1090) begin
          buffers_1_13_0 <= buffers_0_53_0;
        end else begin
          buffers_1_13_0 <= buffers_0_52_0;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_13_1 <= buffers_0_55_1;
    end else begin
      if (_T_1092) begin
        buffers_1_13_1 <= buffers_0_54_1;
      end else begin
        if (_T_1090) begin
          buffers_1_13_1 <= buffers_0_53_1;
        end else begin
          buffers_1_13_1 <= buffers_0_52_1;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_13_2 <= buffers_0_55_2;
    end else begin
      if (_T_1092) begin
        buffers_1_13_2 <= buffers_0_54_2;
      end else begin
        if (_T_1090) begin
          buffers_1_13_2 <= buffers_0_53_2;
        end else begin
          buffers_1_13_2 <= buffers_0_52_2;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_13_3 <= buffers_0_55_3;
    end else begin
      if (_T_1092) begin
        buffers_1_13_3 <= buffers_0_54_3;
      end else begin
        if (_T_1090) begin
          buffers_1_13_3 <= buffers_0_53_3;
        end else begin
          buffers_1_13_3 <= buffers_0_52_3;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_14_0 <= buffers_0_59_0;
    end else begin
      if (_T_1092) begin
        buffers_1_14_0 <= buffers_0_58_0;
      end else begin
        if (_T_1090) begin
          buffers_1_14_0 <= buffers_0_57_0;
        end else begin
          buffers_1_14_0 <= buffers_0_56_0;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_14_1 <= buffers_0_59_1;
    end else begin
      if (_T_1092) begin
        buffers_1_14_1 <= buffers_0_58_1;
      end else begin
        if (_T_1090) begin
          buffers_1_14_1 <= buffers_0_57_1;
        end else begin
          buffers_1_14_1 <= buffers_0_56_1;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_14_2 <= buffers_0_59_2;
    end else begin
      if (_T_1092) begin
        buffers_1_14_2 <= buffers_0_58_2;
      end else begin
        if (_T_1090) begin
          buffers_1_14_2 <= buffers_0_57_2;
        end else begin
          buffers_1_14_2 <= buffers_0_56_2;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_14_3 <= buffers_0_59_3;
    end else begin
      if (_T_1092) begin
        buffers_1_14_3 <= buffers_0_58_3;
      end else begin
        if (_T_1090) begin
          buffers_1_14_3 <= buffers_0_57_3;
        end else begin
          buffers_1_14_3 <= buffers_0_56_3;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_15_0 <= buffers_0_63_0;
    end else begin
      if (_T_1092) begin
        buffers_1_15_0 <= buffers_0_62_0;
      end else begin
        if (_T_1090) begin
          buffers_1_15_0 <= buffers_0_61_0;
        end else begin
          buffers_1_15_0 <= buffers_0_60_0;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_15_1 <= buffers_0_63_1;
    end else begin
      if (_T_1092) begin
        buffers_1_15_1 <= buffers_0_62_1;
      end else begin
        if (_T_1090) begin
          buffers_1_15_1 <= buffers_0_61_1;
        end else begin
          buffers_1_15_1 <= buffers_0_60_1;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_15_2 <= buffers_0_63_2;
    end else begin
      if (_T_1092) begin
        buffers_1_15_2 <= buffers_0_62_2;
      end else begin
        if (_T_1090) begin
          buffers_1_15_2 <= buffers_0_61_2;
        end else begin
          buffers_1_15_2 <= buffers_0_60_2;
        end
      end
    end
    if (_T_1094) begin
      buffers_1_15_3 <= buffers_0_63_3;
    end else begin
      if (_T_1092) begin
        buffers_1_15_3 <= buffers_0_62_3;
      end else begin
        if (_T_1090) begin
          buffers_1_15_3 <= buffers_0_61_3;
        end else begin
          buffers_1_15_3 <= buffers_0_60_3;
        end
      end
    end
    if (_T_1782) begin
      buffers_2_0_0 <= buffers_1_3_0;
    end else begin
      if (_T_1780) begin
        buffers_2_0_0 <= buffers_1_2_0;
      end else begin
        if (_T_1778) begin
          buffers_2_0_0 <= buffers_1_1_0;
        end else begin
          buffers_2_0_0 <= buffers_1_0_0;
        end
      end
    end
    if (_T_1782) begin
      buffers_2_0_1 <= buffers_1_3_1;
    end else begin
      if (_T_1780) begin
        buffers_2_0_1 <= buffers_1_2_1;
      end else begin
        if (_T_1778) begin
          buffers_2_0_1 <= buffers_1_1_1;
        end else begin
          buffers_2_0_1 <= buffers_1_0_1;
        end
      end
    end
    if (_T_1782) begin
      buffers_2_0_2 <= buffers_1_3_2;
    end else begin
      if (_T_1780) begin
        buffers_2_0_2 <= buffers_1_2_2;
      end else begin
        if (_T_1778) begin
          buffers_2_0_2 <= buffers_1_1_2;
        end else begin
          buffers_2_0_2 <= buffers_1_0_2;
        end
      end
    end
    if (_T_1782) begin
      buffers_2_0_3 <= buffers_1_3_3;
    end else begin
      if (_T_1780) begin
        buffers_2_0_3 <= buffers_1_2_3;
      end else begin
        if (_T_1778) begin
          buffers_2_0_3 <= buffers_1_1_3;
        end else begin
          buffers_2_0_3 <= buffers_1_0_3;
        end
      end
    end
    if (_T_1782) begin
      buffers_2_1_0 <= buffers_1_7_0;
    end else begin
      if (_T_1780) begin
        buffers_2_1_0 <= buffers_1_6_0;
      end else begin
        if (_T_1778) begin
          buffers_2_1_0 <= buffers_1_5_0;
        end else begin
          buffers_2_1_0 <= buffers_1_4_0;
        end
      end
    end
    if (_T_1782) begin
      buffers_2_1_1 <= buffers_1_7_1;
    end else begin
      if (_T_1780) begin
        buffers_2_1_1 <= buffers_1_6_1;
      end else begin
        if (_T_1778) begin
          buffers_2_1_1 <= buffers_1_5_1;
        end else begin
          buffers_2_1_1 <= buffers_1_4_1;
        end
      end
    end
    if (_T_1782) begin
      buffers_2_1_2 <= buffers_1_7_2;
    end else begin
      if (_T_1780) begin
        buffers_2_1_2 <= buffers_1_6_2;
      end else begin
        if (_T_1778) begin
          buffers_2_1_2 <= buffers_1_5_2;
        end else begin
          buffers_2_1_2 <= buffers_1_4_2;
        end
      end
    end
    if (_T_1782) begin
      buffers_2_1_3 <= buffers_1_7_3;
    end else begin
      if (_T_1780) begin
        buffers_2_1_3 <= buffers_1_6_3;
      end else begin
        if (_T_1778) begin
          buffers_2_1_3 <= buffers_1_5_3;
        end else begin
          buffers_2_1_3 <= buffers_1_4_3;
        end
      end
    end
    if (_T_1782) begin
      buffers_2_2_0 <= buffers_1_11_0;
    end else begin
      if (_T_1780) begin
        buffers_2_2_0 <= buffers_1_10_0;
      end else begin
        if (_T_1778) begin
          buffers_2_2_0 <= buffers_1_9_0;
        end else begin
          buffers_2_2_0 <= buffers_1_8_0;
        end
      end
    end
    if (_T_1782) begin
      buffers_2_2_1 <= buffers_1_11_1;
    end else begin
      if (_T_1780) begin
        buffers_2_2_1 <= buffers_1_10_1;
      end else begin
        if (_T_1778) begin
          buffers_2_2_1 <= buffers_1_9_1;
        end else begin
          buffers_2_2_1 <= buffers_1_8_1;
        end
      end
    end
    if (_T_1782) begin
      buffers_2_2_2 <= buffers_1_11_2;
    end else begin
      if (_T_1780) begin
        buffers_2_2_2 <= buffers_1_10_2;
      end else begin
        if (_T_1778) begin
          buffers_2_2_2 <= buffers_1_9_2;
        end else begin
          buffers_2_2_2 <= buffers_1_8_2;
        end
      end
    end
    if (_T_1782) begin
      buffers_2_2_3 <= buffers_1_11_3;
    end else begin
      if (_T_1780) begin
        buffers_2_2_3 <= buffers_1_10_3;
      end else begin
        if (_T_1778) begin
          buffers_2_2_3 <= buffers_1_9_3;
        end else begin
          buffers_2_2_3 <= buffers_1_8_3;
        end
      end
    end
    if (_T_1782) begin
      buffers_2_3_0 <= buffers_1_15_0;
    end else begin
      if (_T_1780) begin
        buffers_2_3_0 <= buffers_1_14_0;
      end else begin
        if (_T_1778) begin
          buffers_2_3_0 <= buffers_1_13_0;
        end else begin
          buffers_2_3_0 <= buffers_1_12_0;
        end
      end
    end
    if (_T_1782) begin
      buffers_2_3_1 <= buffers_1_15_1;
    end else begin
      if (_T_1780) begin
        buffers_2_3_1 <= buffers_1_14_1;
      end else begin
        if (_T_1778) begin
          buffers_2_3_1 <= buffers_1_13_1;
        end else begin
          buffers_2_3_1 <= buffers_1_12_1;
        end
      end
    end
    if (_T_1782) begin
      buffers_2_3_2 <= buffers_1_15_2;
    end else begin
      if (_T_1780) begin
        buffers_2_3_2 <= buffers_1_14_2;
      end else begin
        if (_T_1778) begin
          buffers_2_3_2 <= buffers_1_13_2;
        end else begin
          buffers_2_3_2 <= buffers_1_12_2;
        end
      end
    end
    if (_T_1782) begin
      buffers_2_3_3 <= buffers_1_15_3;
    end else begin
      if (_T_1780) begin
        buffers_2_3_3 <= buffers_1_14_3;
      end else begin
        if (_T_1778) begin
          buffers_2_3_3 <= buffers_1_13_3;
        end else begin
          buffers_2_3_3 <= buffers_1_12_3;
        end
      end
    end
    if (_T_1954) begin
      buffers_3_0_0 <= buffers_2_3_0;
    end else begin
      if (_T_1952) begin
        buffers_3_0_0 <= buffers_2_2_0;
      end else begin
        if (_T_1950) begin
          buffers_3_0_0 <= buffers_2_1_0;
        end else begin
          buffers_3_0_0 <= buffers_2_0_0;
        end
      end
    end
    if (_T_1954) begin
      buffers_3_0_1 <= buffers_2_3_1;
    end else begin
      if (_T_1952) begin
        buffers_3_0_1 <= buffers_2_2_1;
      end else begin
        if (_T_1950) begin
          buffers_3_0_1 <= buffers_2_1_1;
        end else begin
          buffers_3_0_1 <= buffers_2_0_1;
        end
      end
    end
    if (_T_1954) begin
      buffers_3_0_2 <= buffers_2_3_2;
    end else begin
      if (_T_1952) begin
        buffers_3_0_2 <= buffers_2_2_2;
      end else begin
        if (_T_1950) begin
          buffers_3_0_2 <= buffers_2_1_2;
        end else begin
          buffers_3_0_2 <= buffers_2_0_2;
        end
      end
    end
    if (_T_1954) begin
      buffers_3_0_3 <= buffers_2_3_3;
    end else begin
      if (_T_1952) begin
        buffers_3_0_3 <= buffers_2_2_3;
      end else begin
        if (_T_1950) begin
          buffers_3_0_3 <= buffers_2_1_3;
        end else begin
          buffers_3_0_3 <= buffers_2_0_3;
        end
      end
    end
    if (reset) begin
      _T_1988 <= 1'h0;
    end else begin
      _T_1988 <= _T_1052;
    end
    if (reset) begin
      _T_1990 <= 1'h0;
    end else begin
      _T_1990 <= _T_1988;
    end
    if (reset) begin
      vld <= 1'h0;
    end else begin
      vld <= _T_1990;
    end
    if (reset) begin
      lastVld <= 1'h0;
    end else begin
      lastVld <= vld;
    end
  end
endmodule
module FanoutAWS(
  input         clock,
  input  [15:0] io_in,
  output [15:0] io_out_0,
  output [15:0] io_out_1,
  output [15:0] io_out_2,
  output [15:0] io_out_3,
  output [15:0] io_out_4,
  output [15:0] io_out_5,
  output [15:0] io_out_6,
  output [15:0] io_out_7,
  output [15:0] io_out_8,
  output [15:0] io_out_9,
  output [15:0] io_out_10,
  output [15:0] io_out_11,
  output [15:0] io_out_12,
  output [15:0] io_out_13,
  output [15:0] io_out_14,
  output [15:0] io_out_15,
  output [15:0] io_out_16,
  output [15:0] io_out_17,
  output [15:0] io_out_18,
  output [15:0] io_out_19,
  output [15:0] io_out_20,
  output [15:0] io_out_21,
  output [15:0] io_out_22,
  output [15:0] io_out_23,
  output [15:0] io_out_24,
  output [15:0] io_out_25,
  output [15:0] io_out_26,
  output [15:0] io_out_27,
  output [15:0] io_out_28,
  output [15:0] io_out_29,
  output [15:0] io_out_30,
  output [15:0] io_out_31,
  output [15:0] io_out_32,
  output [15:0] io_out_33,
  output [15:0] io_out_34,
  output [15:0] io_out_35,
  output [15:0] io_out_36,
  output [15:0] io_out_37,
  output [15:0] io_out_38,
  output [15:0] io_out_39,
  output [15:0] io_out_40,
  output [15:0] io_out_41,
  output [15:0] io_out_42,
  output [15:0] io_out_43,
  output [15:0] io_out_44,
  output [15:0] io_out_45,
  output [15:0] io_out_46,
  output [15:0] io_out_47,
  output [15:0] io_out_48,
  output [15:0] io_out_49,
  output [15:0] io_out_50,
  output [15:0] io_out_51,
  output [15:0] io_out_52,
  output [15:0] io_out_53,
  output [15:0] io_out_54,
  output [15:0] io_out_55,
  output [15:0] io_out_56,
  output [15:0] io_out_57,
  output [15:0] io_out_58,
  output [15:0] io_out_59,
  output [15:0] io_out_60,
  output [15:0] io_out_61,
  output [15:0] io_out_62,
  output [15:0] io_out_63,
  output [15:0] io_out_64,
  output [15:0] io_out_65,
  output [15:0] io_out_66,
  output [15:0] io_out_67,
  output [15:0] io_out_68,
  output [15:0] io_out_69,
  output [15:0] io_out_70,
  output [15:0] io_out_71,
  output [15:0] io_out_72,
  output [15:0] io_out_73,
  output [15:0] io_out_74,
  output [15:0] io_out_75,
  output [15:0] io_out_76,
  output [15:0] io_out_77,
  output [15:0] io_out_78,
  output [15:0] io_out_79,
  output [15:0] io_out_80,
  output [15:0] io_out_81,
  output [15:0] io_out_82,
  output [15:0] io_out_83,
  output [15:0] io_out_84,
  output [15:0] io_out_85,
  output [15:0] io_out_86,
  output [15:0] io_out_87,
  output [15:0] io_out_88,
  output [15:0] io_out_89,
  output [15:0] io_out_90,
  output [15:0] io_out_91,
  output [15:0] io_out_92,
  output [15:0] io_out_93,
  output [15:0] io_out_94,
  output [15:0] io_out_95,
  output [15:0] io_out_96,
  output [15:0] io_out_97,
  output [15:0] io_out_98,
  output [15:0] io_out_99,
  output [15:0] io_out_100,
  output [15:0] io_out_101,
  output [15:0] io_out_102,
  output [15:0] io_out_103,
  output [15:0] io_out_104,
  output [15:0] io_out_105,
  output [15:0] io_out_106,
  output [15:0] io_out_107,
  output [15:0] io_out_108,
  output [15:0] io_out_109,
  output [15:0] io_out_110,
  output [15:0] io_out_111,
  output [15:0] io_out_112,
  output [15:0] io_out_113,
  output [15:0] io_out_114,
  output [15:0] io_out_115,
  output [15:0] io_out_116,
  output [15:0] io_out_117,
  output [15:0] io_out_118,
  output [15:0] io_out_119,
  output [15:0] io_out_120,
  output [15:0] io_out_121,
  output [15:0] io_out_122,
  output [15:0] io_out_123,
  output [15:0] io_out_124,
  output [15:0] io_out_125,
  output [15:0] io_out_126,
  output [15:0] io_out_127
);
  reg [15:0] dataVecs_1_0; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_0;
  reg [15:0] dataVecs_1_1; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_1;
  reg [15:0] dataVecs_1_2; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_2;
  reg [15:0] dataVecs_1_3; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_3;
  reg [15:0] dataVecs_1_4; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_4;
  reg [15:0] dataVecs_2_0; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_5;
  reg [15:0] dataVecs_2_1; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_6;
  reg [15:0] dataVecs_2_2; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_7;
  reg [15:0] dataVecs_2_3; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_8;
  reg [15:0] dataVecs_2_4; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_9;
  reg [15:0] dataVecs_2_5; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_10;
  reg [15:0] dataVecs_2_6; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_11;
  reg [15:0] dataVecs_2_7; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_12;
  reg [15:0] dataVecs_2_8; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_13;
  reg [15:0] dataVecs_2_9; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_14;
  reg [15:0] dataVecs_2_10; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_15;
  reg [15:0] dataVecs_2_11; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_16;
  reg [15:0] dataVecs_2_12; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_17;
  reg [15:0] dataVecs_2_13; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_18;
  reg [15:0] dataVecs_2_14; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_19;
  reg [15:0] dataVecs_2_15; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_20;
  reg [15:0] dataVecs_2_16; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_21;
  reg [15:0] dataVecs_2_17; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_22;
  reg [15:0] dataVecs_2_18; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_23;
  reg [15:0] dataVecs_2_19; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_24;
  reg [15:0] dataVecs_2_20; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_25;
  reg [15:0] dataVecs_2_21; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_26;
  reg [15:0] dataVecs_2_22; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_27;
  reg [15:0] dataVecs_2_23; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_28;
  reg [15:0] dataVecs_2_24; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_29;
  reg [15:0] dataVecs_3_0; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_30;
  reg [15:0] dataVecs_3_1; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_31;
  reg [15:0] dataVecs_3_2; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_32;
  reg [15:0] dataVecs_3_3; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_33;
  reg [15:0] dataVecs_3_4; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_34;
  reg [15:0] dataVecs_3_5; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_35;
  reg [15:0] dataVecs_3_6; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_36;
  reg [15:0] dataVecs_3_7; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_37;
  reg [15:0] dataVecs_3_8; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_38;
  reg [15:0] dataVecs_3_9; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_39;
  reg [15:0] dataVecs_3_10; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_40;
  reg [15:0] dataVecs_3_11; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_41;
  reg [15:0] dataVecs_3_12; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_42;
  reg [15:0] dataVecs_3_13; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_43;
  reg [15:0] dataVecs_3_14; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_44;
  reg [15:0] dataVecs_3_15; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_45;
  reg [15:0] dataVecs_3_16; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_46;
  reg [15:0] dataVecs_3_17; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_47;
  reg [15:0] dataVecs_3_18; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_48;
  reg [15:0] dataVecs_3_19; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_49;
  reg [15:0] dataVecs_3_20; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_50;
  reg [15:0] dataVecs_3_21; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_51;
  reg [15:0] dataVecs_3_22; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_52;
  reg [15:0] dataVecs_3_23; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_53;
  reg [15:0] dataVecs_3_24; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_54;
  reg [15:0] dataVecs_3_25; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_55;
  reg [15:0] dataVecs_3_26; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_56;
  reg [15:0] dataVecs_3_27; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_57;
  reg [15:0] dataVecs_3_28; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_58;
  reg [15:0] dataVecs_3_29; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_59;
  reg [15:0] dataVecs_3_30; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_60;
  reg [15:0] dataVecs_3_31; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_61;
  reg [15:0] dataVecs_3_32; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_62;
  reg [15:0] dataVecs_3_33; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_63;
  reg [15:0] dataVecs_3_34; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_64;
  reg [15:0] dataVecs_3_35; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_65;
  reg [15:0] dataVecs_3_36; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_66;
  reg [15:0] dataVecs_3_37; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_67;
  reg [15:0] dataVecs_3_38; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_68;
  reg [15:0] dataVecs_3_39; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_69;
  reg [15:0] dataVecs_3_40; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_70;
  reg [15:0] dataVecs_3_41; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_71;
  reg [15:0] dataVecs_3_42; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_72;
  reg [15:0] dataVecs_3_43; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_73;
  reg [15:0] dataVecs_3_44; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_74;
  reg [15:0] dataVecs_3_45; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_75;
  reg [15:0] dataVecs_3_46; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_76;
  reg [15:0] dataVecs_3_47; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_77;
  reg [15:0] dataVecs_3_48; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_78;
  reg [15:0] dataVecs_3_49; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_79;
  reg [15:0] dataVecs_3_50; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_80;
  reg [15:0] dataVecs_3_51; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_81;
  reg [15:0] dataVecs_3_52; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_82;
  reg [15:0] dataVecs_3_53; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_83;
  reg [15:0] dataVecs_3_54; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_84;
  reg [15:0] dataVecs_3_55; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_85;
  reg [15:0] dataVecs_3_56; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_86;
  reg [15:0] dataVecs_3_57; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_87;
  reg [15:0] dataVecs_3_58; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_88;
  reg [15:0] dataVecs_3_59; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_89;
  reg [15:0] dataVecs_3_60; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_90;
  reg [15:0] dataVecs_3_61; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_91;
  reg [15:0] dataVecs_3_62; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_92;
  reg [15:0] dataVecs_3_63; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_93;
  reg [15:0] dataVecs_3_64; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_94;
  reg [15:0] dataVecs_3_65; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_95;
  reg [15:0] dataVecs_3_66; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_96;
  reg [15:0] dataVecs_3_67; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_97;
  reg [15:0] dataVecs_3_68; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_98;
  reg [15:0] dataVecs_3_69; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_99;
  reg [15:0] dataVecs_3_70; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_100;
  reg [15:0] dataVecs_3_71; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_101;
  reg [15:0] dataVecs_3_72; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_102;
  reg [15:0] dataVecs_3_73; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_103;
  reg [15:0] dataVecs_3_74; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_104;
  reg [15:0] dataVecs_3_75; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_105;
  reg [15:0] dataVecs_3_76; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_106;
  reg [15:0] dataVecs_3_77; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_107;
  reg [15:0] dataVecs_3_78; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_108;
  reg [15:0] dataVecs_3_79; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_109;
  reg [15:0] dataVecs_3_80; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_110;
  reg [15:0] dataVecs_3_81; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_111;
  reg [15:0] dataVecs_3_82; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_112;
  reg [15:0] dataVecs_3_83; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_113;
  reg [15:0] dataVecs_3_84; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_114;
  reg [15:0] dataVecs_3_85; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_115;
  reg [15:0] dataVecs_3_86; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_116;
  reg [15:0] dataVecs_3_87; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_117;
  reg [15:0] dataVecs_3_88; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_118;
  reg [15:0] dataVecs_3_89; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_119;
  reg [15:0] dataVecs_3_90; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_120;
  reg [15:0] dataVecs_3_91; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_121;
  reg [15:0] dataVecs_3_92; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_122;
  reg [15:0] dataVecs_3_93; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_123;
  reg [15:0] dataVecs_3_94; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_124;
  reg [15:0] dataVecs_3_95; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_125;
  reg [15:0] dataVecs_3_96; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_126;
  reg [15:0] dataVecs_3_97; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_127;
  reg [15:0] dataVecs_3_98; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_128;
  reg [15:0] dataVecs_3_99; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_129;
  reg [15:0] dataVecs_3_100; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_130;
  reg [15:0] dataVecs_3_101; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_131;
  reg [15:0] dataVecs_3_102; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_132;
  reg [15:0] dataVecs_3_103; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_133;
  reg [15:0] dataVecs_3_104; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_134;
  reg [15:0] dataVecs_3_105; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_135;
  reg [15:0] dataVecs_3_106; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_136;
  reg [15:0] dataVecs_3_107; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_137;
  reg [15:0] dataVecs_3_108; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_138;
  reg [15:0] dataVecs_3_109; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_139;
  reg [15:0] dataVecs_3_110; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_140;
  reg [15:0] dataVecs_3_111; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_141;
  reg [15:0] dataVecs_3_112; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_142;
  reg [15:0] dataVecs_3_113; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_143;
  reg [15:0] dataVecs_3_114; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_144;
  reg [15:0] dataVecs_3_115; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_145;
  reg [15:0] dataVecs_3_116; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_146;
  reg [15:0] dataVecs_3_117; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_147;
  reg [15:0] dataVecs_3_118; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_148;
  reg [15:0] dataVecs_3_119; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_149;
  reg [15:0] dataVecs_3_120; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_150;
  reg [15:0] dataVecs_3_121; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_151;
  reg [15:0] dataVecs_3_122; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_152;
  reg [15:0] dataVecs_3_123; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_153;
  reg [15:0] dataVecs_3_124; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_154;
  reg [15:0] dataVecs_3_125; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_155;
  reg [15:0] dataVecs_3_126; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_156;
  reg [15:0] dataVecs_3_127; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_157;
  assign io_out_0 = dataVecs_3_0;
  assign io_out_1 = dataVecs_3_1;
  assign io_out_2 = dataVecs_3_2;
  assign io_out_3 = dataVecs_3_3;
  assign io_out_4 = dataVecs_3_4;
  assign io_out_5 = dataVecs_3_5;
  assign io_out_6 = dataVecs_3_6;
  assign io_out_7 = dataVecs_3_7;
  assign io_out_8 = dataVecs_3_8;
  assign io_out_9 = dataVecs_3_9;
  assign io_out_10 = dataVecs_3_10;
  assign io_out_11 = dataVecs_3_11;
  assign io_out_12 = dataVecs_3_12;
  assign io_out_13 = dataVecs_3_13;
  assign io_out_14 = dataVecs_3_14;
  assign io_out_15 = dataVecs_3_15;
  assign io_out_16 = dataVecs_3_16;
  assign io_out_17 = dataVecs_3_17;
  assign io_out_18 = dataVecs_3_18;
  assign io_out_19 = dataVecs_3_19;
  assign io_out_20 = dataVecs_3_20;
  assign io_out_21 = dataVecs_3_21;
  assign io_out_22 = dataVecs_3_22;
  assign io_out_23 = dataVecs_3_23;
  assign io_out_24 = dataVecs_3_24;
  assign io_out_25 = dataVecs_3_25;
  assign io_out_26 = dataVecs_3_26;
  assign io_out_27 = dataVecs_3_27;
  assign io_out_28 = dataVecs_3_28;
  assign io_out_29 = dataVecs_3_29;
  assign io_out_30 = dataVecs_3_30;
  assign io_out_31 = dataVecs_3_31;
  assign io_out_32 = dataVecs_3_32;
  assign io_out_33 = dataVecs_3_33;
  assign io_out_34 = dataVecs_3_34;
  assign io_out_35 = dataVecs_3_35;
  assign io_out_36 = dataVecs_3_36;
  assign io_out_37 = dataVecs_3_37;
  assign io_out_38 = dataVecs_3_38;
  assign io_out_39 = dataVecs_3_39;
  assign io_out_40 = dataVecs_3_40;
  assign io_out_41 = dataVecs_3_41;
  assign io_out_42 = dataVecs_3_42;
  assign io_out_43 = dataVecs_3_43;
  assign io_out_44 = dataVecs_3_44;
  assign io_out_45 = dataVecs_3_45;
  assign io_out_46 = dataVecs_3_46;
  assign io_out_47 = dataVecs_3_47;
  assign io_out_48 = dataVecs_3_48;
  assign io_out_49 = dataVecs_3_49;
  assign io_out_50 = dataVecs_3_50;
  assign io_out_51 = dataVecs_3_51;
  assign io_out_52 = dataVecs_3_52;
  assign io_out_53 = dataVecs_3_53;
  assign io_out_54 = dataVecs_3_54;
  assign io_out_55 = dataVecs_3_55;
  assign io_out_56 = dataVecs_3_56;
  assign io_out_57 = dataVecs_3_57;
  assign io_out_58 = dataVecs_3_58;
  assign io_out_59 = dataVecs_3_59;
  assign io_out_60 = dataVecs_3_60;
  assign io_out_61 = dataVecs_3_61;
  assign io_out_62 = dataVecs_3_62;
  assign io_out_63 = dataVecs_3_63;
  assign io_out_64 = dataVecs_3_64;
  assign io_out_65 = dataVecs_3_65;
  assign io_out_66 = dataVecs_3_66;
  assign io_out_67 = dataVecs_3_67;
  assign io_out_68 = dataVecs_3_68;
  assign io_out_69 = dataVecs_3_69;
  assign io_out_70 = dataVecs_3_70;
  assign io_out_71 = dataVecs_3_71;
  assign io_out_72 = dataVecs_3_72;
  assign io_out_73 = dataVecs_3_73;
  assign io_out_74 = dataVecs_3_74;
  assign io_out_75 = dataVecs_3_75;
  assign io_out_76 = dataVecs_3_76;
  assign io_out_77 = dataVecs_3_77;
  assign io_out_78 = dataVecs_3_78;
  assign io_out_79 = dataVecs_3_79;
  assign io_out_80 = dataVecs_3_80;
  assign io_out_81 = dataVecs_3_81;
  assign io_out_82 = dataVecs_3_82;
  assign io_out_83 = dataVecs_3_83;
  assign io_out_84 = dataVecs_3_84;
  assign io_out_85 = dataVecs_3_85;
  assign io_out_86 = dataVecs_3_86;
  assign io_out_87 = dataVecs_3_87;
  assign io_out_88 = dataVecs_3_88;
  assign io_out_89 = dataVecs_3_89;
  assign io_out_90 = dataVecs_3_90;
  assign io_out_91 = dataVecs_3_91;
  assign io_out_92 = dataVecs_3_92;
  assign io_out_93 = dataVecs_3_93;
  assign io_out_94 = dataVecs_3_94;
  assign io_out_95 = dataVecs_3_95;
  assign io_out_96 = dataVecs_3_96;
  assign io_out_97 = dataVecs_3_97;
  assign io_out_98 = dataVecs_3_98;
  assign io_out_99 = dataVecs_3_99;
  assign io_out_100 = dataVecs_3_100;
  assign io_out_101 = dataVecs_3_101;
  assign io_out_102 = dataVecs_3_102;
  assign io_out_103 = dataVecs_3_103;
  assign io_out_104 = dataVecs_3_104;
  assign io_out_105 = dataVecs_3_105;
  assign io_out_106 = dataVecs_3_106;
  assign io_out_107 = dataVecs_3_107;
  assign io_out_108 = dataVecs_3_108;
  assign io_out_109 = dataVecs_3_109;
  assign io_out_110 = dataVecs_3_110;
  assign io_out_111 = dataVecs_3_111;
  assign io_out_112 = dataVecs_3_112;
  assign io_out_113 = dataVecs_3_113;
  assign io_out_114 = dataVecs_3_114;
  assign io_out_115 = dataVecs_3_115;
  assign io_out_116 = dataVecs_3_116;
  assign io_out_117 = dataVecs_3_117;
  assign io_out_118 = dataVecs_3_118;
  assign io_out_119 = dataVecs_3_119;
  assign io_out_120 = dataVecs_3_120;
  assign io_out_121 = dataVecs_3_121;
  assign io_out_122 = dataVecs_3_122;
  assign io_out_123 = dataVecs_3_123;
  assign io_out_124 = dataVecs_3_124;
  assign io_out_125 = dataVecs_3_125;
  assign io_out_126 = dataVecs_3_126;
  assign io_out_127 = dataVecs_3_127;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  dataVecs_1_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  dataVecs_1_1 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  dataVecs_1_2 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  dataVecs_1_3 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  dataVecs_1_4 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  dataVecs_2_0 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  dataVecs_2_1 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  dataVecs_2_2 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  dataVecs_2_3 = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  dataVecs_2_4 = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  dataVecs_2_5 = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  dataVecs_2_6 = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  dataVecs_2_7 = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  dataVecs_2_8 = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  dataVecs_2_9 = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  dataVecs_2_10 = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  dataVecs_2_11 = _RAND_16[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  dataVecs_2_12 = _RAND_17[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  dataVecs_2_13 = _RAND_18[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  dataVecs_2_14 = _RAND_19[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  dataVecs_2_15 = _RAND_20[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  dataVecs_2_16 = _RAND_21[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  dataVecs_2_17 = _RAND_22[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  dataVecs_2_18 = _RAND_23[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  dataVecs_2_19 = _RAND_24[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  dataVecs_2_20 = _RAND_25[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  dataVecs_2_21 = _RAND_26[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  dataVecs_2_22 = _RAND_27[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  dataVecs_2_23 = _RAND_28[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  dataVecs_2_24 = _RAND_29[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  dataVecs_3_0 = _RAND_30[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  dataVecs_3_1 = _RAND_31[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  dataVecs_3_2 = _RAND_32[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{$random}};
  dataVecs_3_3 = _RAND_33[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{$random}};
  dataVecs_3_4 = _RAND_34[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{$random}};
  dataVecs_3_5 = _RAND_35[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{$random}};
  dataVecs_3_6 = _RAND_36[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{$random}};
  dataVecs_3_7 = _RAND_37[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{$random}};
  dataVecs_3_8 = _RAND_38[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{$random}};
  dataVecs_3_9 = _RAND_39[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{$random}};
  dataVecs_3_10 = _RAND_40[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{$random}};
  dataVecs_3_11 = _RAND_41[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{$random}};
  dataVecs_3_12 = _RAND_42[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{$random}};
  dataVecs_3_13 = _RAND_43[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{$random}};
  dataVecs_3_14 = _RAND_44[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{$random}};
  dataVecs_3_15 = _RAND_45[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{$random}};
  dataVecs_3_16 = _RAND_46[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{$random}};
  dataVecs_3_17 = _RAND_47[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{$random}};
  dataVecs_3_18 = _RAND_48[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{$random}};
  dataVecs_3_19 = _RAND_49[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{$random}};
  dataVecs_3_20 = _RAND_50[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{$random}};
  dataVecs_3_21 = _RAND_51[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{$random}};
  dataVecs_3_22 = _RAND_52[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{$random}};
  dataVecs_3_23 = _RAND_53[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{$random}};
  dataVecs_3_24 = _RAND_54[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{$random}};
  dataVecs_3_25 = _RAND_55[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{$random}};
  dataVecs_3_26 = _RAND_56[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{$random}};
  dataVecs_3_27 = _RAND_57[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{$random}};
  dataVecs_3_28 = _RAND_58[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{$random}};
  dataVecs_3_29 = _RAND_59[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{$random}};
  dataVecs_3_30 = _RAND_60[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{$random}};
  dataVecs_3_31 = _RAND_61[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{$random}};
  dataVecs_3_32 = _RAND_62[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{$random}};
  dataVecs_3_33 = _RAND_63[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{$random}};
  dataVecs_3_34 = _RAND_64[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{$random}};
  dataVecs_3_35 = _RAND_65[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{$random}};
  dataVecs_3_36 = _RAND_66[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{$random}};
  dataVecs_3_37 = _RAND_67[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{$random}};
  dataVecs_3_38 = _RAND_68[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{$random}};
  dataVecs_3_39 = _RAND_69[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{$random}};
  dataVecs_3_40 = _RAND_70[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{$random}};
  dataVecs_3_41 = _RAND_71[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{$random}};
  dataVecs_3_42 = _RAND_72[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{$random}};
  dataVecs_3_43 = _RAND_73[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{$random}};
  dataVecs_3_44 = _RAND_74[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{$random}};
  dataVecs_3_45 = _RAND_75[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{$random}};
  dataVecs_3_46 = _RAND_76[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{$random}};
  dataVecs_3_47 = _RAND_77[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{$random}};
  dataVecs_3_48 = _RAND_78[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{$random}};
  dataVecs_3_49 = _RAND_79[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{$random}};
  dataVecs_3_50 = _RAND_80[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{$random}};
  dataVecs_3_51 = _RAND_81[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{$random}};
  dataVecs_3_52 = _RAND_82[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{$random}};
  dataVecs_3_53 = _RAND_83[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{$random}};
  dataVecs_3_54 = _RAND_84[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{$random}};
  dataVecs_3_55 = _RAND_85[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{$random}};
  dataVecs_3_56 = _RAND_86[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{$random}};
  dataVecs_3_57 = _RAND_87[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{$random}};
  dataVecs_3_58 = _RAND_88[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{$random}};
  dataVecs_3_59 = _RAND_89[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{$random}};
  dataVecs_3_60 = _RAND_90[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{$random}};
  dataVecs_3_61 = _RAND_91[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{$random}};
  dataVecs_3_62 = _RAND_92[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{$random}};
  dataVecs_3_63 = _RAND_93[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{$random}};
  dataVecs_3_64 = _RAND_94[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{$random}};
  dataVecs_3_65 = _RAND_95[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{$random}};
  dataVecs_3_66 = _RAND_96[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{$random}};
  dataVecs_3_67 = _RAND_97[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{$random}};
  dataVecs_3_68 = _RAND_98[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{$random}};
  dataVecs_3_69 = _RAND_99[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{$random}};
  dataVecs_3_70 = _RAND_100[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{$random}};
  dataVecs_3_71 = _RAND_101[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{$random}};
  dataVecs_3_72 = _RAND_102[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{$random}};
  dataVecs_3_73 = _RAND_103[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{$random}};
  dataVecs_3_74 = _RAND_104[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{$random}};
  dataVecs_3_75 = _RAND_105[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{$random}};
  dataVecs_3_76 = _RAND_106[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{$random}};
  dataVecs_3_77 = _RAND_107[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{$random}};
  dataVecs_3_78 = _RAND_108[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{$random}};
  dataVecs_3_79 = _RAND_109[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{$random}};
  dataVecs_3_80 = _RAND_110[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{$random}};
  dataVecs_3_81 = _RAND_111[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{$random}};
  dataVecs_3_82 = _RAND_112[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{$random}};
  dataVecs_3_83 = _RAND_113[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{$random}};
  dataVecs_3_84 = _RAND_114[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{$random}};
  dataVecs_3_85 = _RAND_115[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{$random}};
  dataVecs_3_86 = _RAND_116[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{$random}};
  dataVecs_3_87 = _RAND_117[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{$random}};
  dataVecs_3_88 = _RAND_118[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{$random}};
  dataVecs_3_89 = _RAND_119[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{$random}};
  dataVecs_3_90 = _RAND_120[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{$random}};
  dataVecs_3_91 = _RAND_121[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{$random}};
  dataVecs_3_92 = _RAND_122[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{$random}};
  dataVecs_3_93 = _RAND_123[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{$random}};
  dataVecs_3_94 = _RAND_124[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{$random}};
  dataVecs_3_95 = _RAND_125[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{$random}};
  dataVecs_3_96 = _RAND_126[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{$random}};
  dataVecs_3_97 = _RAND_127[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{$random}};
  dataVecs_3_98 = _RAND_128[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{$random}};
  dataVecs_3_99 = _RAND_129[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{$random}};
  dataVecs_3_100 = _RAND_130[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{$random}};
  dataVecs_3_101 = _RAND_131[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{$random}};
  dataVecs_3_102 = _RAND_132[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{$random}};
  dataVecs_3_103 = _RAND_133[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{$random}};
  dataVecs_3_104 = _RAND_134[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{$random}};
  dataVecs_3_105 = _RAND_135[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{$random}};
  dataVecs_3_106 = _RAND_136[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{$random}};
  dataVecs_3_107 = _RAND_137[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{$random}};
  dataVecs_3_108 = _RAND_138[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{$random}};
  dataVecs_3_109 = _RAND_139[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{$random}};
  dataVecs_3_110 = _RAND_140[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{$random}};
  dataVecs_3_111 = _RAND_141[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{$random}};
  dataVecs_3_112 = _RAND_142[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{$random}};
  dataVecs_3_113 = _RAND_143[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{$random}};
  dataVecs_3_114 = _RAND_144[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{$random}};
  dataVecs_3_115 = _RAND_145[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{$random}};
  dataVecs_3_116 = _RAND_146[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{$random}};
  dataVecs_3_117 = _RAND_147[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{$random}};
  dataVecs_3_118 = _RAND_148[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{$random}};
  dataVecs_3_119 = _RAND_149[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{$random}};
  dataVecs_3_120 = _RAND_150[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{$random}};
  dataVecs_3_121 = _RAND_151[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{$random}};
  dataVecs_3_122 = _RAND_152[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{$random}};
  dataVecs_3_123 = _RAND_153[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{$random}};
  dataVecs_3_124 = _RAND_154[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{$random}};
  dataVecs_3_125 = _RAND_155[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{$random}};
  dataVecs_3_126 = _RAND_156[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{$random}};
  dataVecs_3_127 = _RAND_157[15:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    dataVecs_1_0 <= io_in;
    dataVecs_1_1 <= io_in;
    dataVecs_1_2 <= io_in;
    dataVecs_1_3 <= io_in;
    dataVecs_1_4 <= io_in;
    dataVecs_2_0 <= dataVecs_1_0;
    dataVecs_2_1 <= dataVecs_1_1;
    dataVecs_2_2 <= dataVecs_1_2;
    dataVecs_2_3 <= dataVecs_1_3;
    dataVecs_2_4 <= dataVecs_1_4;
    dataVecs_2_5 <= dataVecs_1_0;
    dataVecs_2_6 <= dataVecs_1_1;
    dataVecs_2_7 <= dataVecs_1_2;
    dataVecs_2_8 <= dataVecs_1_3;
    dataVecs_2_9 <= dataVecs_1_4;
    dataVecs_2_10 <= dataVecs_1_0;
    dataVecs_2_11 <= dataVecs_1_1;
    dataVecs_2_12 <= dataVecs_1_2;
    dataVecs_2_13 <= dataVecs_1_3;
    dataVecs_2_14 <= dataVecs_1_4;
    dataVecs_2_15 <= dataVecs_1_0;
    dataVecs_2_16 <= dataVecs_1_1;
    dataVecs_2_17 <= dataVecs_1_2;
    dataVecs_2_18 <= dataVecs_1_3;
    dataVecs_2_19 <= dataVecs_1_4;
    dataVecs_2_20 <= dataVecs_1_0;
    dataVecs_2_21 <= dataVecs_1_1;
    dataVecs_2_22 <= dataVecs_1_2;
    dataVecs_2_23 <= dataVecs_1_3;
    dataVecs_2_24 <= dataVecs_1_4;
    dataVecs_3_0 <= dataVecs_2_0;
    dataVecs_3_1 <= dataVecs_2_1;
    dataVecs_3_2 <= dataVecs_2_2;
    dataVecs_3_3 <= dataVecs_2_3;
    dataVecs_3_4 <= dataVecs_2_4;
    dataVecs_3_5 <= dataVecs_2_5;
    dataVecs_3_6 <= dataVecs_2_6;
    dataVecs_3_7 <= dataVecs_2_7;
    dataVecs_3_8 <= dataVecs_2_8;
    dataVecs_3_9 <= dataVecs_2_9;
    dataVecs_3_10 <= dataVecs_2_10;
    dataVecs_3_11 <= dataVecs_2_11;
    dataVecs_3_12 <= dataVecs_2_12;
    dataVecs_3_13 <= dataVecs_2_13;
    dataVecs_3_14 <= dataVecs_2_14;
    dataVecs_3_15 <= dataVecs_2_15;
    dataVecs_3_16 <= dataVecs_2_16;
    dataVecs_3_17 <= dataVecs_2_17;
    dataVecs_3_18 <= dataVecs_2_18;
    dataVecs_3_19 <= dataVecs_2_19;
    dataVecs_3_20 <= dataVecs_2_20;
    dataVecs_3_21 <= dataVecs_2_21;
    dataVecs_3_22 <= dataVecs_2_22;
    dataVecs_3_23 <= dataVecs_2_23;
    dataVecs_3_24 <= dataVecs_2_24;
    dataVecs_3_25 <= dataVecs_2_0;
    dataVecs_3_26 <= dataVecs_2_1;
    dataVecs_3_27 <= dataVecs_2_2;
    dataVecs_3_28 <= dataVecs_2_3;
    dataVecs_3_29 <= dataVecs_2_4;
    dataVecs_3_30 <= dataVecs_2_5;
    dataVecs_3_31 <= dataVecs_2_6;
    dataVecs_3_32 <= dataVecs_2_7;
    dataVecs_3_33 <= dataVecs_2_8;
    dataVecs_3_34 <= dataVecs_2_9;
    dataVecs_3_35 <= dataVecs_2_10;
    dataVecs_3_36 <= dataVecs_2_11;
    dataVecs_3_37 <= dataVecs_2_12;
    dataVecs_3_38 <= dataVecs_2_13;
    dataVecs_3_39 <= dataVecs_2_14;
    dataVecs_3_40 <= dataVecs_2_15;
    dataVecs_3_41 <= dataVecs_2_16;
    dataVecs_3_42 <= dataVecs_2_17;
    dataVecs_3_43 <= dataVecs_2_18;
    dataVecs_3_44 <= dataVecs_2_19;
    dataVecs_3_45 <= dataVecs_2_20;
    dataVecs_3_46 <= dataVecs_2_21;
    dataVecs_3_47 <= dataVecs_2_22;
    dataVecs_3_48 <= dataVecs_2_23;
    dataVecs_3_49 <= dataVecs_2_24;
    dataVecs_3_50 <= dataVecs_2_0;
    dataVecs_3_51 <= dataVecs_2_1;
    dataVecs_3_52 <= dataVecs_2_2;
    dataVecs_3_53 <= dataVecs_2_3;
    dataVecs_3_54 <= dataVecs_2_4;
    dataVecs_3_55 <= dataVecs_2_5;
    dataVecs_3_56 <= dataVecs_2_6;
    dataVecs_3_57 <= dataVecs_2_7;
    dataVecs_3_58 <= dataVecs_2_8;
    dataVecs_3_59 <= dataVecs_2_9;
    dataVecs_3_60 <= dataVecs_2_10;
    dataVecs_3_61 <= dataVecs_2_11;
    dataVecs_3_62 <= dataVecs_2_12;
    dataVecs_3_63 <= dataVecs_2_13;
    dataVecs_3_64 <= dataVecs_2_14;
    dataVecs_3_65 <= dataVecs_2_15;
    dataVecs_3_66 <= dataVecs_2_16;
    dataVecs_3_67 <= dataVecs_2_17;
    dataVecs_3_68 <= dataVecs_2_18;
    dataVecs_3_69 <= dataVecs_2_19;
    dataVecs_3_70 <= dataVecs_2_20;
    dataVecs_3_71 <= dataVecs_2_21;
    dataVecs_3_72 <= dataVecs_2_22;
    dataVecs_3_73 <= dataVecs_2_23;
    dataVecs_3_74 <= dataVecs_2_24;
    dataVecs_3_75 <= dataVecs_2_0;
    dataVecs_3_76 <= dataVecs_2_1;
    dataVecs_3_77 <= dataVecs_2_2;
    dataVecs_3_78 <= dataVecs_2_3;
    dataVecs_3_79 <= dataVecs_2_4;
    dataVecs_3_80 <= dataVecs_2_5;
    dataVecs_3_81 <= dataVecs_2_6;
    dataVecs_3_82 <= dataVecs_2_7;
    dataVecs_3_83 <= dataVecs_2_8;
    dataVecs_3_84 <= dataVecs_2_9;
    dataVecs_3_85 <= dataVecs_2_10;
    dataVecs_3_86 <= dataVecs_2_11;
    dataVecs_3_87 <= dataVecs_2_12;
    dataVecs_3_88 <= dataVecs_2_13;
    dataVecs_3_89 <= dataVecs_2_14;
    dataVecs_3_90 <= dataVecs_2_15;
    dataVecs_3_91 <= dataVecs_2_16;
    dataVecs_3_92 <= dataVecs_2_17;
    dataVecs_3_93 <= dataVecs_2_18;
    dataVecs_3_94 <= dataVecs_2_19;
    dataVecs_3_95 <= dataVecs_2_20;
    dataVecs_3_96 <= dataVecs_2_21;
    dataVecs_3_97 <= dataVecs_2_22;
    dataVecs_3_98 <= dataVecs_2_23;
    dataVecs_3_99 <= dataVecs_2_24;
    dataVecs_3_100 <= dataVecs_2_0;
    dataVecs_3_101 <= dataVecs_2_1;
    dataVecs_3_102 <= dataVecs_2_2;
    dataVecs_3_103 <= dataVecs_2_3;
    dataVecs_3_104 <= dataVecs_2_4;
    dataVecs_3_105 <= dataVecs_2_5;
    dataVecs_3_106 <= dataVecs_2_6;
    dataVecs_3_107 <= dataVecs_2_7;
    dataVecs_3_108 <= dataVecs_2_8;
    dataVecs_3_109 <= dataVecs_2_9;
    dataVecs_3_110 <= dataVecs_2_10;
    dataVecs_3_111 <= dataVecs_2_11;
    dataVecs_3_112 <= dataVecs_2_12;
    dataVecs_3_113 <= dataVecs_2_13;
    dataVecs_3_114 <= dataVecs_2_14;
    dataVecs_3_115 <= dataVecs_2_15;
    dataVecs_3_116 <= dataVecs_2_16;
    dataVecs_3_117 <= dataVecs_2_17;
    dataVecs_3_118 <= dataVecs_2_18;
    dataVecs_3_119 <= dataVecs_2_19;
    dataVecs_3_120 <= dataVecs_2_20;
    dataVecs_3_121 <= dataVecs_2_21;
    dataVecs_3_122 <= dataVecs_2_22;
    dataVecs_3_123 <= dataVecs_2_23;
    dataVecs_3_124 <= dataVecs_2_24;
    dataVecs_3_125 <= dataVecs_2_0;
    dataVecs_3_126 <= dataVecs_2_1;
    dataVecs_3_127 <= dataVecs_2_2;
  end
endmodule
module GenericAddSub16(
  input         clock,
  input  [15:0] io_x_i,
  input  [15:0] io_y_i,
  input         io_x_i_neg,
  input         io_x_i_zero,
  input         io_y_i_neg,
  input         io_y_i_zero,
  output [15:0] io_sum_o
);
  reg [15:0] x_i_reg; // @[GenericAddSub16.scala 29:20]
  reg [31:0] _RAND_0;
  reg [15:0] y_i_reg; // @[GenericAddSub16.scala 30:20]
  reg [31:0] _RAND_1;
  reg  x_i_neg_reg; // @[GenericAddSub16.scala 40:28]
  reg [31:0] _RAND_2;
  reg  y_i_neg_reg; // @[GenericAddSub16.scala 41:28]
  reg [31:0] _RAND_3;
  wire  Xilinx_GenericAddSub_16_dss_c_o; // @[GenericAddSub16.scala 56:25]
  wire [15:0] Xilinx_GenericAddSub_16_dss_sum_o; // @[GenericAddSub16.scala 56:25]
  wire  Xilinx_GenericAddSub_16_dss_neg_y_i; // @[GenericAddSub16.scala 56:25]
  wire  Xilinx_GenericAddSub_16_dss_neg_x_i; // @[GenericAddSub16.scala 56:25]
  wire [15:0] Xilinx_GenericAddSub_16_dss_y_i; // @[GenericAddSub16.scala 56:25]
  wire [15:0] Xilinx_GenericAddSub_16_dss_x_i; // @[GenericAddSub16.scala 56:25]
  reg [15:0] _T_16; // @[GenericAddSub16.scala 61:24]
  reg [31:0] _RAND_4;
  wire [15:0] _GEN_0; // @[GenericAddSub16.scala 34:24]
  wire [15:0] _GEN_1; // @[GenericAddSub16.scala 37:24]
  Xilinx_GenericAddSub_16_dss Xilinx_GenericAddSub_16_dss ( // @[GenericAddSub16.scala 56:25]
    .c_o(Xilinx_GenericAddSub_16_dss_c_o),
    .sum_o(Xilinx_GenericAddSub_16_dss_sum_o),
    .neg_y_i(Xilinx_GenericAddSub_16_dss_neg_y_i),
    .neg_x_i(Xilinx_GenericAddSub_16_dss_neg_x_i),
    .y_i(Xilinx_GenericAddSub_16_dss_y_i),
    .x_i(Xilinx_GenericAddSub_16_dss_x_i)
  );
  assign _GEN_0 = io_x_i_zero ? $signed(16'sh0) : $signed(io_x_i); // @[GenericAddSub16.scala 34:24]
  assign _GEN_1 = io_y_i_zero ? $signed(16'sh0) : $signed(io_y_i); // @[GenericAddSub16.scala 37:24]
  assign io_sum_o = _T_16;
  assign Xilinx_GenericAddSub_16_dss_neg_y_i = y_i_neg_reg;
  assign Xilinx_GenericAddSub_16_dss_neg_x_i = x_i_neg_reg;
  assign Xilinx_GenericAddSub_16_dss_y_i = y_i_reg;
  assign Xilinx_GenericAddSub_16_dss_x_i = x_i_reg;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  x_i_reg = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  y_i_reg = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  x_i_neg_reg = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  y_i_neg_reg = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  _T_16 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (io_x_i_zero) begin
      x_i_reg <= 16'sh0;
    end else begin
      x_i_reg <= io_x_i;
    end
    if (io_y_i_zero) begin
      y_i_reg <= 16'sh0;
    end else begin
      y_i_reg <= io_y_i;
    end
    x_i_neg_reg <= io_x_i_neg;
    y_i_neg_reg <= io_y_i_neg;
    _T_16 <= Xilinx_GenericAddSub_16_dss_sum_o;
  end
endmodule
module MultiplyAccumulate(
  input         clock,
  input  [15:0] io_activations_0,
  input  [15:0] io_activations_1,
  input  [15:0] io_activations_2,
  input  [15:0] io_activations_3,
  input  [7:0]  io_weights,
  output [15:0] io_sum
);
  wire  GenericAddSub16_clock; // @[DenseLayer.scala 29:29]
  wire [15:0] GenericAddSub16_io_x_i; // @[DenseLayer.scala 29:29]
  wire [15:0] GenericAddSub16_io_y_i; // @[DenseLayer.scala 29:29]
  wire  GenericAddSub16_io_x_i_neg; // @[DenseLayer.scala 29:29]
  wire  GenericAddSub16_io_x_i_zero; // @[DenseLayer.scala 29:29]
  wire  GenericAddSub16_io_y_i_neg; // @[DenseLayer.scala 29:29]
  wire  GenericAddSub16_io_y_i_zero; // @[DenseLayer.scala 29:29]
  wire [15:0] GenericAddSub16_io_sum_o; // @[DenseLayer.scala 29:29]
  wire  GenericAddSub16_1_clock; // @[DenseLayer.scala 29:29]
  wire [15:0] GenericAddSub16_1_io_x_i; // @[DenseLayer.scala 29:29]
  wire [15:0] GenericAddSub16_1_io_y_i; // @[DenseLayer.scala 29:29]
  wire  GenericAddSub16_1_io_x_i_neg; // @[DenseLayer.scala 29:29]
  wire  GenericAddSub16_1_io_x_i_zero; // @[DenseLayer.scala 29:29]
  wire  GenericAddSub16_1_io_y_i_neg; // @[DenseLayer.scala 29:29]
  wire  GenericAddSub16_1_io_y_i_zero; // @[DenseLayer.scala 29:29]
  wire [15:0] GenericAddSub16_1_io_sum_o; // @[DenseLayer.scala 29:29]
  reg [15:0] numsToSum_0; // @[DenseLayer.scala 68:14]
  reg [31:0] _RAND_0;
  wire  _T_12; // @[DenseLayer.scala 25:35]
  wire  _T_14; // @[DenseLayer.scala 25:24]
  wire  _T_15; // @[DenseLayer.scala 26:33]
  wire  _T_16; // @[DenseLayer.scala 27:35]
  wire  _T_18; // @[DenseLayer.scala 27:24]
  wire  _T_19; // @[DenseLayer.scala 28:33]
  wire  _T_20; // @[DenseLayer.scala 25:35]
  wire  _T_22; // @[DenseLayer.scala 25:24]
  wire  _T_23; // @[DenseLayer.scala 26:33]
  wire  _T_24; // @[DenseLayer.scala 27:35]
  wire  _T_26; // @[DenseLayer.scala 27:24]
  wire  _T_27; // @[DenseLayer.scala 28:33]
  wire [16:0] _T_28; // @[DenseLayer.scala 67:33]
  wire [15:0] _T_29; // @[DenseLayer.scala 67:33]
  wire [15:0] _T_30; // @[DenseLayer.scala 67:33]
  GenericAddSub16 GenericAddSub16 ( // @[DenseLayer.scala 29:29]
    .clock(GenericAddSub16_clock),
    .io_x_i(GenericAddSub16_io_x_i),
    .io_y_i(GenericAddSub16_io_y_i),
    .io_x_i_neg(GenericAddSub16_io_x_i_neg),
    .io_x_i_zero(GenericAddSub16_io_x_i_zero),
    .io_y_i_neg(GenericAddSub16_io_y_i_neg),
    .io_y_i_zero(GenericAddSub16_io_y_i_zero),
    .io_sum_o(GenericAddSub16_io_sum_o)
  );
  GenericAddSub16 GenericAddSub16_1 ( // @[DenseLayer.scala 29:29]
    .clock(GenericAddSub16_1_clock),
    .io_x_i(GenericAddSub16_1_io_x_i),
    .io_y_i(GenericAddSub16_1_io_y_i),
    .io_x_i_neg(GenericAddSub16_1_io_x_i_neg),
    .io_x_i_zero(GenericAddSub16_1_io_x_i_zero),
    .io_y_i_neg(GenericAddSub16_1_io_y_i_neg),
    .io_y_i_zero(GenericAddSub16_1_io_y_i_zero),
    .io_sum_o(GenericAddSub16_1_io_sum_o)
  );
  assign _T_12 = io_weights[0]; // @[DenseLayer.scala 25:35]
  assign _T_14 = _T_12 == 1'h0; // @[DenseLayer.scala 25:24]
  assign _T_15 = io_weights[1]; // @[DenseLayer.scala 26:33]
  assign _T_16 = io_weights[2]; // @[DenseLayer.scala 27:35]
  assign _T_18 = _T_16 == 1'h0; // @[DenseLayer.scala 27:24]
  assign _T_19 = io_weights[3]; // @[DenseLayer.scala 28:33]
  assign _T_20 = io_weights[4]; // @[DenseLayer.scala 25:35]
  assign _T_22 = _T_20 == 1'h0; // @[DenseLayer.scala 25:24]
  assign _T_23 = io_weights[5]; // @[DenseLayer.scala 26:33]
  assign _T_24 = io_weights[6]; // @[DenseLayer.scala 27:35]
  assign _T_26 = _T_24 == 1'h0; // @[DenseLayer.scala 27:24]
  assign _T_27 = io_weights[7]; // @[DenseLayer.scala 28:33]
  assign _T_28 = $signed(GenericAddSub16_io_sum_o) + $signed(GenericAddSub16_1_io_sum_o); // @[DenseLayer.scala 67:33]
  assign _T_29 = _T_28[15:0]; // @[DenseLayer.scala 67:33]
  assign _T_30 = $signed(_T_29); // @[DenseLayer.scala 67:33]
  assign io_sum = numsToSum_0;
  assign GenericAddSub16_clock = clock;
  assign GenericAddSub16_io_x_i = io_activations_0;
  assign GenericAddSub16_io_y_i = io_activations_1;
  assign GenericAddSub16_io_x_i_neg = _T_15;
  assign GenericAddSub16_io_x_i_zero = _T_14;
  assign GenericAddSub16_io_y_i_neg = _T_19;
  assign GenericAddSub16_io_y_i_zero = _T_18;
  assign GenericAddSub16_1_clock = clock;
  assign GenericAddSub16_1_io_x_i = io_activations_2;
  assign GenericAddSub16_1_io_y_i = io_activations_3;
  assign GenericAddSub16_1_io_x_i_neg = _T_23;
  assign GenericAddSub16_1_io_x_i_zero = _T_22;
  assign GenericAddSub16_1_io_y_i_neg = _T_27;
  assign GenericAddSub16_1_io_y_i_zero = _T_26;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  numsToSum_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    numsToSum_0 <= _T_30;
  end
endmodule
module DenseLayer(
  input         clock,
  input         reset,
  input         io_dataIn_valid,
  input  [15:0] io_dataIn_bits_0,
  input  [15:0] io_dataIn_bits_1,
  input  [15:0] io_dataIn_bits_2,
  input  [15:0] io_dataIn_bits_3,
  output        io_dataOut_valid,
  output [15:0] io_dataOut_bits_0,
  output [15:0] io_dataOut_bits_1,
  output [15:0] io_dataOut_bits_2,
  output [15:0] io_dataOut_bits_3,
  output [15:0] io_dataOut_bits_4,
  output [15:0] io_dataOut_bits_5,
  output [15:0] io_dataOut_bits_6,
  output [15:0] io_dataOut_bits_7,
  output [15:0] io_dataOut_bits_8,
  output [15:0] io_dataOut_bits_9,
  output [15:0] io_dataOut_bits_10,
  output [15:0] io_dataOut_bits_11,
  output [15:0] io_dataOut_bits_12,
  output [15:0] io_dataOut_bits_13,
  output [15:0] io_dataOut_bits_14,
  output [15:0] io_dataOut_bits_15,
  output [15:0] io_dataOut_bits_16,
  output [15:0] io_dataOut_bits_17,
  output [15:0] io_dataOut_bits_18,
  output [15:0] io_dataOut_bits_19,
  output [15:0] io_dataOut_bits_20,
  output [15:0] io_dataOut_bits_21,
  output [15:0] io_dataOut_bits_22,
  output [15:0] io_dataOut_bits_23,
  output [15:0] io_dataOut_bits_24,
  output [15:0] io_dataOut_bits_25,
  output [15:0] io_dataOut_bits_26,
  output [15:0] io_dataOut_bits_27,
  output [15:0] io_dataOut_bits_28,
  output [15:0] io_dataOut_bits_29,
  output [15:0] io_dataOut_bits_30,
  output [15:0] io_dataOut_bits_31,
  output [15:0] io_dataOut_bits_32,
  output [15:0] io_dataOut_bits_33,
  output [15:0] io_dataOut_bits_34,
  output [15:0] io_dataOut_bits_35,
  output [15:0] io_dataOut_bits_36,
  output [15:0] io_dataOut_bits_37,
  output [15:0] io_dataOut_bits_38,
  output [15:0] io_dataOut_bits_39,
  output [15:0] io_dataOut_bits_40,
  output [15:0] io_dataOut_bits_41,
  output [15:0] io_dataOut_bits_42,
  output [15:0] io_dataOut_bits_43,
  output [15:0] io_dataOut_bits_44,
  output [15:0] io_dataOut_bits_45,
  output [15:0] io_dataOut_bits_46,
  output [15:0] io_dataOut_bits_47,
  output [15:0] io_dataOut_bits_48,
  output [15:0] io_dataOut_bits_49,
  output [15:0] io_dataOut_bits_50,
  output [15:0] io_dataOut_bits_51,
  output [15:0] io_dataOut_bits_52,
  output [15:0] io_dataOut_bits_53,
  output [15:0] io_dataOut_bits_54,
  output [15:0] io_dataOut_bits_55,
  output [15:0] io_dataOut_bits_56,
  output [15:0] io_dataOut_bits_57,
  output [15:0] io_dataOut_bits_58,
  output [15:0] io_dataOut_bits_59,
  output [15:0] io_dataOut_bits_60,
  output [15:0] io_dataOut_bits_61,
  output [15:0] io_dataOut_bits_62,
  output [15:0] io_dataOut_bits_63,
  output [15:0] io_dataOut_bits_64,
  output [15:0] io_dataOut_bits_65,
  output [15:0] io_dataOut_bits_66,
  output [15:0] io_dataOut_bits_67,
  output [15:0] io_dataOut_bits_68,
  output [15:0] io_dataOut_bits_69,
  output [15:0] io_dataOut_bits_70,
  output [15:0] io_dataOut_bits_71,
  output [15:0] io_dataOut_bits_72,
  output [15:0] io_dataOut_bits_73,
  output [15:0] io_dataOut_bits_74,
  output [15:0] io_dataOut_bits_75,
  output [15:0] io_dataOut_bits_76,
  output [15:0] io_dataOut_bits_77,
  output [15:0] io_dataOut_bits_78,
  output [15:0] io_dataOut_bits_79,
  output [15:0] io_dataOut_bits_80,
  output [15:0] io_dataOut_bits_81,
  output [15:0] io_dataOut_bits_82,
  output [15:0] io_dataOut_bits_83,
  output [15:0] io_dataOut_bits_84,
  output [15:0] io_dataOut_bits_85,
  output [15:0] io_dataOut_bits_86,
  output [15:0] io_dataOut_bits_87,
  output [15:0] io_dataOut_bits_88,
  output [15:0] io_dataOut_bits_89,
  output [15:0] io_dataOut_bits_90,
  output [15:0] io_dataOut_bits_91,
  output [15:0] io_dataOut_bits_92,
  output [15:0] io_dataOut_bits_93,
  output [15:0] io_dataOut_bits_94,
  output [15:0] io_dataOut_bits_95,
  output [15:0] io_dataOut_bits_96,
  output [15:0] io_dataOut_bits_97,
  output [15:0] io_dataOut_bits_98,
  output [15:0] io_dataOut_bits_99,
  output [15:0] io_dataOut_bits_100,
  output [15:0] io_dataOut_bits_101,
  output [15:0] io_dataOut_bits_102,
  output [15:0] io_dataOut_bits_103,
  output [15:0] io_dataOut_bits_104,
  output [15:0] io_dataOut_bits_105,
  output [15:0] io_dataOut_bits_106,
  output [15:0] io_dataOut_bits_107,
  output [15:0] io_dataOut_bits_108,
  output [15:0] io_dataOut_bits_109,
  output [15:0] io_dataOut_bits_110,
  output [15:0] io_dataOut_bits_111,
  output [15:0] io_dataOut_bits_112,
  output [15:0] io_dataOut_bits_113,
  output [15:0] io_dataOut_bits_114,
  output [15:0] io_dataOut_bits_115,
  output [15:0] io_dataOut_bits_116,
  output [15:0] io_dataOut_bits_117,
  output [15:0] io_dataOut_bits_118,
  output [15:0] io_dataOut_bits_119,
  output [15:0] io_dataOut_bits_120,
  output [15:0] io_dataOut_bits_121,
  output [15:0] io_dataOut_bits_122,
  output [15:0] io_dataOut_bits_123,
  output [15:0] io_dataOut_bits_124,
  output [15:0] io_dataOut_bits_125,
  output [15:0] io_dataOut_bits_126,
  output [15:0] io_dataOut_bits_127
);
  reg [9:0] cntr; // @[DenseLayer.scala 88:21]
  reg [31:0] _RAND_0;
  wire [1023:0] weightsRAM_out; // @[DenseLayer.scala 96:34]
  wire [9:0] weightsRAM_readAddr; // @[DenseLayer.scala 96:34]
  wire  weightsRAM_clock; // @[DenseLayer.scala 96:34]
  reg [9:0] _T_293; // @[DenseLayer.scala 97:36]
  reg [31:0] _RAND_1;
  reg [15:0] currActs_0; // @[DenseLayer.scala 102:25]
  reg [31:0] _RAND_2;
  reg [15:0] currActs_1; // @[DenseLayer.scala 102:25]
  reg [31:0] _RAND_3;
  reg [15:0] currActs_2; // @[DenseLayer.scala 102:25]
  reg [31:0] _RAND_4;
  reg [15:0] currActs_3; // @[DenseLayer.scala 102:25]
  reg [31:0] _RAND_5;
  reg [7:0] _T_711_0; // @[Reg.scala 11:16]
  reg [31:0] _RAND_6;
  reg [7:0] _T_711_1; // @[Reg.scala 11:16]
  reg [31:0] _RAND_7;
  reg [7:0] _T_711_2; // @[Reg.scala 11:16]
  reg [31:0] _RAND_8;
  reg [7:0] _T_711_3; // @[Reg.scala 11:16]
  reg [31:0] _RAND_9;
  reg [7:0] _T_711_4; // @[Reg.scala 11:16]
  reg [31:0] _RAND_10;
  reg [7:0] _T_711_5; // @[Reg.scala 11:16]
  reg [31:0] _RAND_11;
  reg [7:0] _T_711_6; // @[Reg.scala 11:16]
  reg [31:0] _RAND_12;
  reg [7:0] _T_711_7; // @[Reg.scala 11:16]
  reg [31:0] _RAND_13;
  reg [7:0] _T_711_8; // @[Reg.scala 11:16]
  reg [31:0] _RAND_14;
  reg [7:0] _T_711_9; // @[Reg.scala 11:16]
  reg [31:0] _RAND_15;
  reg [7:0] _T_711_10; // @[Reg.scala 11:16]
  reg [31:0] _RAND_16;
  reg [7:0] _T_711_11; // @[Reg.scala 11:16]
  reg [31:0] _RAND_17;
  reg [7:0] _T_711_12; // @[Reg.scala 11:16]
  reg [31:0] _RAND_18;
  reg [7:0] _T_711_13; // @[Reg.scala 11:16]
  reg [31:0] _RAND_19;
  reg [7:0] _T_711_14; // @[Reg.scala 11:16]
  reg [31:0] _RAND_20;
  reg [7:0] _T_711_15; // @[Reg.scala 11:16]
  reg [31:0] _RAND_21;
  reg [7:0] _T_711_16; // @[Reg.scala 11:16]
  reg [31:0] _RAND_22;
  reg [7:0] _T_711_17; // @[Reg.scala 11:16]
  reg [31:0] _RAND_23;
  reg [7:0] _T_711_18; // @[Reg.scala 11:16]
  reg [31:0] _RAND_24;
  reg [7:0] _T_711_19; // @[Reg.scala 11:16]
  reg [31:0] _RAND_25;
  reg [7:0] _T_711_20; // @[Reg.scala 11:16]
  reg [31:0] _RAND_26;
  reg [7:0] _T_711_21; // @[Reg.scala 11:16]
  reg [31:0] _RAND_27;
  reg [7:0] _T_711_22; // @[Reg.scala 11:16]
  reg [31:0] _RAND_28;
  reg [7:0] _T_711_23; // @[Reg.scala 11:16]
  reg [31:0] _RAND_29;
  reg [7:0] _T_711_24; // @[Reg.scala 11:16]
  reg [31:0] _RAND_30;
  reg [7:0] _T_711_25; // @[Reg.scala 11:16]
  reg [31:0] _RAND_31;
  reg [7:0] _T_711_26; // @[Reg.scala 11:16]
  reg [31:0] _RAND_32;
  reg [7:0] _T_711_27; // @[Reg.scala 11:16]
  reg [31:0] _RAND_33;
  reg [7:0] _T_711_28; // @[Reg.scala 11:16]
  reg [31:0] _RAND_34;
  reg [7:0] _T_711_29; // @[Reg.scala 11:16]
  reg [31:0] _RAND_35;
  reg [7:0] _T_711_30; // @[Reg.scala 11:16]
  reg [31:0] _RAND_36;
  reg [7:0] _T_711_31; // @[Reg.scala 11:16]
  reg [31:0] _RAND_37;
  reg [7:0] _T_711_32; // @[Reg.scala 11:16]
  reg [31:0] _RAND_38;
  reg [7:0] _T_711_33; // @[Reg.scala 11:16]
  reg [31:0] _RAND_39;
  reg [7:0] _T_711_34; // @[Reg.scala 11:16]
  reg [31:0] _RAND_40;
  reg [7:0] _T_711_35; // @[Reg.scala 11:16]
  reg [31:0] _RAND_41;
  reg [7:0] _T_711_36; // @[Reg.scala 11:16]
  reg [31:0] _RAND_42;
  reg [7:0] _T_711_37; // @[Reg.scala 11:16]
  reg [31:0] _RAND_43;
  reg [7:0] _T_711_38; // @[Reg.scala 11:16]
  reg [31:0] _RAND_44;
  reg [7:0] _T_711_39; // @[Reg.scala 11:16]
  reg [31:0] _RAND_45;
  reg [7:0] _T_711_40; // @[Reg.scala 11:16]
  reg [31:0] _RAND_46;
  reg [7:0] _T_711_41; // @[Reg.scala 11:16]
  reg [31:0] _RAND_47;
  reg [7:0] _T_711_42; // @[Reg.scala 11:16]
  reg [31:0] _RAND_48;
  reg [7:0] _T_711_43; // @[Reg.scala 11:16]
  reg [31:0] _RAND_49;
  reg [7:0] _T_711_44; // @[Reg.scala 11:16]
  reg [31:0] _RAND_50;
  reg [7:0] _T_711_45; // @[Reg.scala 11:16]
  reg [31:0] _RAND_51;
  reg [7:0] _T_711_46; // @[Reg.scala 11:16]
  reg [31:0] _RAND_52;
  reg [7:0] _T_711_47; // @[Reg.scala 11:16]
  reg [31:0] _RAND_53;
  reg [7:0] _T_711_48; // @[Reg.scala 11:16]
  reg [31:0] _RAND_54;
  reg [7:0] _T_711_49; // @[Reg.scala 11:16]
  reg [31:0] _RAND_55;
  reg [7:0] _T_711_50; // @[Reg.scala 11:16]
  reg [31:0] _RAND_56;
  reg [7:0] _T_711_51; // @[Reg.scala 11:16]
  reg [31:0] _RAND_57;
  reg [7:0] _T_711_52; // @[Reg.scala 11:16]
  reg [31:0] _RAND_58;
  reg [7:0] _T_711_53; // @[Reg.scala 11:16]
  reg [31:0] _RAND_59;
  reg [7:0] _T_711_54; // @[Reg.scala 11:16]
  reg [31:0] _RAND_60;
  reg [7:0] _T_711_55; // @[Reg.scala 11:16]
  reg [31:0] _RAND_61;
  reg [7:0] _T_711_56; // @[Reg.scala 11:16]
  reg [31:0] _RAND_62;
  reg [7:0] _T_711_57; // @[Reg.scala 11:16]
  reg [31:0] _RAND_63;
  reg [7:0] _T_711_58; // @[Reg.scala 11:16]
  reg [31:0] _RAND_64;
  reg [7:0] _T_711_59; // @[Reg.scala 11:16]
  reg [31:0] _RAND_65;
  reg [7:0] _T_711_60; // @[Reg.scala 11:16]
  reg [31:0] _RAND_66;
  reg [7:0] _T_711_61; // @[Reg.scala 11:16]
  reg [31:0] _RAND_67;
  reg [7:0] _T_711_62; // @[Reg.scala 11:16]
  reg [31:0] _RAND_68;
  reg [7:0] _T_711_63; // @[Reg.scala 11:16]
  reg [31:0] _RAND_69;
  reg [7:0] _T_711_64; // @[Reg.scala 11:16]
  reg [31:0] _RAND_70;
  reg [7:0] _T_711_65; // @[Reg.scala 11:16]
  reg [31:0] _RAND_71;
  reg [7:0] _T_711_66; // @[Reg.scala 11:16]
  reg [31:0] _RAND_72;
  reg [7:0] _T_711_67; // @[Reg.scala 11:16]
  reg [31:0] _RAND_73;
  reg [7:0] _T_711_68; // @[Reg.scala 11:16]
  reg [31:0] _RAND_74;
  reg [7:0] _T_711_69; // @[Reg.scala 11:16]
  reg [31:0] _RAND_75;
  reg [7:0] _T_711_70; // @[Reg.scala 11:16]
  reg [31:0] _RAND_76;
  reg [7:0] _T_711_71; // @[Reg.scala 11:16]
  reg [31:0] _RAND_77;
  reg [7:0] _T_711_72; // @[Reg.scala 11:16]
  reg [31:0] _RAND_78;
  reg [7:0] _T_711_73; // @[Reg.scala 11:16]
  reg [31:0] _RAND_79;
  reg [7:0] _T_711_74; // @[Reg.scala 11:16]
  reg [31:0] _RAND_80;
  reg [7:0] _T_711_75; // @[Reg.scala 11:16]
  reg [31:0] _RAND_81;
  reg [7:0] _T_711_76; // @[Reg.scala 11:16]
  reg [31:0] _RAND_82;
  reg [7:0] _T_711_77; // @[Reg.scala 11:16]
  reg [31:0] _RAND_83;
  reg [7:0] _T_711_78; // @[Reg.scala 11:16]
  reg [31:0] _RAND_84;
  reg [7:0] _T_711_79; // @[Reg.scala 11:16]
  reg [31:0] _RAND_85;
  reg [7:0] _T_711_80; // @[Reg.scala 11:16]
  reg [31:0] _RAND_86;
  reg [7:0] _T_711_81; // @[Reg.scala 11:16]
  reg [31:0] _RAND_87;
  reg [7:0] _T_711_82; // @[Reg.scala 11:16]
  reg [31:0] _RAND_88;
  reg [7:0] _T_711_83; // @[Reg.scala 11:16]
  reg [31:0] _RAND_89;
  reg [7:0] _T_711_84; // @[Reg.scala 11:16]
  reg [31:0] _RAND_90;
  reg [7:0] _T_711_85; // @[Reg.scala 11:16]
  reg [31:0] _RAND_91;
  reg [7:0] _T_711_86; // @[Reg.scala 11:16]
  reg [31:0] _RAND_92;
  reg [7:0] _T_711_87; // @[Reg.scala 11:16]
  reg [31:0] _RAND_93;
  reg [7:0] _T_711_88; // @[Reg.scala 11:16]
  reg [31:0] _RAND_94;
  reg [7:0] _T_711_89; // @[Reg.scala 11:16]
  reg [31:0] _RAND_95;
  reg [7:0] _T_711_90; // @[Reg.scala 11:16]
  reg [31:0] _RAND_96;
  reg [7:0] _T_711_91; // @[Reg.scala 11:16]
  reg [31:0] _RAND_97;
  reg [7:0] _T_711_92; // @[Reg.scala 11:16]
  reg [31:0] _RAND_98;
  reg [7:0] _T_711_93; // @[Reg.scala 11:16]
  reg [31:0] _RAND_99;
  reg [7:0] _T_711_94; // @[Reg.scala 11:16]
  reg [31:0] _RAND_100;
  reg [7:0] _T_711_95; // @[Reg.scala 11:16]
  reg [31:0] _RAND_101;
  reg [7:0] _T_711_96; // @[Reg.scala 11:16]
  reg [31:0] _RAND_102;
  reg [7:0] _T_711_97; // @[Reg.scala 11:16]
  reg [31:0] _RAND_103;
  reg [7:0] _T_711_98; // @[Reg.scala 11:16]
  reg [31:0] _RAND_104;
  reg [7:0] _T_711_99; // @[Reg.scala 11:16]
  reg [31:0] _RAND_105;
  reg [7:0] _T_711_100; // @[Reg.scala 11:16]
  reg [31:0] _RAND_106;
  reg [7:0] _T_711_101; // @[Reg.scala 11:16]
  reg [31:0] _RAND_107;
  reg [7:0] _T_711_102; // @[Reg.scala 11:16]
  reg [31:0] _RAND_108;
  reg [7:0] _T_711_103; // @[Reg.scala 11:16]
  reg [31:0] _RAND_109;
  reg [7:0] _T_711_104; // @[Reg.scala 11:16]
  reg [31:0] _RAND_110;
  reg [7:0] _T_711_105; // @[Reg.scala 11:16]
  reg [31:0] _RAND_111;
  reg [7:0] _T_711_106; // @[Reg.scala 11:16]
  reg [31:0] _RAND_112;
  reg [7:0] _T_711_107; // @[Reg.scala 11:16]
  reg [31:0] _RAND_113;
  reg [7:0] _T_711_108; // @[Reg.scala 11:16]
  reg [31:0] _RAND_114;
  reg [7:0] _T_711_109; // @[Reg.scala 11:16]
  reg [31:0] _RAND_115;
  reg [7:0] _T_711_110; // @[Reg.scala 11:16]
  reg [31:0] _RAND_116;
  reg [7:0] _T_711_111; // @[Reg.scala 11:16]
  reg [31:0] _RAND_117;
  reg [7:0] _T_711_112; // @[Reg.scala 11:16]
  reg [31:0] _RAND_118;
  reg [7:0] _T_711_113; // @[Reg.scala 11:16]
  reg [31:0] _RAND_119;
  reg [7:0] _T_711_114; // @[Reg.scala 11:16]
  reg [31:0] _RAND_120;
  reg [7:0] _T_711_115; // @[Reg.scala 11:16]
  reg [31:0] _RAND_121;
  reg [7:0] _T_711_116; // @[Reg.scala 11:16]
  reg [31:0] _RAND_122;
  reg [7:0] _T_711_117; // @[Reg.scala 11:16]
  reg [31:0] _RAND_123;
  reg [7:0] _T_711_118; // @[Reg.scala 11:16]
  reg [31:0] _RAND_124;
  reg [7:0] _T_711_119; // @[Reg.scala 11:16]
  reg [31:0] _RAND_125;
  reg [7:0] _T_711_120; // @[Reg.scala 11:16]
  reg [31:0] _RAND_126;
  reg [7:0] _T_711_121; // @[Reg.scala 11:16]
  reg [31:0] _RAND_127;
  reg [7:0] _T_711_122; // @[Reg.scala 11:16]
  reg [31:0] _RAND_128;
  reg [7:0] _T_711_123; // @[Reg.scala 11:16]
  reg [31:0] _RAND_129;
  reg [7:0] _T_711_124; // @[Reg.scala 11:16]
  reg [31:0] _RAND_130;
  reg [7:0] _T_711_125; // @[Reg.scala 11:16]
  reg [31:0] _RAND_131;
  reg [7:0] _T_711_126; // @[Reg.scala 11:16]
  reg [31:0] _RAND_132;
  reg [7:0] _T_711_127; // @[Reg.scala 11:16]
  reg [31:0] _RAND_133;
  reg [7:0] delayWeights_0; // @[Reg.scala 11:16]
  reg [31:0] _RAND_134;
  reg [7:0] delayWeights_1; // @[Reg.scala 11:16]
  reg [31:0] _RAND_135;
  reg [7:0] delayWeights_2; // @[Reg.scala 11:16]
  reg [31:0] _RAND_136;
  reg [7:0] delayWeights_3; // @[Reg.scala 11:16]
  reg [31:0] _RAND_137;
  reg [7:0] delayWeights_4; // @[Reg.scala 11:16]
  reg [31:0] _RAND_138;
  reg [7:0] delayWeights_5; // @[Reg.scala 11:16]
  reg [31:0] _RAND_139;
  reg [7:0] delayWeights_6; // @[Reg.scala 11:16]
  reg [31:0] _RAND_140;
  reg [7:0] delayWeights_7; // @[Reg.scala 11:16]
  reg [31:0] _RAND_141;
  reg [7:0] delayWeights_8; // @[Reg.scala 11:16]
  reg [31:0] _RAND_142;
  reg [7:0] delayWeights_9; // @[Reg.scala 11:16]
  reg [31:0] _RAND_143;
  reg [7:0] delayWeights_10; // @[Reg.scala 11:16]
  reg [31:0] _RAND_144;
  reg [7:0] delayWeights_11; // @[Reg.scala 11:16]
  reg [31:0] _RAND_145;
  reg [7:0] delayWeights_12; // @[Reg.scala 11:16]
  reg [31:0] _RAND_146;
  reg [7:0] delayWeights_13; // @[Reg.scala 11:16]
  reg [31:0] _RAND_147;
  reg [7:0] delayWeights_14; // @[Reg.scala 11:16]
  reg [31:0] _RAND_148;
  reg [7:0] delayWeights_15; // @[Reg.scala 11:16]
  reg [31:0] _RAND_149;
  reg [7:0] delayWeights_16; // @[Reg.scala 11:16]
  reg [31:0] _RAND_150;
  reg [7:0] delayWeights_17; // @[Reg.scala 11:16]
  reg [31:0] _RAND_151;
  reg [7:0] delayWeights_18; // @[Reg.scala 11:16]
  reg [31:0] _RAND_152;
  reg [7:0] delayWeights_19; // @[Reg.scala 11:16]
  reg [31:0] _RAND_153;
  reg [7:0] delayWeights_20; // @[Reg.scala 11:16]
  reg [31:0] _RAND_154;
  reg [7:0] delayWeights_21; // @[Reg.scala 11:16]
  reg [31:0] _RAND_155;
  reg [7:0] delayWeights_22; // @[Reg.scala 11:16]
  reg [31:0] _RAND_156;
  reg [7:0] delayWeights_23; // @[Reg.scala 11:16]
  reg [31:0] _RAND_157;
  reg [7:0] delayWeights_24; // @[Reg.scala 11:16]
  reg [31:0] _RAND_158;
  reg [7:0] delayWeights_25; // @[Reg.scala 11:16]
  reg [31:0] _RAND_159;
  reg [7:0] delayWeights_26; // @[Reg.scala 11:16]
  reg [31:0] _RAND_160;
  reg [7:0] delayWeights_27; // @[Reg.scala 11:16]
  reg [31:0] _RAND_161;
  reg [7:0] delayWeights_28; // @[Reg.scala 11:16]
  reg [31:0] _RAND_162;
  reg [7:0] delayWeights_29; // @[Reg.scala 11:16]
  reg [31:0] _RAND_163;
  reg [7:0] delayWeights_30; // @[Reg.scala 11:16]
  reg [31:0] _RAND_164;
  reg [7:0] delayWeights_31; // @[Reg.scala 11:16]
  reg [31:0] _RAND_165;
  reg [7:0] delayWeights_32; // @[Reg.scala 11:16]
  reg [31:0] _RAND_166;
  reg [7:0] delayWeights_33; // @[Reg.scala 11:16]
  reg [31:0] _RAND_167;
  reg [7:0] delayWeights_34; // @[Reg.scala 11:16]
  reg [31:0] _RAND_168;
  reg [7:0] delayWeights_35; // @[Reg.scala 11:16]
  reg [31:0] _RAND_169;
  reg [7:0] delayWeights_36; // @[Reg.scala 11:16]
  reg [31:0] _RAND_170;
  reg [7:0] delayWeights_37; // @[Reg.scala 11:16]
  reg [31:0] _RAND_171;
  reg [7:0] delayWeights_38; // @[Reg.scala 11:16]
  reg [31:0] _RAND_172;
  reg [7:0] delayWeights_39; // @[Reg.scala 11:16]
  reg [31:0] _RAND_173;
  reg [7:0] delayWeights_40; // @[Reg.scala 11:16]
  reg [31:0] _RAND_174;
  reg [7:0] delayWeights_41; // @[Reg.scala 11:16]
  reg [31:0] _RAND_175;
  reg [7:0] delayWeights_42; // @[Reg.scala 11:16]
  reg [31:0] _RAND_176;
  reg [7:0] delayWeights_43; // @[Reg.scala 11:16]
  reg [31:0] _RAND_177;
  reg [7:0] delayWeights_44; // @[Reg.scala 11:16]
  reg [31:0] _RAND_178;
  reg [7:0] delayWeights_45; // @[Reg.scala 11:16]
  reg [31:0] _RAND_179;
  reg [7:0] delayWeights_46; // @[Reg.scala 11:16]
  reg [31:0] _RAND_180;
  reg [7:0] delayWeights_47; // @[Reg.scala 11:16]
  reg [31:0] _RAND_181;
  reg [7:0] delayWeights_48; // @[Reg.scala 11:16]
  reg [31:0] _RAND_182;
  reg [7:0] delayWeights_49; // @[Reg.scala 11:16]
  reg [31:0] _RAND_183;
  reg [7:0] delayWeights_50; // @[Reg.scala 11:16]
  reg [31:0] _RAND_184;
  reg [7:0] delayWeights_51; // @[Reg.scala 11:16]
  reg [31:0] _RAND_185;
  reg [7:0] delayWeights_52; // @[Reg.scala 11:16]
  reg [31:0] _RAND_186;
  reg [7:0] delayWeights_53; // @[Reg.scala 11:16]
  reg [31:0] _RAND_187;
  reg [7:0] delayWeights_54; // @[Reg.scala 11:16]
  reg [31:0] _RAND_188;
  reg [7:0] delayWeights_55; // @[Reg.scala 11:16]
  reg [31:0] _RAND_189;
  reg [7:0] delayWeights_56; // @[Reg.scala 11:16]
  reg [31:0] _RAND_190;
  reg [7:0] delayWeights_57; // @[Reg.scala 11:16]
  reg [31:0] _RAND_191;
  reg [7:0] delayWeights_58; // @[Reg.scala 11:16]
  reg [31:0] _RAND_192;
  reg [7:0] delayWeights_59; // @[Reg.scala 11:16]
  reg [31:0] _RAND_193;
  reg [7:0] delayWeights_60; // @[Reg.scala 11:16]
  reg [31:0] _RAND_194;
  reg [7:0] delayWeights_61; // @[Reg.scala 11:16]
  reg [31:0] _RAND_195;
  reg [7:0] delayWeights_62; // @[Reg.scala 11:16]
  reg [31:0] _RAND_196;
  reg [7:0] delayWeights_63; // @[Reg.scala 11:16]
  reg [31:0] _RAND_197;
  reg [7:0] delayWeights_64; // @[Reg.scala 11:16]
  reg [31:0] _RAND_198;
  reg [7:0] delayWeights_65; // @[Reg.scala 11:16]
  reg [31:0] _RAND_199;
  reg [7:0] delayWeights_66; // @[Reg.scala 11:16]
  reg [31:0] _RAND_200;
  reg [7:0] delayWeights_67; // @[Reg.scala 11:16]
  reg [31:0] _RAND_201;
  reg [7:0] delayWeights_68; // @[Reg.scala 11:16]
  reg [31:0] _RAND_202;
  reg [7:0] delayWeights_69; // @[Reg.scala 11:16]
  reg [31:0] _RAND_203;
  reg [7:0] delayWeights_70; // @[Reg.scala 11:16]
  reg [31:0] _RAND_204;
  reg [7:0] delayWeights_71; // @[Reg.scala 11:16]
  reg [31:0] _RAND_205;
  reg [7:0] delayWeights_72; // @[Reg.scala 11:16]
  reg [31:0] _RAND_206;
  reg [7:0] delayWeights_73; // @[Reg.scala 11:16]
  reg [31:0] _RAND_207;
  reg [7:0] delayWeights_74; // @[Reg.scala 11:16]
  reg [31:0] _RAND_208;
  reg [7:0] delayWeights_75; // @[Reg.scala 11:16]
  reg [31:0] _RAND_209;
  reg [7:0] delayWeights_76; // @[Reg.scala 11:16]
  reg [31:0] _RAND_210;
  reg [7:0] delayWeights_77; // @[Reg.scala 11:16]
  reg [31:0] _RAND_211;
  reg [7:0] delayWeights_78; // @[Reg.scala 11:16]
  reg [31:0] _RAND_212;
  reg [7:0] delayWeights_79; // @[Reg.scala 11:16]
  reg [31:0] _RAND_213;
  reg [7:0] delayWeights_80; // @[Reg.scala 11:16]
  reg [31:0] _RAND_214;
  reg [7:0] delayWeights_81; // @[Reg.scala 11:16]
  reg [31:0] _RAND_215;
  reg [7:0] delayWeights_82; // @[Reg.scala 11:16]
  reg [31:0] _RAND_216;
  reg [7:0] delayWeights_83; // @[Reg.scala 11:16]
  reg [31:0] _RAND_217;
  reg [7:0] delayWeights_84; // @[Reg.scala 11:16]
  reg [31:0] _RAND_218;
  reg [7:0] delayWeights_85; // @[Reg.scala 11:16]
  reg [31:0] _RAND_219;
  reg [7:0] delayWeights_86; // @[Reg.scala 11:16]
  reg [31:0] _RAND_220;
  reg [7:0] delayWeights_87; // @[Reg.scala 11:16]
  reg [31:0] _RAND_221;
  reg [7:0] delayWeights_88; // @[Reg.scala 11:16]
  reg [31:0] _RAND_222;
  reg [7:0] delayWeights_89; // @[Reg.scala 11:16]
  reg [31:0] _RAND_223;
  reg [7:0] delayWeights_90; // @[Reg.scala 11:16]
  reg [31:0] _RAND_224;
  reg [7:0] delayWeights_91; // @[Reg.scala 11:16]
  reg [31:0] _RAND_225;
  reg [7:0] delayWeights_92; // @[Reg.scala 11:16]
  reg [31:0] _RAND_226;
  reg [7:0] delayWeights_93; // @[Reg.scala 11:16]
  reg [31:0] _RAND_227;
  reg [7:0] delayWeights_94; // @[Reg.scala 11:16]
  reg [31:0] _RAND_228;
  reg [7:0] delayWeights_95; // @[Reg.scala 11:16]
  reg [31:0] _RAND_229;
  reg [7:0] delayWeights_96; // @[Reg.scala 11:16]
  reg [31:0] _RAND_230;
  reg [7:0] delayWeights_97; // @[Reg.scala 11:16]
  reg [31:0] _RAND_231;
  reg [7:0] delayWeights_98; // @[Reg.scala 11:16]
  reg [31:0] _RAND_232;
  reg [7:0] delayWeights_99; // @[Reg.scala 11:16]
  reg [31:0] _RAND_233;
  reg [7:0] delayWeights_100; // @[Reg.scala 11:16]
  reg [31:0] _RAND_234;
  reg [7:0] delayWeights_101; // @[Reg.scala 11:16]
  reg [31:0] _RAND_235;
  reg [7:0] delayWeights_102; // @[Reg.scala 11:16]
  reg [31:0] _RAND_236;
  reg [7:0] delayWeights_103; // @[Reg.scala 11:16]
  reg [31:0] _RAND_237;
  reg [7:0] delayWeights_104; // @[Reg.scala 11:16]
  reg [31:0] _RAND_238;
  reg [7:0] delayWeights_105; // @[Reg.scala 11:16]
  reg [31:0] _RAND_239;
  reg [7:0] delayWeights_106; // @[Reg.scala 11:16]
  reg [31:0] _RAND_240;
  reg [7:0] delayWeights_107; // @[Reg.scala 11:16]
  reg [31:0] _RAND_241;
  reg [7:0] delayWeights_108; // @[Reg.scala 11:16]
  reg [31:0] _RAND_242;
  reg [7:0] delayWeights_109; // @[Reg.scala 11:16]
  reg [31:0] _RAND_243;
  reg [7:0] delayWeights_110; // @[Reg.scala 11:16]
  reg [31:0] _RAND_244;
  reg [7:0] delayWeights_111; // @[Reg.scala 11:16]
  reg [31:0] _RAND_245;
  reg [7:0] delayWeights_112; // @[Reg.scala 11:16]
  reg [31:0] _RAND_246;
  reg [7:0] delayWeights_113; // @[Reg.scala 11:16]
  reg [31:0] _RAND_247;
  reg [7:0] delayWeights_114; // @[Reg.scala 11:16]
  reg [31:0] _RAND_248;
  reg [7:0] delayWeights_115; // @[Reg.scala 11:16]
  reg [31:0] _RAND_249;
  reg [7:0] delayWeights_116; // @[Reg.scala 11:16]
  reg [31:0] _RAND_250;
  reg [7:0] delayWeights_117; // @[Reg.scala 11:16]
  reg [31:0] _RAND_251;
  reg [7:0] delayWeights_118; // @[Reg.scala 11:16]
  reg [31:0] _RAND_252;
  reg [7:0] delayWeights_119; // @[Reg.scala 11:16]
  reg [31:0] _RAND_253;
  reg [7:0] delayWeights_120; // @[Reg.scala 11:16]
  reg [31:0] _RAND_254;
  reg [7:0] delayWeights_121; // @[Reg.scala 11:16]
  reg [31:0] _RAND_255;
  reg [7:0] delayWeights_122; // @[Reg.scala 11:16]
  reg [31:0] _RAND_256;
  reg [7:0] delayWeights_123; // @[Reg.scala 11:16]
  reg [31:0] _RAND_257;
  reg [7:0] delayWeights_124; // @[Reg.scala 11:16]
  reg [31:0] _RAND_258;
  reg [7:0] delayWeights_125; // @[Reg.scala 11:16]
  reg [31:0] _RAND_259;
  reg [7:0] delayWeights_126; // @[Reg.scala 11:16]
  reg [31:0] _RAND_260;
  reg [7:0] delayWeights_127; // @[Reg.scala 11:16]
  reg [31:0] _RAND_261;
  wire  FanoutAWS_clock; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_in; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_0; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_1; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_2; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_3; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_4; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_5; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_6; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_7; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_8; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_9; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_10; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_11; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_12; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_13; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_14; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_15; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_16; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_17; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_18; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_19; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_20; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_21; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_22; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_23; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_24; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_25; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_26; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_27; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_28; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_29; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_30; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_31; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_32; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_33; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_34; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_35; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_36; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_37; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_38; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_39; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_40; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_41; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_42; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_43; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_44; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_45; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_46; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_47; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_48; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_49; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_50; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_51; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_52; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_53; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_54; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_55; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_56; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_57; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_58; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_59; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_60; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_61; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_62; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_63; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_64; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_65; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_66; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_67; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_68; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_69; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_70; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_71; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_72; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_73; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_74; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_75; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_76; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_77; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_78; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_79; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_80; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_81; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_82; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_83; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_84; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_85; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_86; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_87; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_88; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_89; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_90; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_91; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_92; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_93; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_94; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_95; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_96; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_97; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_98; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_99; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_100; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_101; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_102; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_103; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_104; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_105; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_106; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_107; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_108; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_109; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_110; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_111; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_112; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_113; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_114; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_115; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_116; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_117; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_118; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_119; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_120; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_121; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_122; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_123; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_124; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_125; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_126; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_127; // @[FanoutAWS.scala 16:26]
  wire  FanoutAWS_1_clock; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_in; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_0; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_1; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_2; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_3; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_4; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_5; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_6; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_7; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_8; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_9; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_10; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_11; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_12; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_13; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_14; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_15; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_16; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_17; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_18; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_19; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_20; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_21; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_22; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_23; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_24; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_25; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_26; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_27; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_28; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_29; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_30; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_31; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_32; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_33; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_34; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_35; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_36; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_37; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_38; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_39; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_40; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_41; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_42; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_43; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_44; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_45; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_46; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_47; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_48; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_49; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_50; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_51; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_52; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_53; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_54; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_55; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_56; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_57; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_58; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_59; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_60; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_61; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_62; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_63; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_64; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_65; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_66; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_67; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_68; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_69; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_70; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_71; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_72; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_73; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_74; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_75; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_76; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_77; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_78; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_79; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_80; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_81; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_82; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_83; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_84; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_85; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_86; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_87; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_88; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_89; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_90; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_91; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_92; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_93; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_94; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_95; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_96; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_97; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_98; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_99; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_100; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_101; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_102; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_103; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_104; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_105; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_106; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_107; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_108; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_109; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_110; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_111; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_112; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_113; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_114; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_115; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_116; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_117; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_118; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_119; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_120; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_121; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_122; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_123; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_124; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_125; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_126; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_1_io_out_127; // @[FanoutAWS.scala 16:26]
  wire  FanoutAWS_2_clock; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_in; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_0; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_1; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_2; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_3; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_4; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_5; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_6; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_7; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_8; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_9; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_10; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_11; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_12; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_13; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_14; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_15; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_16; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_17; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_18; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_19; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_20; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_21; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_22; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_23; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_24; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_25; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_26; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_27; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_28; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_29; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_30; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_31; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_32; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_33; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_34; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_35; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_36; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_37; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_38; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_39; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_40; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_41; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_42; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_43; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_44; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_45; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_46; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_47; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_48; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_49; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_50; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_51; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_52; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_53; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_54; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_55; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_56; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_57; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_58; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_59; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_60; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_61; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_62; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_63; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_64; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_65; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_66; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_67; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_68; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_69; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_70; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_71; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_72; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_73; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_74; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_75; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_76; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_77; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_78; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_79; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_80; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_81; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_82; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_83; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_84; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_85; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_86; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_87; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_88; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_89; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_90; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_91; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_92; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_93; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_94; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_95; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_96; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_97; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_98; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_99; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_100; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_101; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_102; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_103; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_104; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_105; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_106; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_107; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_108; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_109; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_110; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_111; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_112; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_113; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_114; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_115; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_116; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_117; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_118; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_119; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_120; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_121; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_122; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_123; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_124; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_125; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_126; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_2_io_out_127; // @[FanoutAWS.scala 16:26]
  wire  FanoutAWS_3_clock; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_in; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_0; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_1; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_2; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_3; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_4; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_5; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_6; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_7; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_8; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_9; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_10; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_11; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_12; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_13; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_14; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_15; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_16; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_17; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_18; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_19; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_20; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_21; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_22; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_23; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_24; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_25; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_26; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_27; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_28; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_29; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_30; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_31; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_32; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_33; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_34; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_35; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_36; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_37; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_38; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_39; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_40; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_41; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_42; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_43; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_44; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_45; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_46; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_47; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_48; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_49; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_50; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_51; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_52; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_53; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_54; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_55; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_56; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_57; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_58; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_59; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_60; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_61; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_62; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_63; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_64; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_65; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_66; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_67; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_68; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_69; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_70; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_71; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_72; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_73; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_74; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_75; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_76; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_77; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_78; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_79; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_80; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_81; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_82; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_83; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_84; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_85; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_86; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_87; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_88; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_89; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_90; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_91; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_92; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_93; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_94; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_95; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_96; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_97; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_98; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_99; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_100; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_101; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_102; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_103; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_104; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_105; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_106; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_107; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_108; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_109; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_110; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_111; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_112; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_113; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_114; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_115; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_116; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_117; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_118; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_119; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_120; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_121; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_122; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_123; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_124; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_125; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_126; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_3_io_out_127; // @[FanoutAWS.scala 16:26]
  wire  MultiplyAccumulate_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_1_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_1_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_1_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_1_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_1_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_1_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_1_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_2_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_2_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_2_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_2_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_2_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_2_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_2_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_3_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_3_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_3_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_3_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_3_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_3_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_3_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_4_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_4_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_4_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_4_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_4_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_4_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_4_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_5_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_5_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_5_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_5_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_5_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_5_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_5_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_6_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_6_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_6_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_6_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_6_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_6_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_6_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_7_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_7_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_7_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_7_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_7_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_7_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_7_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_8_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_8_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_8_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_8_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_8_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_8_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_8_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_9_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_9_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_9_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_9_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_9_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_9_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_9_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_10_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_10_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_10_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_10_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_10_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_10_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_10_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_11_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_11_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_11_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_11_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_11_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_11_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_11_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_12_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_12_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_12_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_12_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_12_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_12_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_12_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_13_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_13_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_13_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_13_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_13_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_13_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_13_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_14_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_14_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_14_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_14_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_14_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_14_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_14_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_15_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_15_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_15_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_15_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_15_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_15_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_15_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_16_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_16_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_16_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_16_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_16_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_16_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_16_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_17_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_17_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_17_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_17_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_17_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_17_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_17_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_18_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_18_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_18_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_18_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_18_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_18_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_18_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_19_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_19_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_19_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_19_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_19_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_19_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_19_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_20_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_20_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_20_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_20_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_20_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_20_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_20_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_21_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_21_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_21_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_21_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_21_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_21_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_21_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_22_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_22_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_22_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_22_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_22_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_22_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_22_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_23_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_23_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_23_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_23_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_23_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_23_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_23_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_24_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_24_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_24_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_24_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_24_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_24_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_24_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_25_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_25_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_25_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_25_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_25_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_25_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_25_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_26_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_26_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_26_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_26_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_26_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_26_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_26_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_27_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_27_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_27_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_27_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_27_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_27_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_27_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_28_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_28_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_28_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_28_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_28_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_28_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_28_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_29_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_29_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_29_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_29_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_29_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_29_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_29_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_30_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_30_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_30_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_30_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_30_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_30_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_30_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_31_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_31_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_31_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_31_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_31_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_31_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_31_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_32_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_32_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_32_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_32_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_32_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_32_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_32_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_33_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_33_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_33_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_33_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_33_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_33_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_33_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_34_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_34_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_34_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_34_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_34_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_34_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_34_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_35_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_35_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_35_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_35_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_35_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_35_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_35_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_36_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_36_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_36_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_36_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_36_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_36_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_36_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_37_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_37_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_37_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_37_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_37_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_37_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_37_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_38_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_38_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_38_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_38_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_38_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_38_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_38_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_39_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_39_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_39_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_39_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_39_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_39_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_39_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_40_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_40_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_40_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_40_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_40_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_40_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_40_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_41_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_41_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_41_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_41_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_41_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_41_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_41_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_42_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_42_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_42_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_42_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_42_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_42_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_42_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_43_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_43_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_43_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_43_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_43_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_43_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_43_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_44_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_44_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_44_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_44_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_44_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_44_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_44_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_45_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_45_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_45_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_45_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_45_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_45_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_45_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_46_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_46_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_46_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_46_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_46_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_46_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_46_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_47_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_47_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_47_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_47_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_47_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_47_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_47_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_48_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_48_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_48_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_48_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_48_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_48_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_48_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_49_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_49_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_49_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_49_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_49_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_49_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_49_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_50_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_50_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_50_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_50_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_50_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_50_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_50_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_51_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_51_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_51_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_51_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_51_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_51_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_51_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_52_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_52_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_52_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_52_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_52_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_52_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_52_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_53_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_53_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_53_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_53_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_53_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_53_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_53_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_54_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_54_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_54_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_54_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_54_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_54_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_54_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_55_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_55_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_55_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_55_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_55_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_55_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_55_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_56_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_56_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_56_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_56_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_56_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_56_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_56_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_57_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_57_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_57_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_57_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_57_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_57_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_57_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_58_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_58_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_58_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_58_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_58_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_58_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_58_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_59_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_59_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_59_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_59_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_59_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_59_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_59_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_60_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_60_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_60_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_60_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_60_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_60_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_60_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_61_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_61_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_61_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_61_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_61_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_61_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_61_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_62_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_62_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_62_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_62_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_62_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_62_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_62_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_63_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_63_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_63_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_63_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_63_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_63_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_63_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_64_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_64_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_64_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_64_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_64_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_64_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_64_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_65_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_65_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_65_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_65_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_65_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_65_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_65_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_66_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_66_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_66_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_66_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_66_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_66_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_66_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_67_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_67_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_67_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_67_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_67_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_67_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_67_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_68_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_68_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_68_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_68_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_68_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_68_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_68_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_69_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_69_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_69_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_69_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_69_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_69_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_69_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_70_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_70_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_70_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_70_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_70_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_70_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_70_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_71_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_71_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_71_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_71_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_71_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_71_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_71_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_72_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_72_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_72_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_72_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_72_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_72_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_72_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_73_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_73_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_73_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_73_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_73_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_73_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_73_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_74_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_74_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_74_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_74_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_74_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_74_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_74_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_75_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_75_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_75_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_75_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_75_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_75_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_75_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_76_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_76_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_76_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_76_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_76_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_76_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_76_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_77_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_77_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_77_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_77_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_77_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_77_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_77_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_78_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_78_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_78_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_78_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_78_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_78_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_78_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_79_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_79_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_79_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_79_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_79_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_79_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_79_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_80_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_80_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_80_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_80_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_80_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_80_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_80_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_81_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_81_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_81_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_81_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_81_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_81_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_81_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_82_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_82_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_82_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_82_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_82_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_82_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_82_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_83_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_83_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_83_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_83_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_83_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_83_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_83_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_84_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_84_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_84_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_84_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_84_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_84_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_84_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_85_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_85_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_85_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_85_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_85_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_85_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_85_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_86_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_86_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_86_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_86_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_86_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_86_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_86_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_87_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_87_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_87_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_87_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_87_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_87_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_87_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_88_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_88_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_88_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_88_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_88_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_88_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_88_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_89_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_89_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_89_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_89_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_89_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_89_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_89_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_90_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_90_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_90_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_90_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_90_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_90_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_90_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_91_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_91_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_91_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_91_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_91_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_91_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_91_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_92_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_92_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_92_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_92_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_92_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_92_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_92_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_93_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_93_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_93_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_93_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_93_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_93_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_93_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_94_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_94_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_94_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_94_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_94_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_94_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_94_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_95_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_95_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_95_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_95_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_95_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_95_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_95_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_96_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_96_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_96_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_96_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_96_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_96_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_96_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_97_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_97_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_97_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_97_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_97_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_97_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_97_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_98_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_98_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_98_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_98_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_98_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_98_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_98_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_99_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_99_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_99_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_99_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_99_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_99_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_99_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_100_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_100_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_100_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_100_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_100_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_100_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_100_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_101_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_101_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_101_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_101_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_101_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_101_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_101_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_102_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_102_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_102_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_102_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_102_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_102_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_102_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_103_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_103_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_103_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_103_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_103_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_103_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_103_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_104_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_104_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_104_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_104_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_104_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_104_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_104_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_105_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_105_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_105_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_105_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_105_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_105_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_105_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_106_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_106_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_106_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_106_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_106_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_106_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_106_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_107_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_107_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_107_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_107_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_107_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_107_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_107_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_108_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_108_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_108_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_108_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_108_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_108_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_108_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_109_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_109_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_109_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_109_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_109_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_109_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_109_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_110_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_110_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_110_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_110_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_110_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_110_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_110_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_111_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_111_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_111_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_111_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_111_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_111_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_111_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_112_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_112_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_112_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_112_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_112_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_112_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_112_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_113_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_113_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_113_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_113_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_113_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_113_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_113_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_114_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_114_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_114_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_114_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_114_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_114_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_114_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_115_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_115_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_115_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_115_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_115_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_115_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_115_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_116_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_116_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_116_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_116_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_116_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_116_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_116_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_117_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_117_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_117_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_117_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_117_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_117_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_117_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_118_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_118_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_118_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_118_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_118_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_118_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_118_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_119_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_119_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_119_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_119_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_119_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_119_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_119_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_120_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_120_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_120_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_120_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_120_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_120_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_120_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_121_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_121_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_121_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_121_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_121_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_121_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_121_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_122_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_122_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_122_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_122_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_122_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_122_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_122_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_123_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_123_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_123_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_123_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_123_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_123_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_123_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_124_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_124_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_124_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_124_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_124_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_124_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_124_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_125_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_125_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_125_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_125_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_125_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_125_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_125_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_126_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_126_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_126_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_126_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_126_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_126_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_126_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_127_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_127_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_127_io_activations_1; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_127_io_activations_2; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_127_io_activations_3; // @[DenseLayer.scala 111:21]
  wire [7:0] MultiplyAccumulate_127_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_127_io_sum; // @[DenseLayer.scala 111:21]
  reg [15:0] cummulativeSums_0; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_262;
  reg [15:0] cummulativeSums_1; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_263;
  reg [15:0] cummulativeSums_2; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_264;
  reg [15:0] cummulativeSums_3; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_265;
  reg [15:0] cummulativeSums_4; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_266;
  reg [15:0] cummulativeSums_5; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_267;
  reg [15:0] cummulativeSums_6; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_268;
  reg [15:0] cummulativeSums_7; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_269;
  reg [15:0] cummulativeSums_8; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_270;
  reg [15:0] cummulativeSums_9; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_271;
  reg [15:0] cummulativeSums_10; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_272;
  reg [15:0] cummulativeSums_11; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_273;
  reg [15:0] cummulativeSums_12; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_274;
  reg [15:0] cummulativeSums_13; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_275;
  reg [15:0] cummulativeSums_14; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_276;
  reg [15:0] cummulativeSums_15; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_277;
  reg [15:0] cummulativeSums_16; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_278;
  reg [15:0] cummulativeSums_17; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_279;
  reg [15:0] cummulativeSums_18; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_280;
  reg [15:0] cummulativeSums_19; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_281;
  reg [15:0] cummulativeSums_20; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_282;
  reg [15:0] cummulativeSums_21; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_283;
  reg [15:0] cummulativeSums_22; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_284;
  reg [15:0] cummulativeSums_23; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_285;
  reg [15:0] cummulativeSums_24; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_286;
  reg [15:0] cummulativeSums_25; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_287;
  reg [15:0] cummulativeSums_26; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_288;
  reg [15:0] cummulativeSums_27; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_289;
  reg [15:0] cummulativeSums_28; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_290;
  reg [15:0] cummulativeSums_29; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_291;
  reg [15:0] cummulativeSums_30; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_292;
  reg [15:0] cummulativeSums_31; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_293;
  reg [15:0] cummulativeSums_32; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_294;
  reg [15:0] cummulativeSums_33; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_295;
  reg [15:0] cummulativeSums_34; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_296;
  reg [15:0] cummulativeSums_35; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_297;
  reg [15:0] cummulativeSums_36; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_298;
  reg [15:0] cummulativeSums_37; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_299;
  reg [15:0] cummulativeSums_38; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_300;
  reg [15:0] cummulativeSums_39; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_301;
  reg [15:0] cummulativeSums_40; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_302;
  reg [15:0] cummulativeSums_41; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_303;
  reg [15:0] cummulativeSums_42; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_304;
  reg [15:0] cummulativeSums_43; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_305;
  reg [15:0] cummulativeSums_44; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_306;
  reg [15:0] cummulativeSums_45; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_307;
  reg [15:0] cummulativeSums_46; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_308;
  reg [15:0] cummulativeSums_47; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_309;
  reg [15:0] cummulativeSums_48; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_310;
  reg [15:0] cummulativeSums_49; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_311;
  reg [15:0] cummulativeSums_50; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_312;
  reg [15:0] cummulativeSums_51; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_313;
  reg [15:0] cummulativeSums_52; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_314;
  reg [15:0] cummulativeSums_53; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_315;
  reg [15:0] cummulativeSums_54; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_316;
  reg [15:0] cummulativeSums_55; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_317;
  reg [15:0] cummulativeSums_56; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_318;
  reg [15:0] cummulativeSums_57; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_319;
  reg [15:0] cummulativeSums_58; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_320;
  reg [15:0] cummulativeSums_59; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_321;
  reg [15:0] cummulativeSums_60; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_322;
  reg [15:0] cummulativeSums_61; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_323;
  reg [15:0] cummulativeSums_62; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_324;
  reg [15:0] cummulativeSums_63; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_325;
  reg [15:0] cummulativeSums_64; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_326;
  reg [15:0] cummulativeSums_65; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_327;
  reg [15:0] cummulativeSums_66; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_328;
  reg [15:0] cummulativeSums_67; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_329;
  reg [15:0] cummulativeSums_68; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_330;
  reg [15:0] cummulativeSums_69; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_331;
  reg [15:0] cummulativeSums_70; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_332;
  reg [15:0] cummulativeSums_71; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_333;
  reg [15:0] cummulativeSums_72; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_334;
  reg [15:0] cummulativeSums_73; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_335;
  reg [15:0] cummulativeSums_74; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_336;
  reg [15:0] cummulativeSums_75; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_337;
  reg [15:0] cummulativeSums_76; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_338;
  reg [15:0] cummulativeSums_77; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_339;
  reg [15:0] cummulativeSums_78; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_340;
  reg [15:0] cummulativeSums_79; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_341;
  reg [15:0] cummulativeSums_80; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_342;
  reg [15:0] cummulativeSums_81; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_343;
  reg [15:0] cummulativeSums_82; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_344;
  reg [15:0] cummulativeSums_83; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_345;
  reg [15:0] cummulativeSums_84; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_346;
  reg [15:0] cummulativeSums_85; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_347;
  reg [15:0] cummulativeSums_86; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_348;
  reg [15:0] cummulativeSums_87; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_349;
  reg [15:0] cummulativeSums_88; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_350;
  reg [15:0] cummulativeSums_89; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_351;
  reg [15:0] cummulativeSums_90; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_352;
  reg [15:0] cummulativeSums_91; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_353;
  reg [15:0] cummulativeSums_92; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_354;
  reg [15:0] cummulativeSums_93; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_355;
  reg [15:0] cummulativeSums_94; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_356;
  reg [15:0] cummulativeSums_95; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_357;
  reg [15:0] cummulativeSums_96; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_358;
  reg [15:0] cummulativeSums_97; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_359;
  reg [15:0] cummulativeSums_98; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_360;
  reg [15:0] cummulativeSums_99; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_361;
  reg [15:0] cummulativeSums_100; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_362;
  reg [15:0] cummulativeSums_101; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_363;
  reg [15:0] cummulativeSums_102; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_364;
  reg [15:0] cummulativeSums_103; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_365;
  reg [15:0] cummulativeSums_104; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_366;
  reg [15:0] cummulativeSums_105; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_367;
  reg [15:0] cummulativeSums_106; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_368;
  reg [15:0] cummulativeSums_107; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_369;
  reg [15:0] cummulativeSums_108; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_370;
  reg [15:0] cummulativeSums_109; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_371;
  reg [15:0] cummulativeSums_110; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_372;
  reg [15:0] cummulativeSums_111; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_373;
  reg [15:0] cummulativeSums_112; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_374;
  reg [15:0] cummulativeSums_113; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_375;
  reg [15:0] cummulativeSums_114; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_376;
  reg [15:0] cummulativeSums_115; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_377;
  reg [15:0] cummulativeSums_116; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_378;
  reg [15:0] cummulativeSums_117; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_379;
  reg [15:0] cummulativeSums_118; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_380;
  reg [15:0] cummulativeSums_119; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_381;
  reg [15:0] cummulativeSums_120; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_382;
  reg [15:0] cummulativeSums_121; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_383;
  reg [15:0] cummulativeSums_122; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_384;
  reg [15:0] cummulativeSums_123; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_385;
  reg [15:0] cummulativeSums_124; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_386;
  reg [15:0] cummulativeSums_125; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_387;
  reg [15:0] cummulativeSums_126; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_388;
  reg [15:0] cummulativeSums_127; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_389;
  reg  _T_2401; // @[Reg.scala 11:16]
  reg [31:0] _RAND_390;
  reg  _T_2403; // @[Reg.scala 11:16]
  reg [31:0] _RAND_391;
  reg  _T_2405; // @[Reg.scala 11:16]
  reg [31:0] _RAND_392;
  reg  _T_2407; // @[Reg.scala 11:16]
  reg [31:0] _RAND_393;
  reg  _T_2409; // @[Reg.scala 11:16]
  reg [31:0] _RAND_394;
  reg  _T_2411; // @[Reg.scala 11:16]
  reg [31:0] _RAND_395;
  reg  rst; // @[Reg.scala 11:16]
  reg [31:0] _RAND_396;
  reg  done; // @[DenseLayer.scala 122:21]
  reg [31:0] _RAND_397;
  reg  _T_2422; // @[Reg.scala 11:16]
  reg [31:0] _RAND_398;
  reg  _T_2424; // @[Reg.scala 11:16]
  reg [31:0] _RAND_399;
  reg  _T_2426; // @[Reg.scala 11:16]
  reg [31:0] _RAND_400;
  reg  _T_2428; // @[Reg.scala 11:16]
  reg [31:0] _RAND_401;
  reg  _T_2430; // @[Reg.scala 11:16]
  reg [31:0] _RAND_402;
  reg  _T_2432; // @[Reg.scala 11:16]
  reg [31:0] _RAND_403;
  reg  vld; // @[Reg.scala 11:16]
  reg [31:0] _RAND_404;
  wire [10:0] _T_158; // @[DenseLayer.scala 90:18]
  wire [9:0] _T_159; // @[DenseLayer.scala 90:18]
  wire [9:0] _GEN_0; // @[DenseLayer.scala 89:28]
  wire [7:0] currWeights_0; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_1; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_2; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_3; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_4; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_5; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_6; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_7; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_8; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_9; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_10; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_11; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_12; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_13; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_14; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_15; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_16; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_17; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_18; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_19; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_20; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_21; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_22; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_23; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_24; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_25; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_26; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_27; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_28; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_29; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_30; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_31; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_32; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_33; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_34; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_35; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_36; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_37; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_38; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_39; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_40; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_41; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_42; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_43; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_44; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_45; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_46; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_47; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_48; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_49; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_50; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_51; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_52; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_53; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_54; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_55; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_56; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_57; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_58; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_59; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_60; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_61; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_62; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_63; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_64; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_65; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_66; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_67; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_68; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_69; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_70; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_71; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_72; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_73; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_74; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_75; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_76; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_77; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_78; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_79; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_80; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_81; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_82; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_83; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_84; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_85; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_86; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_87; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_88; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_89; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_90; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_91; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_92; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_93; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_94; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_95; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_96; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_97; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_98; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_99; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_100; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_101; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_102; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_103; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_104; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_105; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_106; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_107; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_108; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_109; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_110; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_111; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_112; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_113; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_114; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_115; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_116; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_117; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_118; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_119; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_120; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_121; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_122; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_123; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_124; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_125; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_126; // @[DenseLayer.scala 100:42]
  wire [7:0] currWeights_127; // @[DenseLayer.scala 100:42]
  wire  _T_2398; // @[DenseLayer.scala 121:33]
  wire  _T_2416; // @[DenseLayer.scala 123:16]
  wire  _GEN_264; // @[DenseLayer.scala 123:42]
  wire  _T_2418; // @[DenseLayer.scala 126:14]
  wire  _GEN_265; // @[DenseLayer.scala 126:23]
  wire [16:0] _T_2434; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2435; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2436; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_273; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_274; // @[DenseLayer.scala 135:18]
  wire  _T_2438; // @[DenseLayer.scala 138:16]
  wire [15:0] _GEN_275; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2439; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2440; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2441; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_276; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_277; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_278; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2444; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2445; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2446; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_279; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_280; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_281; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2449; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2450; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2451; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_282; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_283; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_284; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2454; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2455; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2456; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_285; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_286; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_287; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2459; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2460; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2461; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_288; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_289; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_290; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2464; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2465; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2466; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_291; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_292; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_293; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2469; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2470; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2471; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_294; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_295; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_296; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2474; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2475; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2476; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_297; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_298; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_299; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2479; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2480; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2481; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_300; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_301; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_302; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2484; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2485; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2486; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_303; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_304; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_305; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2489; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2490; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2491; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_306; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_307; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_308; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2494; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2495; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2496; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_309; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_310; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_311; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2499; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2500; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2501; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_312; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_313; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_314; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2504; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2505; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2506; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_315; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_316; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_317; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2509; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2510; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2511; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_318; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_319; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_320; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2514; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2515; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2516; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_321; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_322; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_323; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2519; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2520; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2521; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_324; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_325; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_326; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2524; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2525; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2526; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_327; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_328; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_329; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2529; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2530; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2531; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_330; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_331; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_332; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2534; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2535; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2536; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_333; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_334; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_335; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2539; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2540; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2541; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_336; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_337; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_338; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2544; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2545; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2546; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_339; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_340; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_341; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2549; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2550; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2551; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_342; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_343; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_344; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2554; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2555; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2556; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_345; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_346; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_347; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2559; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2560; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2561; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_348; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_349; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_350; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2564; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2565; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2566; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_351; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_352; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_353; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2569; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2570; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2571; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_354; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_355; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_356; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2574; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2575; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2576; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_357; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_358; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_359; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2579; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2580; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2581; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_360; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_361; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_362; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2584; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2585; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2586; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_363; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_364; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_365; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2589; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2590; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2591; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_366; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_367; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_368; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2594; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2595; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2596; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_369; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_370; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_371; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2599; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2600; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2601; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_372; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_373; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_374; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2604; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2605; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2606; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_375; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_376; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_377; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2609; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2610; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2611; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_378; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_379; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_380; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2614; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2615; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2616; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_381; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_382; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_383; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2619; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2620; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2621; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_384; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_385; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_386; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2624; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2625; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2626; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_387; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_388; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_389; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2629; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2630; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2631; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_390; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_391; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_392; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2634; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2635; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2636; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_393; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_394; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_395; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2639; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2640; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2641; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_396; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_397; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_398; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2644; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2645; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2646; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_399; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_400; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_401; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2649; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2650; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2651; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_402; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_403; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_404; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2654; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2655; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2656; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_405; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_406; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_407; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2659; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2660; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2661; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_408; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_409; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_410; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2664; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2665; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2666; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_411; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_412; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_413; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2669; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2670; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2671; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_414; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_415; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_416; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2674; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2675; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2676; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_417; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_418; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_419; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2679; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2680; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2681; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_420; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_421; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_422; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2684; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2685; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2686; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_423; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_424; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_425; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2689; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2690; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2691; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_426; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_427; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_428; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2694; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2695; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2696; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_429; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_430; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_431; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2699; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2700; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2701; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_432; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_433; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_434; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2704; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2705; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2706; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_435; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_436; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_437; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2709; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2710; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2711; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_438; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_439; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_440; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2714; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2715; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2716; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_441; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_442; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_443; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2719; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2720; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2721; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_444; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_445; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_446; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2724; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2725; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2726; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_447; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_448; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_449; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2729; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2730; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2731; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_450; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_451; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_452; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2734; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2735; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2736; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_453; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_454; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_455; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2739; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2740; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2741; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_456; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_457; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_458; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2744; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2745; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2746; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_459; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_460; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_461; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2749; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2750; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2751; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_462; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_463; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_464; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2754; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2755; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2756; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_465; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_466; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_467; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2759; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2760; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2761; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_468; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_469; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_470; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2764; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2765; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2766; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_471; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_472; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_473; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2769; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2770; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2771; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_474; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_475; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_476; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2774; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2775; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2776; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_477; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_478; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_479; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2779; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2780; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2781; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_480; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_481; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_482; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2784; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2785; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2786; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_483; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_484; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_485; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2789; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2790; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2791; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_486; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_487; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_488; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2794; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2795; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2796; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_489; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_490; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_491; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2799; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2800; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2801; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_492; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_493; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_494; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2804; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2805; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2806; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_495; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_496; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_497; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2809; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2810; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2811; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_498; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_499; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_500; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2814; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2815; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2816; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_501; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_502; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_503; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2819; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2820; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2821; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_504; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_505; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_506; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2824; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2825; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2826; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_507; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_508; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_509; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2829; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2830; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2831; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_510; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_511; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_512; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2834; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2835; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2836; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_513; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_514; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_515; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2839; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2840; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2841; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_516; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_517; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_518; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2844; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2845; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2846; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_519; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_520; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_521; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2849; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2850; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2851; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_522; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_523; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_524; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2854; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2855; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2856; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_525; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_526; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_527; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2859; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2860; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2861; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_528; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_529; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_530; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2864; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2865; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2866; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_531; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_532; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_533; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2869; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2870; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2871; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_534; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_535; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_536; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2874; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2875; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2876; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_537; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_538; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_539; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2879; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2880; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2881; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_540; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_541; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_542; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2884; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2885; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2886; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_543; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_544; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_545; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2889; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2890; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2891; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_546; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_547; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_548; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2894; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2895; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2896; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_549; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_550; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_551; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2899; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2900; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2901; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_552; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_553; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_554; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2904; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2905; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2906; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_555; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_556; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_557; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2909; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2910; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2911; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_558; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_559; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_560; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2914; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2915; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2916; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_561; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_562; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_563; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2919; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2920; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2921; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_564; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_565; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_566; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2924; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2925; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2926; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_567; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_568; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_569; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2929; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2930; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2931; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_570; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_571; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_572; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2934; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2935; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2936; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_573; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_574; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_575; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2939; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2940; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2941; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_576; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_577; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_578; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2944; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2945; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2946; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_579; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_580; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_581; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2949; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2950; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2951; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_582; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_583; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_584; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2954; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2955; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2956; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_585; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_586; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_587; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2959; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2960; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2961; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_588; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_589; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_590; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2964; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2965; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2966; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_591; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_592; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_593; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2969; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2970; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2971; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_594; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_595; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_596; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2974; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2975; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2976; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_597; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_598; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_599; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2979; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2980; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2981; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_600; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_601; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_602; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2984; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2985; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2986; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_603; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_604; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_605; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2989; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2990; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2991; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_606; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_607; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_608; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2994; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2995; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_2996; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_609; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_610; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_611; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_2999; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_3000; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_3001; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_612; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_613; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_614; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_3004; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_3005; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_3006; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_615; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_616; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_617; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_3009; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_3010; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_3011; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_618; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_619; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_620; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_3014; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_3015; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_3016; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_621; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_622; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_623; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_3019; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_3020; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_3021; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_624; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_625; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_626; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_3024; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_3025; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_3026; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_627; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_628; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_629; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_3029; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_3030; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_3031; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_630; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_631; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_632; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_3034; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_3035; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_3036; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_633; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_634; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_635; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_3039; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_3040; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_3041; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_636; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_637; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_638; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_3044; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_3045; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_3046; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_639; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_640; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_641; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_3049; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_3050; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_3051; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_642; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_643; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_644; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_3054; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_3055; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_3056; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_645; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_646; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_647; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_3059; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_3060; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_3061; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_648; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_649; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_650; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_3064; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_3065; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_3066; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_651; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_652; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_653; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_3069; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_3070; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_3071; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_654; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_655; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_656; // @[DenseLayer.scala 138:24]
  DenseBlackBox3f4b5cb0a2 weightsRAM ( // @[DenseLayer.scala 96:34]
    .out(weightsRAM_out),
    .readAddr(weightsRAM_readAddr),
    .clock(weightsRAM_clock)
  );
  FanoutAWS FanoutAWS ( // @[FanoutAWS.scala 16:26]
    .clock(FanoutAWS_clock),
    .io_in(FanoutAWS_io_in),
    .io_out_0(FanoutAWS_io_out_0),
    .io_out_1(FanoutAWS_io_out_1),
    .io_out_2(FanoutAWS_io_out_2),
    .io_out_3(FanoutAWS_io_out_3),
    .io_out_4(FanoutAWS_io_out_4),
    .io_out_5(FanoutAWS_io_out_5),
    .io_out_6(FanoutAWS_io_out_6),
    .io_out_7(FanoutAWS_io_out_7),
    .io_out_8(FanoutAWS_io_out_8),
    .io_out_9(FanoutAWS_io_out_9),
    .io_out_10(FanoutAWS_io_out_10),
    .io_out_11(FanoutAWS_io_out_11),
    .io_out_12(FanoutAWS_io_out_12),
    .io_out_13(FanoutAWS_io_out_13),
    .io_out_14(FanoutAWS_io_out_14),
    .io_out_15(FanoutAWS_io_out_15),
    .io_out_16(FanoutAWS_io_out_16),
    .io_out_17(FanoutAWS_io_out_17),
    .io_out_18(FanoutAWS_io_out_18),
    .io_out_19(FanoutAWS_io_out_19),
    .io_out_20(FanoutAWS_io_out_20),
    .io_out_21(FanoutAWS_io_out_21),
    .io_out_22(FanoutAWS_io_out_22),
    .io_out_23(FanoutAWS_io_out_23),
    .io_out_24(FanoutAWS_io_out_24),
    .io_out_25(FanoutAWS_io_out_25),
    .io_out_26(FanoutAWS_io_out_26),
    .io_out_27(FanoutAWS_io_out_27),
    .io_out_28(FanoutAWS_io_out_28),
    .io_out_29(FanoutAWS_io_out_29),
    .io_out_30(FanoutAWS_io_out_30),
    .io_out_31(FanoutAWS_io_out_31),
    .io_out_32(FanoutAWS_io_out_32),
    .io_out_33(FanoutAWS_io_out_33),
    .io_out_34(FanoutAWS_io_out_34),
    .io_out_35(FanoutAWS_io_out_35),
    .io_out_36(FanoutAWS_io_out_36),
    .io_out_37(FanoutAWS_io_out_37),
    .io_out_38(FanoutAWS_io_out_38),
    .io_out_39(FanoutAWS_io_out_39),
    .io_out_40(FanoutAWS_io_out_40),
    .io_out_41(FanoutAWS_io_out_41),
    .io_out_42(FanoutAWS_io_out_42),
    .io_out_43(FanoutAWS_io_out_43),
    .io_out_44(FanoutAWS_io_out_44),
    .io_out_45(FanoutAWS_io_out_45),
    .io_out_46(FanoutAWS_io_out_46),
    .io_out_47(FanoutAWS_io_out_47),
    .io_out_48(FanoutAWS_io_out_48),
    .io_out_49(FanoutAWS_io_out_49),
    .io_out_50(FanoutAWS_io_out_50),
    .io_out_51(FanoutAWS_io_out_51),
    .io_out_52(FanoutAWS_io_out_52),
    .io_out_53(FanoutAWS_io_out_53),
    .io_out_54(FanoutAWS_io_out_54),
    .io_out_55(FanoutAWS_io_out_55),
    .io_out_56(FanoutAWS_io_out_56),
    .io_out_57(FanoutAWS_io_out_57),
    .io_out_58(FanoutAWS_io_out_58),
    .io_out_59(FanoutAWS_io_out_59),
    .io_out_60(FanoutAWS_io_out_60),
    .io_out_61(FanoutAWS_io_out_61),
    .io_out_62(FanoutAWS_io_out_62),
    .io_out_63(FanoutAWS_io_out_63),
    .io_out_64(FanoutAWS_io_out_64),
    .io_out_65(FanoutAWS_io_out_65),
    .io_out_66(FanoutAWS_io_out_66),
    .io_out_67(FanoutAWS_io_out_67),
    .io_out_68(FanoutAWS_io_out_68),
    .io_out_69(FanoutAWS_io_out_69),
    .io_out_70(FanoutAWS_io_out_70),
    .io_out_71(FanoutAWS_io_out_71),
    .io_out_72(FanoutAWS_io_out_72),
    .io_out_73(FanoutAWS_io_out_73),
    .io_out_74(FanoutAWS_io_out_74),
    .io_out_75(FanoutAWS_io_out_75),
    .io_out_76(FanoutAWS_io_out_76),
    .io_out_77(FanoutAWS_io_out_77),
    .io_out_78(FanoutAWS_io_out_78),
    .io_out_79(FanoutAWS_io_out_79),
    .io_out_80(FanoutAWS_io_out_80),
    .io_out_81(FanoutAWS_io_out_81),
    .io_out_82(FanoutAWS_io_out_82),
    .io_out_83(FanoutAWS_io_out_83),
    .io_out_84(FanoutAWS_io_out_84),
    .io_out_85(FanoutAWS_io_out_85),
    .io_out_86(FanoutAWS_io_out_86),
    .io_out_87(FanoutAWS_io_out_87),
    .io_out_88(FanoutAWS_io_out_88),
    .io_out_89(FanoutAWS_io_out_89),
    .io_out_90(FanoutAWS_io_out_90),
    .io_out_91(FanoutAWS_io_out_91),
    .io_out_92(FanoutAWS_io_out_92),
    .io_out_93(FanoutAWS_io_out_93),
    .io_out_94(FanoutAWS_io_out_94),
    .io_out_95(FanoutAWS_io_out_95),
    .io_out_96(FanoutAWS_io_out_96),
    .io_out_97(FanoutAWS_io_out_97),
    .io_out_98(FanoutAWS_io_out_98),
    .io_out_99(FanoutAWS_io_out_99),
    .io_out_100(FanoutAWS_io_out_100),
    .io_out_101(FanoutAWS_io_out_101),
    .io_out_102(FanoutAWS_io_out_102),
    .io_out_103(FanoutAWS_io_out_103),
    .io_out_104(FanoutAWS_io_out_104),
    .io_out_105(FanoutAWS_io_out_105),
    .io_out_106(FanoutAWS_io_out_106),
    .io_out_107(FanoutAWS_io_out_107),
    .io_out_108(FanoutAWS_io_out_108),
    .io_out_109(FanoutAWS_io_out_109),
    .io_out_110(FanoutAWS_io_out_110),
    .io_out_111(FanoutAWS_io_out_111),
    .io_out_112(FanoutAWS_io_out_112),
    .io_out_113(FanoutAWS_io_out_113),
    .io_out_114(FanoutAWS_io_out_114),
    .io_out_115(FanoutAWS_io_out_115),
    .io_out_116(FanoutAWS_io_out_116),
    .io_out_117(FanoutAWS_io_out_117),
    .io_out_118(FanoutAWS_io_out_118),
    .io_out_119(FanoutAWS_io_out_119),
    .io_out_120(FanoutAWS_io_out_120),
    .io_out_121(FanoutAWS_io_out_121),
    .io_out_122(FanoutAWS_io_out_122),
    .io_out_123(FanoutAWS_io_out_123),
    .io_out_124(FanoutAWS_io_out_124),
    .io_out_125(FanoutAWS_io_out_125),
    .io_out_126(FanoutAWS_io_out_126),
    .io_out_127(FanoutAWS_io_out_127)
  );
  FanoutAWS FanoutAWS_1 ( // @[FanoutAWS.scala 16:26]
    .clock(FanoutAWS_1_clock),
    .io_in(FanoutAWS_1_io_in),
    .io_out_0(FanoutAWS_1_io_out_0),
    .io_out_1(FanoutAWS_1_io_out_1),
    .io_out_2(FanoutAWS_1_io_out_2),
    .io_out_3(FanoutAWS_1_io_out_3),
    .io_out_4(FanoutAWS_1_io_out_4),
    .io_out_5(FanoutAWS_1_io_out_5),
    .io_out_6(FanoutAWS_1_io_out_6),
    .io_out_7(FanoutAWS_1_io_out_7),
    .io_out_8(FanoutAWS_1_io_out_8),
    .io_out_9(FanoutAWS_1_io_out_9),
    .io_out_10(FanoutAWS_1_io_out_10),
    .io_out_11(FanoutAWS_1_io_out_11),
    .io_out_12(FanoutAWS_1_io_out_12),
    .io_out_13(FanoutAWS_1_io_out_13),
    .io_out_14(FanoutAWS_1_io_out_14),
    .io_out_15(FanoutAWS_1_io_out_15),
    .io_out_16(FanoutAWS_1_io_out_16),
    .io_out_17(FanoutAWS_1_io_out_17),
    .io_out_18(FanoutAWS_1_io_out_18),
    .io_out_19(FanoutAWS_1_io_out_19),
    .io_out_20(FanoutAWS_1_io_out_20),
    .io_out_21(FanoutAWS_1_io_out_21),
    .io_out_22(FanoutAWS_1_io_out_22),
    .io_out_23(FanoutAWS_1_io_out_23),
    .io_out_24(FanoutAWS_1_io_out_24),
    .io_out_25(FanoutAWS_1_io_out_25),
    .io_out_26(FanoutAWS_1_io_out_26),
    .io_out_27(FanoutAWS_1_io_out_27),
    .io_out_28(FanoutAWS_1_io_out_28),
    .io_out_29(FanoutAWS_1_io_out_29),
    .io_out_30(FanoutAWS_1_io_out_30),
    .io_out_31(FanoutAWS_1_io_out_31),
    .io_out_32(FanoutAWS_1_io_out_32),
    .io_out_33(FanoutAWS_1_io_out_33),
    .io_out_34(FanoutAWS_1_io_out_34),
    .io_out_35(FanoutAWS_1_io_out_35),
    .io_out_36(FanoutAWS_1_io_out_36),
    .io_out_37(FanoutAWS_1_io_out_37),
    .io_out_38(FanoutAWS_1_io_out_38),
    .io_out_39(FanoutAWS_1_io_out_39),
    .io_out_40(FanoutAWS_1_io_out_40),
    .io_out_41(FanoutAWS_1_io_out_41),
    .io_out_42(FanoutAWS_1_io_out_42),
    .io_out_43(FanoutAWS_1_io_out_43),
    .io_out_44(FanoutAWS_1_io_out_44),
    .io_out_45(FanoutAWS_1_io_out_45),
    .io_out_46(FanoutAWS_1_io_out_46),
    .io_out_47(FanoutAWS_1_io_out_47),
    .io_out_48(FanoutAWS_1_io_out_48),
    .io_out_49(FanoutAWS_1_io_out_49),
    .io_out_50(FanoutAWS_1_io_out_50),
    .io_out_51(FanoutAWS_1_io_out_51),
    .io_out_52(FanoutAWS_1_io_out_52),
    .io_out_53(FanoutAWS_1_io_out_53),
    .io_out_54(FanoutAWS_1_io_out_54),
    .io_out_55(FanoutAWS_1_io_out_55),
    .io_out_56(FanoutAWS_1_io_out_56),
    .io_out_57(FanoutAWS_1_io_out_57),
    .io_out_58(FanoutAWS_1_io_out_58),
    .io_out_59(FanoutAWS_1_io_out_59),
    .io_out_60(FanoutAWS_1_io_out_60),
    .io_out_61(FanoutAWS_1_io_out_61),
    .io_out_62(FanoutAWS_1_io_out_62),
    .io_out_63(FanoutAWS_1_io_out_63),
    .io_out_64(FanoutAWS_1_io_out_64),
    .io_out_65(FanoutAWS_1_io_out_65),
    .io_out_66(FanoutAWS_1_io_out_66),
    .io_out_67(FanoutAWS_1_io_out_67),
    .io_out_68(FanoutAWS_1_io_out_68),
    .io_out_69(FanoutAWS_1_io_out_69),
    .io_out_70(FanoutAWS_1_io_out_70),
    .io_out_71(FanoutAWS_1_io_out_71),
    .io_out_72(FanoutAWS_1_io_out_72),
    .io_out_73(FanoutAWS_1_io_out_73),
    .io_out_74(FanoutAWS_1_io_out_74),
    .io_out_75(FanoutAWS_1_io_out_75),
    .io_out_76(FanoutAWS_1_io_out_76),
    .io_out_77(FanoutAWS_1_io_out_77),
    .io_out_78(FanoutAWS_1_io_out_78),
    .io_out_79(FanoutAWS_1_io_out_79),
    .io_out_80(FanoutAWS_1_io_out_80),
    .io_out_81(FanoutAWS_1_io_out_81),
    .io_out_82(FanoutAWS_1_io_out_82),
    .io_out_83(FanoutAWS_1_io_out_83),
    .io_out_84(FanoutAWS_1_io_out_84),
    .io_out_85(FanoutAWS_1_io_out_85),
    .io_out_86(FanoutAWS_1_io_out_86),
    .io_out_87(FanoutAWS_1_io_out_87),
    .io_out_88(FanoutAWS_1_io_out_88),
    .io_out_89(FanoutAWS_1_io_out_89),
    .io_out_90(FanoutAWS_1_io_out_90),
    .io_out_91(FanoutAWS_1_io_out_91),
    .io_out_92(FanoutAWS_1_io_out_92),
    .io_out_93(FanoutAWS_1_io_out_93),
    .io_out_94(FanoutAWS_1_io_out_94),
    .io_out_95(FanoutAWS_1_io_out_95),
    .io_out_96(FanoutAWS_1_io_out_96),
    .io_out_97(FanoutAWS_1_io_out_97),
    .io_out_98(FanoutAWS_1_io_out_98),
    .io_out_99(FanoutAWS_1_io_out_99),
    .io_out_100(FanoutAWS_1_io_out_100),
    .io_out_101(FanoutAWS_1_io_out_101),
    .io_out_102(FanoutAWS_1_io_out_102),
    .io_out_103(FanoutAWS_1_io_out_103),
    .io_out_104(FanoutAWS_1_io_out_104),
    .io_out_105(FanoutAWS_1_io_out_105),
    .io_out_106(FanoutAWS_1_io_out_106),
    .io_out_107(FanoutAWS_1_io_out_107),
    .io_out_108(FanoutAWS_1_io_out_108),
    .io_out_109(FanoutAWS_1_io_out_109),
    .io_out_110(FanoutAWS_1_io_out_110),
    .io_out_111(FanoutAWS_1_io_out_111),
    .io_out_112(FanoutAWS_1_io_out_112),
    .io_out_113(FanoutAWS_1_io_out_113),
    .io_out_114(FanoutAWS_1_io_out_114),
    .io_out_115(FanoutAWS_1_io_out_115),
    .io_out_116(FanoutAWS_1_io_out_116),
    .io_out_117(FanoutAWS_1_io_out_117),
    .io_out_118(FanoutAWS_1_io_out_118),
    .io_out_119(FanoutAWS_1_io_out_119),
    .io_out_120(FanoutAWS_1_io_out_120),
    .io_out_121(FanoutAWS_1_io_out_121),
    .io_out_122(FanoutAWS_1_io_out_122),
    .io_out_123(FanoutAWS_1_io_out_123),
    .io_out_124(FanoutAWS_1_io_out_124),
    .io_out_125(FanoutAWS_1_io_out_125),
    .io_out_126(FanoutAWS_1_io_out_126),
    .io_out_127(FanoutAWS_1_io_out_127)
  );
  FanoutAWS FanoutAWS_2 ( // @[FanoutAWS.scala 16:26]
    .clock(FanoutAWS_2_clock),
    .io_in(FanoutAWS_2_io_in),
    .io_out_0(FanoutAWS_2_io_out_0),
    .io_out_1(FanoutAWS_2_io_out_1),
    .io_out_2(FanoutAWS_2_io_out_2),
    .io_out_3(FanoutAWS_2_io_out_3),
    .io_out_4(FanoutAWS_2_io_out_4),
    .io_out_5(FanoutAWS_2_io_out_5),
    .io_out_6(FanoutAWS_2_io_out_6),
    .io_out_7(FanoutAWS_2_io_out_7),
    .io_out_8(FanoutAWS_2_io_out_8),
    .io_out_9(FanoutAWS_2_io_out_9),
    .io_out_10(FanoutAWS_2_io_out_10),
    .io_out_11(FanoutAWS_2_io_out_11),
    .io_out_12(FanoutAWS_2_io_out_12),
    .io_out_13(FanoutAWS_2_io_out_13),
    .io_out_14(FanoutAWS_2_io_out_14),
    .io_out_15(FanoutAWS_2_io_out_15),
    .io_out_16(FanoutAWS_2_io_out_16),
    .io_out_17(FanoutAWS_2_io_out_17),
    .io_out_18(FanoutAWS_2_io_out_18),
    .io_out_19(FanoutAWS_2_io_out_19),
    .io_out_20(FanoutAWS_2_io_out_20),
    .io_out_21(FanoutAWS_2_io_out_21),
    .io_out_22(FanoutAWS_2_io_out_22),
    .io_out_23(FanoutAWS_2_io_out_23),
    .io_out_24(FanoutAWS_2_io_out_24),
    .io_out_25(FanoutAWS_2_io_out_25),
    .io_out_26(FanoutAWS_2_io_out_26),
    .io_out_27(FanoutAWS_2_io_out_27),
    .io_out_28(FanoutAWS_2_io_out_28),
    .io_out_29(FanoutAWS_2_io_out_29),
    .io_out_30(FanoutAWS_2_io_out_30),
    .io_out_31(FanoutAWS_2_io_out_31),
    .io_out_32(FanoutAWS_2_io_out_32),
    .io_out_33(FanoutAWS_2_io_out_33),
    .io_out_34(FanoutAWS_2_io_out_34),
    .io_out_35(FanoutAWS_2_io_out_35),
    .io_out_36(FanoutAWS_2_io_out_36),
    .io_out_37(FanoutAWS_2_io_out_37),
    .io_out_38(FanoutAWS_2_io_out_38),
    .io_out_39(FanoutAWS_2_io_out_39),
    .io_out_40(FanoutAWS_2_io_out_40),
    .io_out_41(FanoutAWS_2_io_out_41),
    .io_out_42(FanoutAWS_2_io_out_42),
    .io_out_43(FanoutAWS_2_io_out_43),
    .io_out_44(FanoutAWS_2_io_out_44),
    .io_out_45(FanoutAWS_2_io_out_45),
    .io_out_46(FanoutAWS_2_io_out_46),
    .io_out_47(FanoutAWS_2_io_out_47),
    .io_out_48(FanoutAWS_2_io_out_48),
    .io_out_49(FanoutAWS_2_io_out_49),
    .io_out_50(FanoutAWS_2_io_out_50),
    .io_out_51(FanoutAWS_2_io_out_51),
    .io_out_52(FanoutAWS_2_io_out_52),
    .io_out_53(FanoutAWS_2_io_out_53),
    .io_out_54(FanoutAWS_2_io_out_54),
    .io_out_55(FanoutAWS_2_io_out_55),
    .io_out_56(FanoutAWS_2_io_out_56),
    .io_out_57(FanoutAWS_2_io_out_57),
    .io_out_58(FanoutAWS_2_io_out_58),
    .io_out_59(FanoutAWS_2_io_out_59),
    .io_out_60(FanoutAWS_2_io_out_60),
    .io_out_61(FanoutAWS_2_io_out_61),
    .io_out_62(FanoutAWS_2_io_out_62),
    .io_out_63(FanoutAWS_2_io_out_63),
    .io_out_64(FanoutAWS_2_io_out_64),
    .io_out_65(FanoutAWS_2_io_out_65),
    .io_out_66(FanoutAWS_2_io_out_66),
    .io_out_67(FanoutAWS_2_io_out_67),
    .io_out_68(FanoutAWS_2_io_out_68),
    .io_out_69(FanoutAWS_2_io_out_69),
    .io_out_70(FanoutAWS_2_io_out_70),
    .io_out_71(FanoutAWS_2_io_out_71),
    .io_out_72(FanoutAWS_2_io_out_72),
    .io_out_73(FanoutAWS_2_io_out_73),
    .io_out_74(FanoutAWS_2_io_out_74),
    .io_out_75(FanoutAWS_2_io_out_75),
    .io_out_76(FanoutAWS_2_io_out_76),
    .io_out_77(FanoutAWS_2_io_out_77),
    .io_out_78(FanoutAWS_2_io_out_78),
    .io_out_79(FanoutAWS_2_io_out_79),
    .io_out_80(FanoutAWS_2_io_out_80),
    .io_out_81(FanoutAWS_2_io_out_81),
    .io_out_82(FanoutAWS_2_io_out_82),
    .io_out_83(FanoutAWS_2_io_out_83),
    .io_out_84(FanoutAWS_2_io_out_84),
    .io_out_85(FanoutAWS_2_io_out_85),
    .io_out_86(FanoutAWS_2_io_out_86),
    .io_out_87(FanoutAWS_2_io_out_87),
    .io_out_88(FanoutAWS_2_io_out_88),
    .io_out_89(FanoutAWS_2_io_out_89),
    .io_out_90(FanoutAWS_2_io_out_90),
    .io_out_91(FanoutAWS_2_io_out_91),
    .io_out_92(FanoutAWS_2_io_out_92),
    .io_out_93(FanoutAWS_2_io_out_93),
    .io_out_94(FanoutAWS_2_io_out_94),
    .io_out_95(FanoutAWS_2_io_out_95),
    .io_out_96(FanoutAWS_2_io_out_96),
    .io_out_97(FanoutAWS_2_io_out_97),
    .io_out_98(FanoutAWS_2_io_out_98),
    .io_out_99(FanoutAWS_2_io_out_99),
    .io_out_100(FanoutAWS_2_io_out_100),
    .io_out_101(FanoutAWS_2_io_out_101),
    .io_out_102(FanoutAWS_2_io_out_102),
    .io_out_103(FanoutAWS_2_io_out_103),
    .io_out_104(FanoutAWS_2_io_out_104),
    .io_out_105(FanoutAWS_2_io_out_105),
    .io_out_106(FanoutAWS_2_io_out_106),
    .io_out_107(FanoutAWS_2_io_out_107),
    .io_out_108(FanoutAWS_2_io_out_108),
    .io_out_109(FanoutAWS_2_io_out_109),
    .io_out_110(FanoutAWS_2_io_out_110),
    .io_out_111(FanoutAWS_2_io_out_111),
    .io_out_112(FanoutAWS_2_io_out_112),
    .io_out_113(FanoutAWS_2_io_out_113),
    .io_out_114(FanoutAWS_2_io_out_114),
    .io_out_115(FanoutAWS_2_io_out_115),
    .io_out_116(FanoutAWS_2_io_out_116),
    .io_out_117(FanoutAWS_2_io_out_117),
    .io_out_118(FanoutAWS_2_io_out_118),
    .io_out_119(FanoutAWS_2_io_out_119),
    .io_out_120(FanoutAWS_2_io_out_120),
    .io_out_121(FanoutAWS_2_io_out_121),
    .io_out_122(FanoutAWS_2_io_out_122),
    .io_out_123(FanoutAWS_2_io_out_123),
    .io_out_124(FanoutAWS_2_io_out_124),
    .io_out_125(FanoutAWS_2_io_out_125),
    .io_out_126(FanoutAWS_2_io_out_126),
    .io_out_127(FanoutAWS_2_io_out_127)
  );
  FanoutAWS FanoutAWS_3 ( // @[FanoutAWS.scala 16:26]
    .clock(FanoutAWS_3_clock),
    .io_in(FanoutAWS_3_io_in),
    .io_out_0(FanoutAWS_3_io_out_0),
    .io_out_1(FanoutAWS_3_io_out_1),
    .io_out_2(FanoutAWS_3_io_out_2),
    .io_out_3(FanoutAWS_3_io_out_3),
    .io_out_4(FanoutAWS_3_io_out_4),
    .io_out_5(FanoutAWS_3_io_out_5),
    .io_out_6(FanoutAWS_3_io_out_6),
    .io_out_7(FanoutAWS_3_io_out_7),
    .io_out_8(FanoutAWS_3_io_out_8),
    .io_out_9(FanoutAWS_3_io_out_9),
    .io_out_10(FanoutAWS_3_io_out_10),
    .io_out_11(FanoutAWS_3_io_out_11),
    .io_out_12(FanoutAWS_3_io_out_12),
    .io_out_13(FanoutAWS_3_io_out_13),
    .io_out_14(FanoutAWS_3_io_out_14),
    .io_out_15(FanoutAWS_3_io_out_15),
    .io_out_16(FanoutAWS_3_io_out_16),
    .io_out_17(FanoutAWS_3_io_out_17),
    .io_out_18(FanoutAWS_3_io_out_18),
    .io_out_19(FanoutAWS_3_io_out_19),
    .io_out_20(FanoutAWS_3_io_out_20),
    .io_out_21(FanoutAWS_3_io_out_21),
    .io_out_22(FanoutAWS_3_io_out_22),
    .io_out_23(FanoutAWS_3_io_out_23),
    .io_out_24(FanoutAWS_3_io_out_24),
    .io_out_25(FanoutAWS_3_io_out_25),
    .io_out_26(FanoutAWS_3_io_out_26),
    .io_out_27(FanoutAWS_3_io_out_27),
    .io_out_28(FanoutAWS_3_io_out_28),
    .io_out_29(FanoutAWS_3_io_out_29),
    .io_out_30(FanoutAWS_3_io_out_30),
    .io_out_31(FanoutAWS_3_io_out_31),
    .io_out_32(FanoutAWS_3_io_out_32),
    .io_out_33(FanoutAWS_3_io_out_33),
    .io_out_34(FanoutAWS_3_io_out_34),
    .io_out_35(FanoutAWS_3_io_out_35),
    .io_out_36(FanoutAWS_3_io_out_36),
    .io_out_37(FanoutAWS_3_io_out_37),
    .io_out_38(FanoutAWS_3_io_out_38),
    .io_out_39(FanoutAWS_3_io_out_39),
    .io_out_40(FanoutAWS_3_io_out_40),
    .io_out_41(FanoutAWS_3_io_out_41),
    .io_out_42(FanoutAWS_3_io_out_42),
    .io_out_43(FanoutAWS_3_io_out_43),
    .io_out_44(FanoutAWS_3_io_out_44),
    .io_out_45(FanoutAWS_3_io_out_45),
    .io_out_46(FanoutAWS_3_io_out_46),
    .io_out_47(FanoutAWS_3_io_out_47),
    .io_out_48(FanoutAWS_3_io_out_48),
    .io_out_49(FanoutAWS_3_io_out_49),
    .io_out_50(FanoutAWS_3_io_out_50),
    .io_out_51(FanoutAWS_3_io_out_51),
    .io_out_52(FanoutAWS_3_io_out_52),
    .io_out_53(FanoutAWS_3_io_out_53),
    .io_out_54(FanoutAWS_3_io_out_54),
    .io_out_55(FanoutAWS_3_io_out_55),
    .io_out_56(FanoutAWS_3_io_out_56),
    .io_out_57(FanoutAWS_3_io_out_57),
    .io_out_58(FanoutAWS_3_io_out_58),
    .io_out_59(FanoutAWS_3_io_out_59),
    .io_out_60(FanoutAWS_3_io_out_60),
    .io_out_61(FanoutAWS_3_io_out_61),
    .io_out_62(FanoutAWS_3_io_out_62),
    .io_out_63(FanoutAWS_3_io_out_63),
    .io_out_64(FanoutAWS_3_io_out_64),
    .io_out_65(FanoutAWS_3_io_out_65),
    .io_out_66(FanoutAWS_3_io_out_66),
    .io_out_67(FanoutAWS_3_io_out_67),
    .io_out_68(FanoutAWS_3_io_out_68),
    .io_out_69(FanoutAWS_3_io_out_69),
    .io_out_70(FanoutAWS_3_io_out_70),
    .io_out_71(FanoutAWS_3_io_out_71),
    .io_out_72(FanoutAWS_3_io_out_72),
    .io_out_73(FanoutAWS_3_io_out_73),
    .io_out_74(FanoutAWS_3_io_out_74),
    .io_out_75(FanoutAWS_3_io_out_75),
    .io_out_76(FanoutAWS_3_io_out_76),
    .io_out_77(FanoutAWS_3_io_out_77),
    .io_out_78(FanoutAWS_3_io_out_78),
    .io_out_79(FanoutAWS_3_io_out_79),
    .io_out_80(FanoutAWS_3_io_out_80),
    .io_out_81(FanoutAWS_3_io_out_81),
    .io_out_82(FanoutAWS_3_io_out_82),
    .io_out_83(FanoutAWS_3_io_out_83),
    .io_out_84(FanoutAWS_3_io_out_84),
    .io_out_85(FanoutAWS_3_io_out_85),
    .io_out_86(FanoutAWS_3_io_out_86),
    .io_out_87(FanoutAWS_3_io_out_87),
    .io_out_88(FanoutAWS_3_io_out_88),
    .io_out_89(FanoutAWS_3_io_out_89),
    .io_out_90(FanoutAWS_3_io_out_90),
    .io_out_91(FanoutAWS_3_io_out_91),
    .io_out_92(FanoutAWS_3_io_out_92),
    .io_out_93(FanoutAWS_3_io_out_93),
    .io_out_94(FanoutAWS_3_io_out_94),
    .io_out_95(FanoutAWS_3_io_out_95),
    .io_out_96(FanoutAWS_3_io_out_96),
    .io_out_97(FanoutAWS_3_io_out_97),
    .io_out_98(FanoutAWS_3_io_out_98),
    .io_out_99(FanoutAWS_3_io_out_99),
    .io_out_100(FanoutAWS_3_io_out_100),
    .io_out_101(FanoutAWS_3_io_out_101),
    .io_out_102(FanoutAWS_3_io_out_102),
    .io_out_103(FanoutAWS_3_io_out_103),
    .io_out_104(FanoutAWS_3_io_out_104),
    .io_out_105(FanoutAWS_3_io_out_105),
    .io_out_106(FanoutAWS_3_io_out_106),
    .io_out_107(FanoutAWS_3_io_out_107),
    .io_out_108(FanoutAWS_3_io_out_108),
    .io_out_109(FanoutAWS_3_io_out_109),
    .io_out_110(FanoutAWS_3_io_out_110),
    .io_out_111(FanoutAWS_3_io_out_111),
    .io_out_112(FanoutAWS_3_io_out_112),
    .io_out_113(FanoutAWS_3_io_out_113),
    .io_out_114(FanoutAWS_3_io_out_114),
    .io_out_115(FanoutAWS_3_io_out_115),
    .io_out_116(FanoutAWS_3_io_out_116),
    .io_out_117(FanoutAWS_3_io_out_117),
    .io_out_118(FanoutAWS_3_io_out_118),
    .io_out_119(FanoutAWS_3_io_out_119),
    .io_out_120(FanoutAWS_3_io_out_120),
    .io_out_121(FanoutAWS_3_io_out_121),
    .io_out_122(FanoutAWS_3_io_out_122),
    .io_out_123(FanoutAWS_3_io_out_123),
    .io_out_124(FanoutAWS_3_io_out_124),
    .io_out_125(FanoutAWS_3_io_out_125),
    .io_out_126(FanoutAWS_3_io_out_126),
    .io_out_127(FanoutAWS_3_io_out_127)
  );
  MultiplyAccumulate MultiplyAccumulate ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_clock),
    .io_activations_0(MultiplyAccumulate_io_activations_0),
    .io_activations_1(MultiplyAccumulate_io_activations_1),
    .io_activations_2(MultiplyAccumulate_io_activations_2),
    .io_activations_3(MultiplyAccumulate_io_activations_3),
    .io_weights(MultiplyAccumulate_io_weights),
    .io_sum(MultiplyAccumulate_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_1 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_1_clock),
    .io_activations_0(MultiplyAccumulate_1_io_activations_0),
    .io_activations_1(MultiplyAccumulate_1_io_activations_1),
    .io_activations_2(MultiplyAccumulate_1_io_activations_2),
    .io_activations_3(MultiplyAccumulate_1_io_activations_3),
    .io_weights(MultiplyAccumulate_1_io_weights),
    .io_sum(MultiplyAccumulate_1_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_2 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_2_clock),
    .io_activations_0(MultiplyAccumulate_2_io_activations_0),
    .io_activations_1(MultiplyAccumulate_2_io_activations_1),
    .io_activations_2(MultiplyAccumulate_2_io_activations_2),
    .io_activations_3(MultiplyAccumulate_2_io_activations_3),
    .io_weights(MultiplyAccumulate_2_io_weights),
    .io_sum(MultiplyAccumulate_2_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_3 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_3_clock),
    .io_activations_0(MultiplyAccumulate_3_io_activations_0),
    .io_activations_1(MultiplyAccumulate_3_io_activations_1),
    .io_activations_2(MultiplyAccumulate_3_io_activations_2),
    .io_activations_3(MultiplyAccumulate_3_io_activations_3),
    .io_weights(MultiplyAccumulate_3_io_weights),
    .io_sum(MultiplyAccumulate_3_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_4 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_4_clock),
    .io_activations_0(MultiplyAccumulate_4_io_activations_0),
    .io_activations_1(MultiplyAccumulate_4_io_activations_1),
    .io_activations_2(MultiplyAccumulate_4_io_activations_2),
    .io_activations_3(MultiplyAccumulate_4_io_activations_3),
    .io_weights(MultiplyAccumulate_4_io_weights),
    .io_sum(MultiplyAccumulate_4_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_5 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_5_clock),
    .io_activations_0(MultiplyAccumulate_5_io_activations_0),
    .io_activations_1(MultiplyAccumulate_5_io_activations_1),
    .io_activations_2(MultiplyAccumulate_5_io_activations_2),
    .io_activations_3(MultiplyAccumulate_5_io_activations_3),
    .io_weights(MultiplyAccumulate_5_io_weights),
    .io_sum(MultiplyAccumulate_5_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_6 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_6_clock),
    .io_activations_0(MultiplyAccumulate_6_io_activations_0),
    .io_activations_1(MultiplyAccumulate_6_io_activations_1),
    .io_activations_2(MultiplyAccumulate_6_io_activations_2),
    .io_activations_3(MultiplyAccumulate_6_io_activations_3),
    .io_weights(MultiplyAccumulate_6_io_weights),
    .io_sum(MultiplyAccumulate_6_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_7 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_7_clock),
    .io_activations_0(MultiplyAccumulate_7_io_activations_0),
    .io_activations_1(MultiplyAccumulate_7_io_activations_1),
    .io_activations_2(MultiplyAccumulate_7_io_activations_2),
    .io_activations_3(MultiplyAccumulate_7_io_activations_3),
    .io_weights(MultiplyAccumulate_7_io_weights),
    .io_sum(MultiplyAccumulate_7_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_8 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_8_clock),
    .io_activations_0(MultiplyAccumulate_8_io_activations_0),
    .io_activations_1(MultiplyAccumulate_8_io_activations_1),
    .io_activations_2(MultiplyAccumulate_8_io_activations_2),
    .io_activations_3(MultiplyAccumulate_8_io_activations_3),
    .io_weights(MultiplyAccumulate_8_io_weights),
    .io_sum(MultiplyAccumulate_8_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_9 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_9_clock),
    .io_activations_0(MultiplyAccumulate_9_io_activations_0),
    .io_activations_1(MultiplyAccumulate_9_io_activations_1),
    .io_activations_2(MultiplyAccumulate_9_io_activations_2),
    .io_activations_3(MultiplyAccumulate_9_io_activations_3),
    .io_weights(MultiplyAccumulate_9_io_weights),
    .io_sum(MultiplyAccumulate_9_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_10 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_10_clock),
    .io_activations_0(MultiplyAccumulate_10_io_activations_0),
    .io_activations_1(MultiplyAccumulate_10_io_activations_1),
    .io_activations_2(MultiplyAccumulate_10_io_activations_2),
    .io_activations_3(MultiplyAccumulate_10_io_activations_3),
    .io_weights(MultiplyAccumulate_10_io_weights),
    .io_sum(MultiplyAccumulate_10_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_11 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_11_clock),
    .io_activations_0(MultiplyAccumulate_11_io_activations_0),
    .io_activations_1(MultiplyAccumulate_11_io_activations_1),
    .io_activations_2(MultiplyAccumulate_11_io_activations_2),
    .io_activations_3(MultiplyAccumulate_11_io_activations_3),
    .io_weights(MultiplyAccumulate_11_io_weights),
    .io_sum(MultiplyAccumulate_11_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_12 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_12_clock),
    .io_activations_0(MultiplyAccumulate_12_io_activations_0),
    .io_activations_1(MultiplyAccumulate_12_io_activations_1),
    .io_activations_2(MultiplyAccumulate_12_io_activations_2),
    .io_activations_3(MultiplyAccumulate_12_io_activations_3),
    .io_weights(MultiplyAccumulate_12_io_weights),
    .io_sum(MultiplyAccumulate_12_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_13 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_13_clock),
    .io_activations_0(MultiplyAccumulate_13_io_activations_0),
    .io_activations_1(MultiplyAccumulate_13_io_activations_1),
    .io_activations_2(MultiplyAccumulate_13_io_activations_2),
    .io_activations_3(MultiplyAccumulate_13_io_activations_3),
    .io_weights(MultiplyAccumulate_13_io_weights),
    .io_sum(MultiplyAccumulate_13_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_14 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_14_clock),
    .io_activations_0(MultiplyAccumulate_14_io_activations_0),
    .io_activations_1(MultiplyAccumulate_14_io_activations_1),
    .io_activations_2(MultiplyAccumulate_14_io_activations_2),
    .io_activations_3(MultiplyAccumulate_14_io_activations_3),
    .io_weights(MultiplyAccumulate_14_io_weights),
    .io_sum(MultiplyAccumulate_14_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_15 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_15_clock),
    .io_activations_0(MultiplyAccumulate_15_io_activations_0),
    .io_activations_1(MultiplyAccumulate_15_io_activations_1),
    .io_activations_2(MultiplyAccumulate_15_io_activations_2),
    .io_activations_3(MultiplyAccumulate_15_io_activations_3),
    .io_weights(MultiplyAccumulate_15_io_weights),
    .io_sum(MultiplyAccumulate_15_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_16 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_16_clock),
    .io_activations_0(MultiplyAccumulate_16_io_activations_0),
    .io_activations_1(MultiplyAccumulate_16_io_activations_1),
    .io_activations_2(MultiplyAccumulate_16_io_activations_2),
    .io_activations_3(MultiplyAccumulate_16_io_activations_3),
    .io_weights(MultiplyAccumulate_16_io_weights),
    .io_sum(MultiplyAccumulate_16_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_17 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_17_clock),
    .io_activations_0(MultiplyAccumulate_17_io_activations_0),
    .io_activations_1(MultiplyAccumulate_17_io_activations_1),
    .io_activations_2(MultiplyAccumulate_17_io_activations_2),
    .io_activations_3(MultiplyAccumulate_17_io_activations_3),
    .io_weights(MultiplyAccumulate_17_io_weights),
    .io_sum(MultiplyAccumulate_17_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_18 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_18_clock),
    .io_activations_0(MultiplyAccumulate_18_io_activations_0),
    .io_activations_1(MultiplyAccumulate_18_io_activations_1),
    .io_activations_2(MultiplyAccumulate_18_io_activations_2),
    .io_activations_3(MultiplyAccumulate_18_io_activations_3),
    .io_weights(MultiplyAccumulate_18_io_weights),
    .io_sum(MultiplyAccumulate_18_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_19 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_19_clock),
    .io_activations_0(MultiplyAccumulate_19_io_activations_0),
    .io_activations_1(MultiplyAccumulate_19_io_activations_1),
    .io_activations_2(MultiplyAccumulate_19_io_activations_2),
    .io_activations_3(MultiplyAccumulate_19_io_activations_3),
    .io_weights(MultiplyAccumulate_19_io_weights),
    .io_sum(MultiplyAccumulate_19_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_20 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_20_clock),
    .io_activations_0(MultiplyAccumulate_20_io_activations_0),
    .io_activations_1(MultiplyAccumulate_20_io_activations_1),
    .io_activations_2(MultiplyAccumulate_20_io_activations_2),
    .io_activations_3(MultiplyAccumulate_20_io_activations_3),
    .io_weights(MultiplyAccumulate_20_io_weights),
    .io_sum(MultiplyAccumulate_20_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_21 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_21_clock),
    .io_activations_0(MultiplyAccumulate_21_io_activations_0),
    .io_activations_1(MultiplyAccumulate_21_io_activations_1),
    .io_activations_2(MultiplyAccumulate_21_io_activations_2),
    .io_activations_3(MultiplyAccumulate_21_io_activations_3),
    .io_weights(MultiplyAccumulate_21_io_weights),
    .io_sum(MultiplyAccumulate_21_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_22 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_22_clock),
    .io_activations_0(MultiplyAccumulate_22_io_activations_0),
    .io_activations_1(MultiplyAccumulate_22_io_activations_1),
    .io_activations_2(MultiplyAccumulate_22_io_activations_2),
    .io_activations_3(MultiplyAccumulate_22_io_activations_3),
    .io_weights(MultiplyAccumulate_22_io_weights),
    .io_sum(MultiplyAccumulate_22_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_23 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_23_clock),
    .io_activations_0(MultiplyAccumulate_23_io_activations_0),
    .io_activations_1(MultiplyAccumulate_23_io_activations_1),
    .io_activations_2(MultiplyAccumulate_23_io_activations_2),
    .io_activations_3(MultiplyAccumulate_23_io_activations_3),
    .io_weights(MultiplyAccumulate_23_io_weights),
    .io_sum(MultiplyAccumulate_23_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_24 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_24_clock),
    .io_activations_0(MultiplyAccumulate_24_io_activations_0),
    .io_activations_1(MultiplyAccumulate_24_io_activations_1),
    .io_activations_2(MultiplyAccumulate_24_io_activations_2),
    .io_activations_3(MultiplyAccumulate_24_io_activations_3),
    .io_weights(MultiplyAccumulate_24_io_weights),
    .io_sum(MultiplyAccumulate_24_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_25 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_25_clock),
    .io_activations_0(MultiplyAccumulate_25_io_activations_0),
    .io_activations_1(MultiplyAccumulate_25_io_activations_1),
    .io_activations_2(MultiplyAccumulate_25_io_activations_2),
    .io_activations_3(MultiplyAccumulate_25_io_activations_3),
    .io_weights(MultiplyAccumulate_25_io_weights),
    .io_sum(MultiplyAccumulate_25_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_26 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_26_clock),
    .io_activations_0(MultiplyAccumulate_26_io_activations_0),
    .io_activations_1(MultiplyAccumulate_26_io_activations_1),
    .io_activations_2(MultiplyAccumulate_26_io_activations_2),
    .io_activations_3(MultiplyAccumulate_26_io_activations_3),
    .io_weights(MultiplyAccumulate_26_io_weights),
    .io_sum(MultiplyAccumulate_26_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_27 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_27_clock),
    .io_activations_0(MultiplyAccumulate_27_io_activations_0),
    .io_activations_1(MultiplyAccumulate_27_io_activations_1),
    .io_activations_2(MultiplyAccumulate_27_io_activations_2),
    .io_activations_3(MultiplyAccumulate_27_io_activations_3),
    .io_weights(MultiplyAccumulate_27_io_weights),
    .io_sum(MultiplyAccumulate_27_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_28 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_28_clock),
    .io_activations_0(MultiplyAccumulate_28_io_activations_0),
    .io_activations_1(MultiplyAccumulate_28_io_activations_1),
    .io_activations_2(MultiplyAccumulate_28_io_activations_2),
    .io_activations_3(MultiplyAccumulate_28_io_activations_3),
    .io_weights(MultiplyAccumulate_28_io_weights),
    .io_sum(MultiplyAccumulate_28_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_29 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_29_clock),
    .io_activations_0(MultiplyAccumulate_29_io_activations_0),
    .io_activations_1(MultiplyAccumulate_29_io_activations_1),
    .io_activations_2(MultiplyAccumulate_29_io_activations_2),
    .io_activations_3(MultiplyAccumulate_29_io_activations_3),
    .io_weights(MultiplyAccumulate_29_io_weights),
    .io_sum(MultiplyAccumulate_29_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_30 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_30_clock),
    .io_activations_0(MultiplyAccumulate_30_io_activations_0),
    .io_activations_1(MultiplyAccumulate_30_io_activations_1),
    .io_activations_2(MultiplyAccumulate_30_io_activations_2),
    .io_activations_3(MultiplyAccumulate_30_io_activations_3),
    .io_weights(MultiplyAccumulate_30_io_weights),
    .io_sum(MultiplyAccumulate_30_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_31 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_31_clock),
    .io_activations_0(MultiplyAccumulate_31_io_activations_0),
    .io_activations_1(MultiplyAccumulate_31_io_activations_1),
    .io_activations_2(MultiplyAccumulate_31_io_activations_2),
    .io_activations_3(MultiplyAccumulate_31_io_activations_3),
    .io_weights(MultiplyAccumulate_31_io_weights),
    .io_sum(MultiplyAccumulate_31_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_32 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_32_clock),
    .io_activations_0(MultiplyAccumulate_32_io_activations_0),
    .io_activations_1(MultiplyAccumulate_32_io_activations_1),
    .io_activations_2(MultiplyAccumulate_32_io_activations_2),
    .io_activations_3(MultiplyAccumulate_32_io_activations_3),
    .io_weights(MultiplyAccumulate_32_io_weights),
    .io_sum(MultiplyAccumulate_32_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_33 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_33_clock),
    .io_activations_0(MultiplyAccumulate_33_io_activations_0),
    .io_activations_1(MultiplyAccumulate_33_io_activations_1),
    .io_activations_2(MultiplyAccumulate_33_io_activations_2),
    .io_activations_3(MultiplyAccumulate_33_io_activations_3),
    .io_weights(MultiplyAccumulate_33_io_weights),
    .io_sum(MultiplyAccumulate_33_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_34 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_34_clock),
    .io_activations_0(MultiplyAccumulate_34_io_activations_0),
    .io_activations_1(MultiplyAccumulate_34_io_activations_1),
    .io_activations_2(MultiplyAccumulate_34_io_activations_2),
    .io_activations_3(MultiplyAccumulate_34_io_activations_3),
    .io_weights(MultiplyAccumulate_34_io_weights),
    .io_sum(MultiplyAccumulate_34_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_35 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_35_clock),
    .io_activations_0(MultiplyAccumulate_35_io_activations_0),
    .io_activations_1(MultiplyAccumulate_35_io_activations_1),
    .io_activations_2(MultiplyAccumulate_35_io_activations_2),
    .io_activations_3(MultiplyAccumulate_35_io_activations_3),
    .io_weights(MultiplyAccumulate_35_io_weights),
    .io_sum(MultiplyAccumulate_35_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_36 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_36_clock),
    .io_activations_0(MultiplyAccumulate_36_io_activations_0),
    .io_activations_1(MultiplyAccumulate_36_io_activations_1),
    .io_activations_2(MultiplyAccumulate_36_io_activations_2),
    .io_activations_3(MultiplyAccumulate_36_io_activations_3),
    .io_weights(MultiplyAccumulate_36_io_weights),
    .io_sum(MultiplyAccumulate_36_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_37 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_37_clock),
    .io_activations_0(MultiplyAccumulate_37_io_activations_0),
    .io_activations_1(MultiplyAccumulate_37_io_activations_1),
    .io_activations_2(MultiplyAccumulate_37_io_activations_2),
    .io_activations_3(MultiplyAccumulate_37_io_activations_3),
    .io_weights(MultiplyAccumulate_37_io_weights),
    .io_sum(MultiplyAccumulate_37_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_38 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_38_clock),
    .io_activations_0(MultiplyAccumulate_38_io_activations_0),
    .io_activations_1(MultiplyAccumulate_38_io_activations_1),
    .io_activations_2(MultiplyAccumulate_38_io_activations_2),
    .io_activations_3(MultiplyAccumulate_38_io_activations_3),
    .io_weights(MultiplyAccumulate_38_io_weights),
    .io_sum(MultiplyAccumulate_38_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_39 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_39_clock),
    .io_activations_0(MultiplyAccumulate_39_io_activations_0),
    .io_activations_1(MultiplyAccumulate_39_io_activations_1),
    .io_activations_2(MultiplyAccumulate_39_io_activations_2),
    .io_activations_3(MultiplyAccumulate_39_io_activations_3),
    .io_weights(MultiplyAccumulate_39_io_weights),
    .io_sum(MultiplyAccumulate_39_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_40 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_40_clock),
    .io_activations_0(MultiplyAccumulate_40_io_activations_0),
    .io_activations_1(MultiplyAccumulate_40_io_activations_1),
    .io_activations_2(MultiplyAccumulate_40_io_activations_2),
    .io_activations_3(MultiplyAccumulate_40_io_activations_3),
    .io_weights(MultiplyAccumulate_40_io_weights),
    .io_sum(MultiplyAccumulate_40_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_41 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_41_clock),
    .io_activations_0(MultiplyAccumulate_41_io_activations_0),
    .io_activations_1(MultiplyAccumulate_41_io_activations_1),
    .io_activations_2(MultiplyAccumulate_41_io_activations_2),
    .io_activations_3(MultiplyAccumulate_41_io_activations_3),
    .io_weights(MultiplyAccumulate_41_io_weights),
    .io_sum(MultiplyAccumulate_41_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_42 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_42_clock),
    .io_activations_0(MultiplyAccumulate_42_io_activations_0),
    .io_activations_1(MultiplyAccumulate_42_io_activations_1),
    .io_activations_2(MultiplyAccumulate_42_io_activations_2),
    .io_activations_3(MultiplyAccumulate_42_io_activations_3),
    .io_weights(MultiplyAccumulate_42_io_weights),
    .io_sum(MultiplyAccumulate_42_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_43 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_43_clock),
    .io_activations_0(MultiplyAccumulate_43_io_activations_0),
    .io_activations_1(MultiplyAccumulate_43_io_activations_1),
    .io_activations_2(MultiplyAccumulate_43_io_activations_2),
    .io_activations_3(MultiplyAccumulate_43_io_activations_3),
    .io_weights(MultiplyAccumulate_43_io_weights),
    .io_sum(MultiplyAccumulate_43_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_44 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_44_clock),
    .io_activations_0(MultiplyAccumulate_44_io_activations_0),
    .io_activations_1(MultiplyAccumulate_44_io_activations_1),
    .io_activations_2(MultiplyAccumulate_44_io_activations_2),
    .io_activations_3(MultiplyAccumulate_44_io_activations_3),
    .io_weights(MultiplyAccumulate_44_io_weights),
    .io_sum(MultiplyAccumulate_44_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_45 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_45_clock),
    .io_activations_0(MultiplyAccumulate_45_io_activations_0),
    .io_activations_1(MultiplyAccumulate_45_io_activations_1),
    .io_activations_2(MultiplyAccumulate_45_io_activations_2),
    .io_activations_3(MultiplyAccumulate_45_io_activations_3),
    .io_weights(MultiplyAccumulate_45_io_weights),
    .io_sum(MultiplyAccumulate_45_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_46 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_46_clock),
    .io_activations_0(MultiplyAccumulate_46_io_activations_0),
    .io_activations_1(MultiplyAccumulate_46_io_activations_1),
    .io_activations_2(MultiplyAccumulate_46_io_activations_2),
    .io_activations_3(MultiplyAccumulate_46_io_activations_3),
    .io_weights(MultiplyAccumulate_46_io_weights),
    .io_sum(MultiplyAccumulate_46_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_47 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_47_clock),
    .io_activations_0(MultiplyAccumulate_47_io_activations_0),
    .io_activations_1(MultiplyAccumulate_47_io_activations_1),
    .io_activations_2(MultiplyAccumulate_47_io_activations_2),
    .io_activations_3(MultiplyAccumulate_47_io_activations_3),
    .io_weights(MultiplyAccumulate_47_io_weights),
    .io_sum(MultiplyAccumulate_47_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_48 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_48_clock),
    .io_activations_0(MultiplyAccumulate_48_io_activations_0),
    .io_activations_1(MultiplyAccumulate_48_io_activations_1),
    .io_activations_2(MultiplyAccumulate_48_io_activations_2),
    .io_activations_3(MultiplyAccumulate_48_io_activations_3),
    .io_weights(MultiplyAccumulate_48_io_weights),
    .io_sum(MultiplyAccumulate_48_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_49 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_49_clock),
    .io_activations_0(MultiplyAccumulate_49_io_activations_0),
    .io_activations_1(MultiplyAccumulate_49_io_activations_1),
    .io_activations_2(MultiplyAccumulate_49_io_activations_2),
    .io_activations_3(MultiplyAccumulate_49_io_activations_3),
    .io_weights(MultiplyAccumulate_49_io_weights),
    .io_sum(MultiplyAccumulate_49_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_50 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_50_clock),
    .io_activations_0(MultiplyAccumulate_50_io_activations_0),
    .io_activations_1(MultiplyAccumulate_50_io_activations_1),
    .io_activations_2(MultiplyAccumulate_50_io_activations_2),
    .io_activations_3(MultiplyAccumulate_50_io_activations_3),
    .io_weights(MultiplyAccumulate_50_io_weights),
    .io_sum(MultiplyAccumulate_50_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_51 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_51_clock),
    .io_activations_0(MultiplyAccumulate_51_io_activations_0),
    .io_activations_1(MultiplyAccumulate_51_io_activations_1),
    .io_activations_2(MultiplyAccumulate_51_io_activations_2),
    .io_activations_3(MultiplyAccumulate_51_io_activations_3),
    .io_weights(MultiplyAccumulate_51_io_weights),
    .io_sum(MultiplyAccumulate_51_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_52 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_52_clock),
    .io_activations_0(MultiplyAccumulate_52_io_activations_0),
    .io_activations_1(MultiplyAccumulate_52_io_activations_1),
    .io_activations_2(MultiplyAccumulate_52_io_activations_2),
    .io_activations_3(MultiplyAccumulate_52_io_activations_3),
    .io_weights(MultiplyAccumulate_52_io_weights),
    .io_sum(MultiplyAccumulate_52_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_53 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_53_clock),
    .io_activations_0(MultiplyAccumulate_53_io_activations_0),
    .io_activations_1(MultiplyAccumulate_53_io_activations_1),
    .io_activations_2(MultiplyAccumulate_53_io_activations_2),
    .io_activations_3(MultiplyAccumulate_53_io_activations_3),
    .io_weights(MultiplyAccumulate_53_io_weights),
    .io_sum(MultiplyAccumulate_53_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_54 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_54_clock),
    .io_activations_0(MultiplyAccumulate_54_io_activations_0),
    .io_activations_1(MultiplyAccumulate_54_io_activations_1),
    .io_activations_2(MultiplyAccumulate_54_io_activations_2),
    .io_activations_3(MultiplyAccumulate_54_io_activations_3),
    .io_weights(MultiplyAccumulate_54_io_weights),
    .io_sum(MultiplyAccumulate_54_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_55 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_55_clock),
    .io_activations_0(MultiplyAccumulate_55_io_activations_0),
    .io_activations_1(MultiplyAccumulate_55_io_activations_1),
    .io_activations_2(MultiplyAccumulate_55_io_activations_2),
    .io_activations_3(MultiplyAccumulate_55_io_activations_3),
    .io_weights(MultiplyAccumulate_55_io_weights),
    .io_sum(MultiplyAccumulate_55_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_56 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_56_clock),
    .io_activations_0(MultiplyAccumulate_56_io_activations_0),
    .io_activations_1(MultiplyAccumulate_56_io_activations_1),
    .io_activations_2(MultiplyAccumulate_56_io_activations_2),
    .io_activations_3(MultiplyAccumulate_56_io_activations_3),
    .io_weights(MultiplyAccumulate_56_io_weights),
    .io_sum(MultiplyAccumulate_56_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_57 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_57_clock),
    .io_activations_0(MultiplyAccumulate_57_io_activations_0),
    .io_activations_1(MultiplyAccumulate_57_io_activations_1),
    .io_activations_2(MultiplyAccumulate_57_io_activations_2),
    .io_activations_3(MultiplyAccumulate_57_io_activations_3),
    .io_weights(MultiplyAccumulate_57_io_weights),
    .io_sum(MultiplyAccumulate_57_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_58 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_58_clock),
    .io_activations_0(MultiplyAccumulate_58_io_activations_0),
    .io_activations_1(MultiplyAccumulate_58_io_activations_1),
    .io_activations_2(MultiplyAccumulate_58_io_activations_2),
    .io_activations_3(MultiplyAccumulate_58_io_activations_3),
    .io_weights(MultiplyAccumulate_58_io_weights),
    .io_sum(MultiplyAccumulate_58_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_59 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_59_clock),
    .io_activations_0(MultiplyAccumulate_59_io_activations_0),
    .io_activations_1(MultiplyAccumulate_59_io_activations_1),
    .io_activations_2(MultiplyAccumulate_59_io_activations_2),
    .io_activations_3(MultiplyAccumulate_59_io_activations_3),
    .io_weights(MultiplyAccumulate_59_io_weights),
    .io_sum(MultiplyAccumulate_59_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_60 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_60_clock),
    .io_activations_0(MultiplyAccumulate_60_io_activations_0),
    .io_activations_1(MultiplyAccumulate_60_io_activations_1),
    .io_activations_2(MultiplyAccumulate_60_io_activations_2),
    .io_activations_3(MultiplyAccumulate_60_io_activations_3),
    .io_weights(MultiplyAccumulate_60_io_weights),
    .io_sum(MultiplyAccumulate_60_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_61 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_61_clock),
    .io_activations_0(MultiplyAccumulate_61_io_activations_0),
    .io_activations_1(MultiplyAccumulate_61_io_activations_1),
    .io_activations_2(MultiplyAccumulate_61_io_activations_2),
    .io_activations_3(MultiplyAccumulate_61_io_activations_3),
    .io_weights(MultiplyAccumulate_61_io_weights),
    .io_sum(MultiplyAccumulate_61_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_62 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_62_clock),
    .io_activations_0(MultiplyAccumulate_62_io_activations_0),
    .io_activations_1(MultiplyAccumulate_62_io_activations_1),
    .io_activations_2(MultiplyAccumulate_62_io_activations_2),
    .io_activations_3(MultiplyAccumulate_62_io_activations_3),
    .io_weights(MultiplyAccumulate_62_io_weights),
    .io_sum(MultiplyAccumulate_62_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_63 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_63_clock),
    .io_activations_0(MultiplyAccumulate_63_io_activations_0),
    .io_activations_1(MultiplyAccumulate_63_io_activations_1),
    .io_activations_2(MultiplyAccumulate_63_io_activations_2),
    .io_activations_3(MultiplyAccumulate_63_io_activations_3),
    .io_weights(MultiplyAccumulate_63_io_weights),
    .io_sum(MultiplyAccumulate_63_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_64 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_64_clock),
    .io_activations_0(MultiplyAccumulate_64_io_activations_0),
    .io_activations_1(MultiplyAccumulate_64_io_activations_1),
    .io_activations_2(MultiplyAccumulate_64_io_activations_2),
    .io_activations_3(MultiplyAccumulate_64_io_activations_3),
    .io_weights(MultiplyAccumulate_64_io_weights),
    .io_sum(MultiplyAccumulate_64_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_65 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_65_clock),
    .io_activations_0(MultiplyAccumulate_65_io_activations_0),
    .io_activations_1(MultiplyAccumulate_65_io_activations_1),
    .io_activations_2(MultiplyAccumulate_65_io_activations_2),
    .io_activations_3(MultiplyAccumulate_65_io_activations_3),
    .io_weights(MultiplyAccumulate_65_io_weights),
    .io_sum(MultiplyAccumulate_65_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_66 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_66_clock),
    .io_activations_0(MultiplyAccumulate_66_io_activations_0),
    .io_activations_1(MultiplyAccumulate_66_io_activations_1),
    .io_activations_2(MultiplyAccumulate_66_io_activations_2),
    .io_activations_3(MultiplyAccumulate_66_io_activations_3),
    .io_weights(MultiplyAccumulate_66_io_weights),
    .io_sum(MultiplyAccumulate_66_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_67 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_67_clock),
    .io_activations_0(MultiplyAccumulate_67_io_activations_0),
    .io_activations_1(MultiplyAccumulate_67_io_activations_1),
    .io_activations_2(MultiplyAccumulate_67_io_activations_2),
    .io_activations_3(MultiplyAccumulate_67_io_activations_3),
    .io_weights(MultiplyAccumulate_67_io_weights),
    .io_sum(MultiplyAccumulate_67_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_68 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_68_clock),
    .io_activations_0(MultiplyAccumulate_68_io_activations_0),
    .io_activations_1(MultiplyAccumulate_68_io_activations_1),
    .io_activations_2(MultiplyAccumulate_68_io_activations_2),
    .io_activations_3(MultiplyAccumulate_68_io_activations_3),
    .io_weights(MultiplyAccumulate_68_io_weights),
    .io_sum(MultiplyAccumulate_68_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_69 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_69_clock),
    .io_activations_0(MultiplyAccumulate_69_io_activations_0),
    .io_activations_1(MultiplyAccumulate_69_io_activations_1),
    .io_activations_2(MultiplyAccumulate_69_io_activations_2),
    .io_activations_3(MultiplyAccumulate_69_io_activations_3),
    .io_weights(MultiplyAccumulate_69_io_weights),
    .io_sum(MultiplyAccumulate_69_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_70 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_70_clock),
    .io_activations_0(MultiplyAccumulate_70_io_activations_0),
    .io_activations_1(MultiplyAccumulate_70_io_activations_1),
    .io_activations_2(MultiplyAccumulate_70_io_activations_2),
    .io_activations_3(MultiplyAccumulate_70_io_activations_3),
    .io_weights(MultiplyAccumulate_70_io_weights),
    .io_sum(MultiplyAccumulate_70_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_71 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_71_clock),
    .io_activations_0(MultiplyAccumulate_71_io_activations_0),
    .io_activations_1(MultiplyAccumulate_71_io_activations_1),
    .io_activations_2(MultiplyAccumulate_71_io_activations_2),
    .io_activations_3(MultiplyAccumulate_71_io_activations_3),
    .io_weights(MultiplyAccumulate_71_io_weights),
    .io_sum(MultiplyAccumulate_71_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_72 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_72_clock),
    .io_activations_0(MultiplyAccumulate_72_io_activations_0),
    .io_activations_1(MultiplyAccumulate_72_io_activations_1),
    .io_activations_2(MultiplyAccumulate_72_io_activations_2),
    .io_activations_3(MultiplyAccumulate_72_io_activations_3),
    .io_weights(MultiplyAccumulate_72_io_weights),
    .io_sum(MultiplyAccumulate_72_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_73 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_73_clock),
    .io_activations_0(MultiplyAccumulate_73_io_activations_0),
    .io_activations_1(MultiplyAccumulate_73_io_activations_1),
    .io_activations_2(MultiplyAccumulate_73_io_activations_2),
    .io_activations_3(MultiplyAccumulate_73_io_activations_3),
    .io_weights(MultiplyAccumulate_73_io_weights),
    .io_sum(MultiplyAccumulate_73_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_74 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_74_clock),
    .io_activations_0(MultiplyAccumulate_74_io_activations_0),
    .io_activations_1(MultiplyAccumulate_74_io_activations_1),
    .io_activations_2(MultiplyAccumulate_74_io_activations_2),
    .io_activations_3(MultiplyAccumulate_74_io_activations_3),
    .io_weights(MultiplyAccumulate_74_io_weights),
    .io_sum(MultiplyAccumulate_74_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_75 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_75_clock),
    .io_activations_0(MultiplyAccumulate_75_io_activations_0),
    .io_activations_1(MultiplyAccumulate_75_io_activations_1),
    .io_activations_2(MultiplyAccumulate_75_io_activations_2),
    .io_activations_3(MultiplyAccumulate_75_io_activations_3),
    .io_weights(MultiplyAccumulate_75_io_weights),
    .io_sum(MultiplyAccumulate_75_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_76 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_76_clock),
    .io_activations_0(MultiplyAccumulate_76_io_activations_0),
    .io_activations_1(MultiplyAccumulate_76_io_activations_1),
    .io_activations_2(MultiplyAccumulate_76_io_activations_2),
    .io_activations_3(MultiplyAccumulate_76_io_activations_3),
    .io_weights(MultiplyAccumulate_76_io_weights),
    .io_sum(MultiplyAccumulate_76_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_77 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_77_clock),
    .io_activations_0(MultiplyAccumulate_77_io_activations_0),
    .io_activations_1(MultiplyAccumulate_77_io_activations_1),
    .io_activations_2(MultiplyAccumulate_77_io_activations_2),
    .io_activations_3(MultiplyAccumulate_77_io_activations_3),
    .io_weights(MultiplyAccumulate_77_io_weights),
    .io_sum(MultiplyAccumulate_77_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_78 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_78_clock),
    .io_activations_0(MultiplyAccumulate_78_io_activations_0),
    .io_activations_1(MultiplyAccumulate_78_io_activations_1),
    .io_activations_2(MultiplyAccumulate_78_io_activations_2),
    .io_activations_3(MultiplyAccumulate_78_io_activations_3),
    .io_weights(MultiplyAccumulate_78_io_weights),
    .io_sum(MultiplyAccumulate_78_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_79 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_79_clock),
    .io_activations_0(MultiplyAccumulate_79_io_activations_0),
    .io_activations_1(MultiplyAccumulate_79_io_activations_1),
    .io_activations_2(MultiplyAccumulate_79_io_activations_2),
    .io_activations_3(MultiplyAccumulate_79_io_activations_3),
    .io_weights(MultiplyAccumulate_79_io_weights),
    .io_sum(MultiplyAccumulate_79_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_80 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_80_clock),
    .io_activations_0(MultiplyAccumulate_80_io_activations_0),
    .io_activations_1(MultiplyAccumulate_80_io_activations_1),
    .io_activations_2(MultiplyAccumulate_80_io_activations_2),
    .io_activations_3(MultiplyAccumulate_80_io_activations_3),
    .io_weights(MultiplyAccumulate_80_io_weights),
    .io_sum(MultiplyAccumulate_80_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_81 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_81_clock),
    .io_activations_0(MultiplyAccumulate_81_io_activations_0),
    .io_activations_1(MultiplyAccumulate_81_io_activations_1),
    .io_activations_2(MultiplyAccumulate_81_io_activations_2),
    .io_activations_3(MultiplyAccumulate_81_io_activations_3),
    .io_weights(MultiplyAccumulate_81_io_weights),
    .io_sum(MultiplyAccumulate_81_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_82 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_82_clock),
    .io_activations_0(MultiplyAccumulate_82_io_activations_0),
    .io_activations_1(MultiplyAccumulate_82_io_activations_1),
    .io_activations_2(MultiplyAccumulate_82_io_activations_2),
    .io_activations_3(MultiplyAccumulate_82_io_activations_3),
    .io_weights(MultiplyAccumulate_82_io_weights),
    .io_sum(MultiplyAccumulate_82_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_83 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_83_clock),
    .io_activations_0(MultiplyAccumulate_83_io_activations_0),
    .io_activations_1(MultiplyAccumulate_83_io_activations_1),
    .io_activations_2(MultiplyAccumulate_83_io_activations_2),
    .io_activations_3(MultiplyAccumulate_83_io_activations_3),
    .io_weights(MultiplyAccumulate_83_io_weights),
    .io_sum(MultiplyAccumulate_83_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_84 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_84_clock),
    .io_activations_0(MultiplyAccumulate_84_io_activations_0),
    .io_activations_1(MultiplyAccumulate_84_io_activations_1),
    .io_activations_2(MultiplyAccumulate_84_io_activations_2),
    .io_activations_3(MultiplyAccumulate_84_io_activations_3),
    .io_weights(MultiplyAccumulate_84_io_weights),
    .io_sum(MultiplyAccumulate_84_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_85 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_85_clock),
    .io_activations_0(MultiplyAccumulate_85_io_activations_0),
    .io_activations_1(MultiplyAccumulate_85_io_activations_1),
    .io_activations_2(MultiplyAccumulate_85_io_activations_2),
    .io_activations_3(MultiplyAccumulate_85_io_activations_3),
    .io_weights(MultiplyAccumulate_85_io_weights),
    .io_sum(MultiplyAccumulate_85_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_86 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_86_clock),
    .io_activations_0(MultiplyAccumulate_86_io_activations_0),
    .io_activations_1(MultiplyAccumulate_86_io_activations_1),
    .io_activations_2(MultiplyAccumulate_86_io_activations_2),
    .io_activations_3(MultiplyAccumulate_86_io_activations_3),
    .io_weights(MultiplyAccumulate_86_io_weights),
    .io_sum(MultiplyAccumulate_86_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_87 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_87_clock),
    .io_activations_0(MultiplyAccumulate_87_io_activations_0),
    .io_activations_1(MultiplyAccumulate_87_io_activations_1),
    .io_activations_2(MultiplyAccumulate_87_io_activations_2),
    .io_activations_3(MultiplyAccumulate_87_io_activations_3),
    .io_weights(MultiplyAccumulate_87_io_weights),
    .io_sum(MultiplyAccumulate_87_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_88 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_88_clock),
    .io_activations_0(MultiplyAccumulate_88_io_activations_0),
    .io_activations_1(MultiplyAccumulate_88_io_activations_1),
    .io_activations_2(MultiplyAccumulate_88_io_activations_2),
    .io_activations_3(MultiplyAccumulate_88_io_activations_3),
    .io_weights(MultiplyAccumulate_88_io_weights),
    .io_sum(MultiplyAccumulate_88_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_89 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_89_clock),
    .io_activations_0(MultiplyAccumulate_89_io_activations_0),
    .io_activations_1(MultiplyAccumulate_89_io_activations_1),
    .io_activations_2(MultiplyAccumulate_89_io_activations_2),
    .io_activations_3(MultiplyAccumulate_89_io_activations_3),
    .io_weights(MultiplyAccumulate_89_io_weights),
    .io_sum(MultiplyAccumulate_89_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_90 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_90_clock),
    .io_activations_0(MultiplyAccumulate_90_io_activations_0),
    .io_activations_1(MultiplyAccumulate_90_io_activations_1),
    .io_activations_2(MultiplyAccumulate_90_io_activations_2),
    .io_activations_3(MultiplyAccumulate_90_io_activations_3),
    .io_weights(MultiplyAccumulate_90_io_weights),
    .io_sum(MultiplyAccumulate_90_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_91 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_91_clock),
    .io_activations_0(MultiplyAccumulate_91_io_activations_0),
    .io_activations_1(MultiplyAccumulate_91_io_activations_1),
    .io_activations_2(MultiplyAccumulate_91_io_activations_2),
    .io_activations_3(MultiplyAccumulate_91_io_activations_3),
    .io_weights(MultiplyAccumulate_91_io_weights),
    .io_sum(MultiplyAccumulate_91_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_92 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_92_clock),
    .io_activations_0(MultiplyAccumulate_92_io_activations_0),
    .io_activations_1(MultiplyAccumulate_92_io_activations_1),
    .io_activations_2(MultiplyAccumulate_92_io_activations_2),
    .io_activations_3(MultiplyAccumulate_92_io_activations_3),
    .io_weights(MultiplyAccumulate_92_io_weights),
    .io_sum(MultiplyAccumulate_92_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_93 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_93_clock),
    .io_activations_0(MultiplyAccumulate_93_io_activations_0),
    .io_activations_1(MultiplyAccumulate_93_io_activations_1),
    .io_activations_2(MultiplyAccumulate_93_io_activations_2),
    .io_activations_3(MultiplyAccumulate_93_io_activations_3),
    .io_weights(MultiplyAccumulate_93_io_weights),
    .io_sum(MultiplyAccumulate_93_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_94 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_94_clock),
    .io_activations_0(MultiplyAccumulate_94_io_activations_0),
    .io_activations_1(MultiplyAccumulate_94_io_activations_1),
    .io_activations_2(MultiplyAccumulate_94_io_activations_2),
    .io_activations_3(MultiplyAccumulate_94_io_activations_3),
    .io_weights(MultiplyAccumulate_94_io_weights),
    .io_sum(MultiplyAccumulate_94_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_95 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_95_clock),
    .io_activations_0(MultiplyAccumulate_95_io_activations_0),
    .io_activations_1(MultiplyAccumulate_95_io_activations_1),
    .io_activations_2(MultiplyAccumulate_95_io_activations_2),
    .io_activations_3(MultiplyAccumulate_95_io_activations_3),
    .io_weights(MultiplyAccumulate_95_io_weights),
    .io_sum(MultiplyAccumulate_95_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_96 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_96_clock),
    .io_activations_0(MultiplyAccumulate_96_io_activations_0),
    .io_activations_1(MultiplyAccumulate_96_io_activations_1),
    .io_activations_2(MultiplyAccumulate_96_io_activations_2),
    .io_activations_3(MultiplyAccumulate_96_io_activations_3),
    .io_weights(MultiplyAccumulate_96_io_weights),
    .io_sum(MultiplyAccumulate_96_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_97 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_97_clock),
    .io_activations_0(MultiplyAccumulate_97_io_activations_0),
    .io_activations_1(MultiplyAccumulate_97_io_activations_1),
    .io_activations_2(MultiplyAccumulate_97_io_activations_2),
    .io_activations_3(MultiplyAccumulate_97_io_activations_3),
    .io_weights(MultiplyAccumulate_97_io_weights),
    .io_sum(MultiplyAccumulate_97_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_98 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_98_clock),
    .io_activations_0(MultiplyAccumulate_98_io_activations_0),
    .io_activations_1(MultiplyAccumulate_98_io_activations_1),
    .io_activations_2(MultiplyAccumulate_98_io_activations_2),
    .io_activations_3(MultiplyAccumulate_98_io_activations_3),
    .io_weights(MultiplyAccumulate_98_io_weights),
    .io_sum(MultiplyAccumulate_98_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_99 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_99_clock),
    .io_activations_0(MultiplyAccumulate_99_io_activations_0),
    .io_activations_1(MultiplyAccumulate_99_io_activations_1),
    .io_activations_2(MultiplyAccumulate_99_io_activations_2),
    .io_activations_3(MultiplyAccumulate_99_io_activations_3),
    .io_weights(MultiplyAccumulate_99_io_weights),
    .io_sum(MultiplyAccumulate_99_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_100 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_100_clock),
    .io_activations_0(MultiplyAccumulate_100_io_activations_0),
    .io_activations_1(MultiplyAccumulate_100_io_activations_1),
    .io_activations_2(MultiplyAccumulate_100_io_activations_2),
    .io_activations_3(MultiplyAccumulate_100_io_activations_3),
    .io_weights(MultiplyAccumulate_100_io_weights),
    .io_sum(MultiplyAccumulate_100_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_101 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_101_clock),
    .io_activations_0(MultiplyAccumulate_101_io_activations_0),
    .io_activations_1(MultiplyAccumulate_101_io_activations_1),
    .io_activations_2(MultiplyAccumulate_101_io_activations_2),
    .io_activations_3(MultiplyAccumulate_101_io_activations_3),
    .io_weights(MultiplyAccumulate_101_io_weights),
    .io_sum(MultiplyAccumulate_101_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_102 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_102_clock),
    .io_activations_0(MultiplyAccumulate_102_io_activations_0),
    .io_activations_1(MultiplyAccumulate_102_io_activations_1),
    .io_activations_2(MultiplyAccumulate_102_io_activations_2),
    .io_activations_3(MultiplyAccumulate_102_io_activations_3),
    .io_weights(MultiplyAccumulate_102_io_weights),
    .io_sum(MultiplyAccumulate_102_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_103 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_103_clock),
    .io_activations_0(MultiplyAccumulate_103_io_activations_0),
    .io_activations_1(MultiplyAccumulate_103_io_activations_1),
    .io_activations_2(MultiplyAccumulate_103_io_activations_2),
    .io_activations_3(MultiplyAccumulate_103_io_activations_3),
    .io_weights(MultiplyAccumulate_103_io_weights),
    .io_sum(MultiplyAccumulate_103_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_104 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_104_clock),
    .io_activations_0(MultiplyAccumulate_104_io_activations_0),
    .io_activations_1(MultiplyAccumulate_104_io_activations_1),
    .io_activations_2(MultiplyAccumulate_104_io_activations_2),
    .io_activations_3(MultiplyAccumulate_104_io_activations_3),
    .io_weights(MultiplyAccumulate_104_io_weights),
    .io_sum(MultiplyAccumulate_104_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_105 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_105_clock),
    .io_activations_0(MultiplyAccumulate_105_io_activations_0),
    .io_activations_1(MultiplyAccumulate_105_io_activations_1),
    .io_activations_2(MultiplyAccumulate_105_io_activations_2),
    .io_activations_3(MultiplyAccumulate_105_io_activations_3),
    .io_weights(MultiplyAccumulate_105_io_weights),
    .io_sum(MultiplyAccumulate_105_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_106 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_106_clock),
    .io_activations_0(MultiplyAccumulate_106_io_activations_0),
    .io_activations_1(MultiplyAccumulate_106_io_activations_1),
    .io_activations_2(MultiplyAccumulate_106_io_activations_2),
    .io_activations_3(MultiplyAccumulate_106_io_activations_3),
    .io_weights(MultiplyAccumulate_106_io_weights),
    .io_sum(MultiplyAccumulate_106_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_107 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_107_clock),
    .io_activations_0(MultiplyAccumulate_107_io_activations_0),
    .io_activations_1(MultiplyAccumulate_107_io_activations_1),
    .io_activations_2(MultiplyAccumulate_107_io_activations_2),
    .io_activations_3(MultiplyAccumulate_107_io_activations_3),
    .io_weights(MultiplyAccumulate_107_io_weights),
    .io_sum(MultiplyAccumulate_107_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_108 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_108_clock),
    .io_activations_0(MultiplyAccumulate_108_io_activations_0),
    .io_activations_1(MultiplyAccumulate_108_io_activations_1),
    .io_activations_2(MultiplyAccumulate_108_io_activations_2),
    .io_activations_3(MultiplyAccumulate_108_io_activations_3),
    .io_weights(MultiplyAccumulate_108_io_weights),
    .io_sum(MultiplyAccumulate_108_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_109 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_109_clock),
    .io_activations_0(MultiplyAccumulate_109_io_activations_0),
    .io_activations_1(MultiplyAccumulate_109_io_activations_1),
    .io_activations_2(MultiplyAccumulate_109_io_activations_2),
    .io_activations_3(MultiplyAccumulate_109_io_activations_3),
    .io_weights(MultiplyAccumulate_109_io_weights),
    .io_sum(MultiplyAccumulate_109_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_110 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_110_clock),
    .io_activations_0(MultiplyAccumulate_110_io_activations_0),
    .io_activations_1(MultiplyAccumulate_110_io_activations_1),
    .io_activations_2(MultiplyAccumulate_110_io_activations_2),
    .io_activations_3(MultiplyAccumulate_110_io_activations_3),
    .io_weights(MultiplyAccumulate_110_io_weights),
    .io_sum(MultiplyAccumulate_110_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_111 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_111_clock),
    .io_activations_0(MultiplyAccumulate_111_io_activations_0),
    .io_activations_1(MultiplyAccumulate_111_io_activations_1),
    .io_activations_2(MultiplyAccumulate_111_io_activations_2),
    .io_activations_3(MultiplyAccumulate_111_io_activations_3),
    .io_weights(MultiplyAccumulate_111_io_weights),
    .io_sum(MultiplyAccumulate_111_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_112 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_112_clock),
    .io_activations_0(MultiplyAccumulate_112_io_activations_0),
    .io_activations_1(MultiplyAccumulate_112_io_activations_1),
    .io_activations_2(MultiplyAccumulate_112_io_activations_2),
    .io_activations_3(MultiplyAccumulate_112_io_activations_3),
    .io_weights(MultiplyAccumulate_112_io_weights),
    .io_sum(MultiplyAccumulate_112_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_113 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_113_clock),
    .io_activations_0(MultiplyAccumulate_113_io_activations_0),
    .io_activations_1(MultiplyAccumulate_113_io_activations_1),
    .io_activations_2(MultiplyAccumulate_113_io_activations_2),
    .io_activations_3(MultiplyAccumulate_113_io_activations_3),
    .io_weights(MultiplyAccumulate_113_io_weights),
    .io_sum(MultiplyAccumulate_113_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_114 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_114_clock),
    .io_activations_0(MultiplyAccumulate_114_io_activations_0),
    .io_activations_1(MultiplyAccumulate_114_io_activations_1),
    .io_activations_2(MultiplyAccumulate_114_io_activations_2),
    .io_activations_3(MultiplyAccumulate_114_io_activations_3),
    .io_weights(MultiplyAccumulate_114_io_weights),
    .io_sum(MultiplyAccumulate_114_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_115 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_115_clock),
    .io_activations_0(MultiplyAccumulate_115_io_activations_0),
    .io_activations_1(MultiplyAccumulate_115_io_activations_1),
    .io_activations_2(MultiplyAccumulate_115_io_activations_2),
    .io_activations_3(MultiplyAccumulate_115_io_activations_3),
    .io_weights(MultiplyAccumulate_115_io_weights),
    .io_sum(MultiplyAccumulate_115_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_116 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_116_clock),
    .io_activations_0(MultiplyAccumulate_116_io_activations_0),
    .io_activations_1(MultiplyAccumulate_116_io_activations_1),
    .io_activations_2(MultiplyAccumulate_116_io_activations_2),
    .io_activations_3(MultiplyAccumulate_116_io_activations_3),
    .io_weights(MultiplyAccumulate_116_io_weights),
    .io_sum(MultiplyAccumulate_116_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_117 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_117_clock),
    .io_activations_0(MultiplyAccumulate_117_io_activations_0),
    .io_activations_1(MultiplyAccumulate_117_io_activations_1),
    .io_activations_2(MultiplyAccumulate_117_io_activations_2),
    .io_activations_3(MultiplyAccumulate_117_io_activations_3),
    .io_weights(MultiplyAccumulate_117_io_weights),
    .io_sum(MultiplyAccumulate_117_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_118 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_118_clock),
    .io_activations_0(MultiplyAccumulate_118_io_activations_0),
    .io_activations_1(MultiplyAccumulate_118_io_activations_1),
    .io_activations_2(MultiplyAccumulate_118_io_activations_2),
    .io_activations_3(MultiplyAccumulate_118_io_activations_3),
    .io_weights(MultiplyAccumulate_118_io_weights),
    .io_sum(MultiplyAccumulate_118_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_119 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_119_clock),
    .io_activations_0(MultiplyAccumulate_119_io_activations_0),
    .io_activations_1(MultiplyAccumulate_119_io_activations_1),
    .io_activations_2(MultiplyAccumulate_119_io_activations_2),
    .io_activations_3(MultiplyAccumulate_119_io_activations_3),
    .io_weights(MultiplyAccumulate_119_io_weights),
    .io_sum(MultiplyAccumulate_119_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_120 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_120_clock),
    .io_activations_0(MultiplyAccumulate_120_io_activations_0),
    .io_activations_1(MultiplyAccumulate_120_io_activations_1),
    .io_activations_2(MultiplyAccumulate_120_io_activations_2),
    .io_activations_3(MultiplyAccumulate_120_io_activations_3),
    .io_weights(MultiplyAccumulate_120_io_weights),
    .io_sum(MultiplyAccumulate_120_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_121 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_121_clock),
    .io_activations_0(MultiplyAccumulate_121_io_activations_0),
    .io_activations_1(MultiplyAccumulate_121_io_activations_1),
    .io_activations_2(MultiplyAccumulate_121_io_activations_2),
    .io_activations_3(MultiplyAccumulate_121_io_activations_3),
    .io_weights(MultiplyAccumulate_121_io_weights),
    .io_sum(MultiplyAccumulate_121_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_122 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_122_clock),
    .io_activations_0(MultiplyAccumulate_122_io_activations_0),
    .io_activations_1(MultiplyAccumulate_122_io_activations_1),
    .io_activations_2(MultiplyAccumulate_122_io_activations_2),
    .io_activations_3(MultiplyAccumulate_122_io_activations_3),
    .io_weights(MultiplyAccumulate_122_io_weights),
    .io_sum(MultiplyAccumulate_122_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_123 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_123_clock),
    .io_activations_0(MultiplyAccumulate_123_io_activations_0),
    .io_activations_1(MultiplyAccumulate_123_io_activations_1),
    .io_activations_2(MultiplyAccumulate_123_io_activations_2),
    .io_activations_3(MultiplyAccumulate_123_io_activations_3),
    .io_weights(MultiplyAccumulate_123_io_weights),
    .io_sum(MultiplyAccumulate_123_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_124 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_124_clock),
    .io_activations_0(MultiplyAccumulate_124_io_activations_0),
    .io_activations_1(MultiplyAccumulate_124_io_activations_1),
    .io_activations_2(MultiplyAccumulate_124_io_activations_2),
    .io_activations_3(MultiplyAccumulate_124_io_activations_3),
    .io_weights(MultiplyAccumulate_124_io_weights),
    .io_sum(MultiplyAccumulate_124_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_125 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_125_clock),
    .io_activations_0(MultiplyAccumulate_125_io_activations_0),
    .io_activations_1(MultiplyAccumulate_125_io_activations_1),
    .io_activations_2(MultiplyAccumulate_125_io_activations_2),
    .io_activations_3(MultiplyAccumulate_125_io_activations_3),
    .io_weights(MultiplyAccumulate_125_io_weights),
    .io_sum(MultiplyAccumulate_125_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_126 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_126_clock),
    .io_activations_0(MultiplyAccumulate_126_io_activations_0),
    .io_activations_1(MultiplyAccumulate_126_io_activations_1),
    .io_activations_2(MultiplyAccumulate_126_io_activations_2),
    .io_activations_3(MultiplyAccumulate_126_io_activations_3),
    .io_weights(MultiplyAccumulate_126_io_weights),
    .io_sum(MultiplyAccumulate_126_io_sum)
  );
  MultiplyAccumulate MultiplyAccumulate_127 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_127_clock),
    .io_activations_0(MultiplyAccumulate_127_io_activations_0),
    .io_activations_1(MultiplyAccumulate_127_io_activations_1),
    .io_activations_2(MultiplyAccumulate_127_io_activations_2),
    .io_activations_3(MultiplyAccumulate_127_io_activations_3),
    .io_weights(MultiplyAccumulate_127_io_weights),
    .io_sum(MultiplyAccumulate_127_io_sum)
  );
  assign _T_158 = cntr + 10'h1; // @[DenseLayer.scala 90:18]
  assign _T_159 = _T_158[9:0]; // @[DenseLayer.scala 90:18]
  assign _GEN_0 = io_dataIn_valid ? _T_159 : cntr; // @[DenseLayer.scala 89:28]
  assign currWeights_0 = weightsRAM_out[7:0]; // @[DenseLayer.scala 100:42]
  assign currWeights_1 = weightsRAM_out[15:8]; // @[DenseLayer.scala 100:42]
  assign currWeights_2 = weightsRAM_out[23:16]; // @[DenseLayer.scala 100:42]
  assign currWeights_3 = weightsRAM_out[31:24]; // @[DenseLayer.scala 100:42]
  assign currWeights_4 = weightsRAM_out[39:32]; // @[DenseLayer.scala 100:42]
  assign currWeights_5 = weightsRAM_out[47:40]; // @[DenseLayer.scala 100:42]
  assign currWeights_6 = weightsRAM_out[55:48]; // @[DenseLayer.scala 100:42]
  assign currWeights_7 = weightsRAM_out[63:56]; // @[DenseLayer.scala 100:42]
  assign currWeights_8 = weightsRAM_out[71:64]; // @[DenseLayer.scala 100:42]
  assign currWeights_9 = weightsRAM_out[79:72]; // @[DenseLayer.scala 100:42]
  assign currWeights_10 = weightsRAM_out[87:80]; // @[DenseLayer.scala 100:42]
  assign currWeights_11 = weightsRAM_out[95:88]; // @[DenseLayer.scala 100:42]
  assign currWeights_12 = weightsRAM_out[103:96]; // @[DenseLayer.scala 100:42]
  assign currWeights_13 = weightsRAM_out[111:104]; // @[DenseLayer.scala 100:42]
  assign currWeights_14 = weightsRAM_out[119:112]; // @[DenseLayer.scala 100:42]
  assign currWeights_15 = weightsRAM_out[127:120]; // @[DenseLayer.scala 100:42]
  assign currWeights_16 = weightsRAM_out[135:128]; // @[DenseLayer.scala 100:42]
  assign currWeights_17 = weightsRAM_out[143:136]; // @[DenseLayer.scala 100:42]
  assign currWeights_18 = weightsRAM_out[151:144]; // @[DenseLayer.scala 100:42]
  assign currWeights_19 = weightsRAM_out[159:152]; // @[DenseLayer.scala 100:42]
  assign currWeights_20 = weightsRAM_out[167:160]; // @[DenseLayer.scala 100:42]
  assign currWeights_21 = weightsRAM_out[175:168]; // @[DenseLayer.scala 100:42]
  assign currWeights_22 = weightsRAM_out[183:176]; // @[DenseLayer.scala 100:42]
  assign currWeights_23 = weightsRAM_out[191:184]; // @[DenseLayer.scala 100:42]
  assign currWeights_24 = weightsRAM_out[199:192]; // @[DenseLayer.scala 100:42]
  assign currWeights_25 = weightsRAM_out[207:200]; // @[DenseLayer.scala 100:42]
  assign currWeights_26 = weightsRAM_out[215:208]; // @[DenseLayer.scala 100:42]
  assign currWeights_27 = weightsRAM_out[223:216]; // @[DenseLayer.scala 100:42]
  assign currWeights_28 = weightsRAM_out[231:224]; // @[DenseLayer.scala 100:42]
  assign currWeights_29 = weightsRAM_out[239:232]; // @[DenseLayer.scala 100:42]
  assign currWeights_30 = weightsRAM_out[247:240]; // @[DenseLayer.scala 100:42]
  assign currWeights_31 = weightsRAM_out[255:248]; // @[DenseLayer.scala 100:42]
  assign currWeights_32 = weightsRAM_out[263:256]; // @[DenseLayer.scala 100:42]
  assign currWeights_33 = weightsRAM_out[271:264]; // @[DenseLayer.scala 100:42]
  assign currWeights_34 = weightsRAM_out[279:272]; // @[DenseLayer.scala 100:42]
  assign currWeights_35 = weightsRAM_out[287:280]; // @[DenseLayer.scala 100:42]
  assign currWeights_36 = weightsRAM_out[295:288]; // @[DenseLayer.scala 100:42]
  assign currWeights_37 = weightsRAM_out[303:296]; // @[DenseLayer.scala 100:42]
  assign currWeights_38 = weightsRAM_out[311:304]; // @[DenseLayer.scala 100:42]
  assign currWeights_39 = weightsRAM_out[319:312]; // @[DenseLayer.scala 100:42]
  assign currWeights_40 = weightsRAM_out[327:320]; // @[DenseLayer.scala 100:42]
  assign currWeights_41 = weightsRAM_out[335:328]; // @[DenseLayer.scala 100:42]
  assign currWeights_42 = weightsRAM_out[343:336]; // @[DenseLayer.scala 100:42]
  assign currWeights_43 = weightsRAM_out[351:344]; // @[DenseLayer.scala 100:42]
  assign currWeights_44 = weightsRAM_out[359:352]; // @[DenseLayer.scala 100:42]
  assign currWeights_45 = weightsRAM_out[367:360]; // @[DenseLayer.scala 100:42]
  assign currWeights_46 = weightsRAM_out[375:368]; // @[DenseLayer.scala 100:42]
  assign currWeights_47 = weightsRAM_out[383:376]; // @[DenseLayer.scala 100:42]
  assign currWeights_48 = weightsRAM_out[391:384]; // @[DenseLayer.scala 100:42]
  assign currWeights_49 = weightsRAM_out[399:392]; // @[DenseLayer.scala 100:42]
  assign currWeights_50 = weightsRAM_out[407:400]; // @[DenseLayer.scala 100:42]
  assign currWeights_51 = weightsRAM_out[415:408]; // @[DenseLayer.scala 100:42]
  assign currWeights_52 = weightsRAM_out[423:416]; // @[DenseLayer.scala 100:42]
  assign currWeights_53 = weightsRAM_out[431:424]; // @[DenseLayer.scala 100:42]
  assign currWeights_54 = weightsRAM_out[439:432]; // @[DenseLayer.scala 100:42]
  assign currWeights_55 = weightsRAM_out[447:440]; // @[DenseLayer.scala 100:42]
  assign currWeights_56 = weightsRAM_out[455:448]; // @[DenseLayer.scala 100:42]
  assign currWeights_57 = weightsRAM_out[463:456]; // @[DenseLayer.scala 100:42]
  assign currWeights_58 = weightsRAM_out[471:464]; // @[DenseLayer.scala 100:42]
  assign currWeights_59 = weightsRAM_out[479:472]; // @[DenseLayer.scala 100:42]
  assign currWeights_60 = weightsRAM_out[487:480]; // @[DenseLayer.scala 100:42]
  assign currWeights_61 = weightsRAM_out[495:488]; // @[DenseLayer.scala 100:42]
  assign currWeights_62 = weightsRAM_out[503:496]; // @[DenseLayer.scala 100:42]
  assign currWeights_63 = weightsRAM_out[511:504]; // @[DenseLayer.scala 100:42]
  assign currWeights_64 = weightsRAM_out[519:512]; // @[DenseLayer.scala 100:42]
  assign currWeights_65 = weightsRAM_out[527:520]; // @[DenseLayer.scala 100:42]
  assign currWeights_66 = weightsRAM_out[535:528]; // @[DenseLayer.scala 100:42]
  assign currWeights_67 = weightsRAM_out[543:536]; // @[DenseLayer.scala 100:42]
  assign currWeights_68 = weightsRAM_out[551:544]; // @[DenseLayer.scala 100:42]
  assign currWeights_69 = weightsRAM_out[559:552]; // @[DenseLayer.scala 100:42]
  assign currWeights_70 = weightsRAM_out[567:560]; // @[DenseLayer.scala 100:42]
  assign currWeights_71 = weightsRAM_out[575:568]; // @[DenseLayer.scala 100:42]
  assign currWeights_72 = weightsRAM_out[583:576]; // @[DenseLayer.scala 100:42]
  assign currWeights_73 = weightsRAM_out[591:584]; // @[DenseLayer.scala 100:42]
  assign currWeights_74 = weightsRAM_out[599:592]; // @[DenseLayer.scala 100:42]
  assign currWeights_75 = weightsRAM_out[607:600]; // @[DenseLayer.scala 100:42]
  assign currWeights_76 = weightsRAM_out[615:608]; // @[DenseLayer.scala 100:42]
  assign currWeights_77 = weightsRAM_out[623:616]; // @[DenseLayer.scala 100:42]
  assign currWeights_78 = weightsRAM_out[631:624]; // @[DenseLayer.scala 100:42]
  assign currWeights_79 = weightsRAM_out[639:632]; // @[DenseLayer.scala 100:42]
  assign currWeights_80 = weightsRAM_out[647:640]; // @[DenseLayer.scala 100:42]
  assign currWeights_81 = weightsRAM_out[655:648]; // @[DenseLayer.scala 100:42]
  assign currWeights_82 = weightsRAM_out[663:656]; // @[DenseLayer.scala 100:42]
  assign currWeights_83 = weightsRAM_out[671:664]; // @[DenseLayer.scala 100:42]
  assign currWeights_84 = weightsRAM_out[679:672]; // @[DenseLayer.scala 100:42]
  assign currWeights_85 = weightsRAM_out[687:680]; // @[DenseLayer.scala 100:42]
  assign currWeights_86 = weightsRAM_out[695:688]; // @[DenseLayer.scala 100:42]
  assign currWeights_87 = weightsRAM_out[703:696]; // @[DenseLayer.scala 100:42]
  assign currWeights_88 = weightsRAM_out[711:704]; // @[DenseLayer.scala 100:42]
  assign currWeights_89 = weightsRAM_out[719:712]; // @[DenseLayer.scala 100:42]
  assign currWeights_90 = weightsRAM_out[727:720]; // @[DenseLayer.scala 100:42]
  assign currWeights_91 = weightsRAM_out[735:728]; // @[DenseLayer.scala 100:42]
  assign currWeights_92 = weightsRAM_out[743:736]; // @[DenseLayer.scala 100:42]
  assign currWeights_93 = weightsRAM_out[751:744]; // @[DenseLayer.scala 100:42]
  assign currWeights_94 = weightsRAM_out[759:752]; // @[DenseLayer.scala 100:42]
  assign currWeights_95 = weightsRAM_out[767:760]; // @[DenseLayer.scala 100:42]
  assign currWeights_96 = weightsRAM_out[775:768]; // @[DenseLayer.scala 100:42]
  assign currWeights_97 = weightsRAM_out[783:776]; // @[DenseLayer.scala 100:42]
  assign currWeights_98 = weightsRAM_out[791:784]; // @[DenseLayer.scala 100:42]
  assign currWeights_99 = weightsRAM_out[799:792]; // @[DenseLayer.scala 100:42]
  assign currWeights_100 = weightsRAM_out[807:800]; // @[DenseLayer.scala 100:42]
  assign currWeights_101 = weightsRAM_out[815:808]; // @[DenseLayer.scala 100:42]
  assign currWeights_102 = weightsRAM_out[823:816]; // @[DenseLayer.scala 100:42]
  assign currWeights_103 = weightsRAM_out[831:824]; // @[DenseLayer.scala 100:42]
  assign currWeights_104 = weightsRAM_out[839:832]; // @[DenseLayer.scala 100:42]
  assign currWeights_105 = weightsRAM_out[847:840]; // @[DenseLayer.scala 100:42]
  assign currWeights_106 = weightsRAM_out[855:848]; // @[DenseLayer.scala 100:42]
  assign currWeights_107 = weightsRAM_out[863:856]; // @[DenseLayer.scala 100:42]
  assign currWeights_108 = weightsRAM_out[871:864]; // @[DenseLayer.scala 100:42]
  assign currWeights_109 = weightsRAM_out[879:872]; // @[DenseLayer.scala 100:42]
  assign currWeights_110 = weightsRAM_out[887:880]; // @[DenseLayer.scala 100:42]
  assign currWeights_111 = weightsRAM_out[895:888]; // @[DenseLayer.scala 100:42]
  assign currWeights_112 = weightsRAM_out[903:896]; // @[DenseLayer.scala 100:42]
  assign currWeights_113 = weightsRAM_out[911:904]; // @[DenseLayer.scala 100:42]
  assign currWeights_114 = weightsRAM_out[919:912]; // @[DenseLayer.scala 100:42]
  assign currWeights_115 = weightsRAM_out[927:920]; // @[DenseLayer.scala 100:42]
  assign currWeights_116 = weightsRAM_out[935:928]; // @[DenseLayer.scala 100:42]
  assign currWeights_117 = weightsRAM_out[943:936]; // @[DenseLayer.scala 100:42]
  assign currWeights_118 = weightsRAM_out[951:944]; // @[DenseLayer.scala 100:42]
  assign currWeights_119 = weightsRAM_out[959:952]; // @[DenseLayer.scala 100:42]
  assign currWeights_120 = weightsRAM_out[967:960]; // @[DenseLayer.scala 100:42]
  assign currWeights_121 = weightsRAM_out[975:968]; // @[DenseLayer.scala 100:42]
  assign currWeights_122 = weightsRAM_out[983:976]; // @[DenseLayer.scala 100:42]
  assign currWeights_123 = weightsRAM_out[991:984]; // @[DenseLayer.scala 100:42]
  assign currWeights_124 = weightsRAM_out[999:992]; // @[DenseLayer.scala 100:42]
  assign currWeights_125 = weightsRAM_out[1007:1000]; // @[DenseLayer.scala 100:42]
  assign currWeights_126 = weightsRAM_out[1015:1008]; // @[DenseLayer.scala 100:42]
  assign currWeights_127 = weightsRAM_out[1023:1016]; // @[DenseLayer.scala 100:42]
  assign _T_2398 = cntr == 10'h0; // @[DenseLayer.scala 121:33]
  assign _T_2416 = cntr == 10'h3ff; // @[DenseLayer.scala 123:16]
  assign _GEN_264 = _T_2416 ? 1'h1 : done; // @[DenseLayer.scala 123:42]
  assign _T_2418 = rst & done; // @[DenseLayer.scala 126:14]
  assign _GEN_265 = _T_2418 ? 1'h0 : _GEN_264; // @[DenseLayer.scala 126:23]
  assign _T_2434 = $signed(cummulativeSums_0) + $signed(MultiplyAccumulate_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2435 = _T_2434[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2436 = $signed(_T_2435); // @[DenseLayer.scala 133:59]
  assign _GEN_273 = vld ? $signed(_T_2436) : $signed(cummulativeSums_0); // @[DenseLayer.scala 132:18]
  assign _GEN_274 = rst ? $signed(16'sh0) : $signed(_GEN_273); // @[DenseLayer.scala 135:18]
  assign _T_2438 = rst & vld; // @[DenseLayer.scala 138:16]
  assign _GEN_275 = _T_2438 ? $signed(MultiplyAccumulate_io_sum) : $signed(_GEN_274); // @[DenseLayer.scala 138:24]
  assign _T_2439 = $signed(cummulativeSums_1) + $signed(MultiplyAccumulate_1_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2440 = _T_2439[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2441 = $signed(_T_2440); // @[DenseLayer.scala 133:59]
  assign _GEN_276 = vld ? $signed(_T_2441) : $signed(cummulativeSums_1); // @[DenseLayer.scala 132:18]
  assign _GEN_277 = rst ? $signed(16'sh0) : $signed(_GEN_276); // @[DenseLayer.scala 135:18]
  assign _GEN_278 = _T_2438 ? $signed(MultiplyAccumulate_1_io_sum) : $signed(_GEN_277); // @[DenseLayer.scala 138:24]
  assign _T_2444 = $signed(cummulativeSums_2) + $signed(MultiplyAccumulate_2_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2445 = _T_2444[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2446 = $signed(_T_2445); // @[DenseLayer.scala 133:59]
  assign _GEN_279 = vld ? $signed(_T_2446) : $signed(cummulativeSums_2); // @[DenseLayer.scala 132:18]
  assign _GEN_280 = rst ? $signed(16'sh0) : $signed(_GEN_279); // @[DenseLayer.scala 135:18]
  assign _GEN_281 = _T_2438 ? $signed(MultiplyAccumulate_2_io_sum) : $signed(_GEN_280); // @[DenseLayer.scala 138:24]
  assign _T_2449 = $signed(cummulativeSums_3) + $signed(MultiplyAccumulate_3_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2450 = _T_2449[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2451 = $signed(_T_2450); // @[DenseLayer.scala 133:59]
  assign _GEN_282 = vld ? $signed(_T_2451) : $signed(cummulativeSums_3); // @[DenseLayer.scala 132:18]
  assign _GEN_283 = rst ? $signed(16'sh0) : $signed(_GEN_282); // @[DenseLayer.scala 135:18]
  assign _GEN_284 = _T_2438 ? $signed(MultiplyAccumulate_3_io_sum) : $signed(_GEN_283); // @[DenseLayer.scala 138:24]
  assign _T_2454 = $signed(cummulativeSums_4) + $signed(MultiplyAccumulate_4_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2455 = _T_2454[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2456 = $signed(_T_2455); // @[DenseLayer.scala 133:59]
  assign _GEN_285 = vld ? $signed(_T_2456) : $signed(cummulativeSums_4); // @[DenseLayer.scala 132:18]
  assign _GEN_286 = rst ? $signed(16'sh0) : $signed(_GEN_285); // @[DenseLayer.scala 135:18]
  assign _GEN_287 = _T_2438 ? $signed(MultiplyAccumulate_4_io_sum) : $signed(_GEN_286); // @[DenseLayer.scala 138:24]
  assign _T_2459 = $signed(cummulativeSums_5) + $signed(MultiplyAccumulate_5_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2460 = _T_2459[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2461 = $signed(_T_2460); // @[DenseLayer.scala 133:59]
  assign _GEN_288 = vld ? $signed(_T_2461) : $signed(cummulativeSums_5); // @[DenseLayer.scala 132:18]
  assign _GEN_289 = rst ? $signed(16'sh0) : $signed(_GEN_288); // @[DenseLayer.scala 135:18]
  assign _GEN_290 = _T_2438 ? $signed(MultiplyAccumulate_5_io_sum) : $signed(_GEN_289); // @[DenseLayer.scala 138:24]
  assign _T_2464 = $signed(cummulativeSums_6) + $signed(MultiplyAccumulate_6_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2465 = _T_2464[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2466 = $signed(_T_2465); // @[DenseLayer.scala 133:59]
  assign _GEN_291 = vld ? $signed(_T_2466) : $signed(cummulativeSums_6); // @[DenseLayer.scala 132:18]
  assign _GEN_292 = rst ? $signed(16'sh0) : $signed(_GEN_291); // @[DenseLayer.scala 135:18]
  assign _GEN_293 = _T_2438 ? $signed(MultiplyAccumulate_6_io_sum) : $signed(_GEN_292); // @[DenseLayer.scala 138:24]
  assign _T_2469 = $signed(cummulativeSums_7) + $signed(MultiplyAccumulate_7_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2470 = _T_2469[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2471 = $signed(_T_2470); // @[DenseLayer.scala 133:59]
  assign _GEN_294 = vld ? $signed(_T_2471) : $signed(cummulativeSums_7); // @[DenseLayer.scala 132:18]
  assign _GEN_295 = rst ? $signed(16'sh0) : $signed(_GEN_294); // @[DenseLayer.scala 135:18]
  assign _GEN_296 = _T_2438 ? $signed(MultiplyAccumulate_7_io_sum) : $signed(_GEN_295); // @[DenseLayer.scala 138:24]
  assign _T_2474 = $signed(cummulativeSums_8) + $signed(MultiplyAccumulate_8_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2475 = _T_2474[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2476 = $signed(_T_2475); // @[DenseLayer.scala 133:59]
  assign _GEN_297 = vld ? $signed(_T_2476) : $signed(cummulativeSums_8); // @[DenseLayer.scala 132:18]
  assign _GEN_298 = rst ? $signed(16'sh0) : $signed(_GEN_297); // @[DenseLayer.scala 135:18]
  assign _GEN_299 = _T_2438 ? $signed(MultiplyAccumulate_8_io_sum) : $signed(_GEN_298); // @[DenseLayer.scala 138:24]
  assign _T_2479 = $signed(cummulativeSums_9) + $signed(MultiplyAccumulate_9_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2480 = _T_2479[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2481 = $signed(_T_2480); // @[DenseLayer.scala 133:59]
  assign _GEN_300 = vld ? $signed(_T_2481) : $signed(cummulativeSums_9); // @[DenseLayer.scala 132:18]
  assign _GEN_301 = rst ? $signed(16'sh0) : $signed(_GEN_300); // @[DenseLayer.scala 135:18]
  assign _GEN_302 = _T_2438 ? $signed(MultiplyAccumulate_9_io_sum) : $signed(_GEN_301); // @[DenseLayer.scala 138:24]
  assign _T_2484 = $signed(cummulativeSums_10) + $signed(MultiplyAccumulate_10_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2485 = _T_2484[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2486 = $signed(_T_2485); // @[DenseLayer.scala 133:59]
  assign _GEN_303 = vld ? $signed(_T_2486) : $signed(cummulativeSums_10); // @[DenseLayer.scala 132:18]
  assign _GEN_304 = rst ? $signed(16'sh0) : $signed(_GEN_303); // @[DenseLayer.scala 135:18]
  assign _GEN_305 = _T_2438 ? $signed(MultiplyAccumulate_10_io_sum) : $signed(_GEN_304); // @[DenseLayer.scala 138:24]
  assign _T_2489 = $signed(cummulativeSums_11) + $signed(MultiplyAccumulate_11_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2490 = _T_2489[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2491 = $signed(_T_2490); // @[DenseLayer.scala 133:59]
  assign _GEN_306 = vld ? $signed(_T_2491) : $signed(cummulativeSums_11); // @[DenseLayer.scala 132:18]
  assign _GEN_307 = rst ? $signed(16'sh0) : $signed(_GEN_306); // @[DenseLayer.scala 135:18]
  assign _GEN_308 = _T_2438 ? $signed(MultiplyAccumulate_11_io_sum) : $signed(_GEN_307); // @[DenseLayer.scala 138:24]
  assign _T_2494 = $signed(cummulativeSums_12) + $signed(MultiplyAccumulate_12_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2495 = _T_2494[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2496 = $signed(_T_2495); // @[DenseLayer.scala 133:59]
  assign _GEN_309 = vld ? $signed(_T_2496) : $signed(cummulativeSums_12); // @[DenseLayer.scala 132:18]
  assign _GEN_310 = rst ? $signed(16'sh0) : $signed(_GEN_309); // @[DenseLayer.scala 135:18]
  assign _GEN_311 = _T_2438 ? $signed(MultiplyAccumulate_12_io_sum) : $signed(_GEN_310); // @[DenseLayer.scala 138:24]
  assign _T_2499 = $signed(cummulativeSums_13) + $signed(MultiplyAccumulate_13_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2500 = _T_2499[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2501 = $signed(_T_2500); // @[DenseLayer.scala 133:59]
  assign _GEN_312 = vld ? $signed(_T_2501) : $signed(cummulativeSums_13); // @[DenseLayer.scala 132:18]
  assign _GEN_313 = rst ? $signed(16'sh0) : $signed(_GEN_312); // @[DenseLayer.scala 135:18]
  assign _GEN_314 = _T_2438 ? $signed(MultiplyAccumulate_13_io_sum) : $signed(_GEN_313); // @[DenseLayer.scala 138:24]
  assign _T_2504 = $signed(cummulativeSums_14) + $signed(MultiplyAccumulate_14_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2505 = _T_2504[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2506 = $signed(_T_2505); // @[DenseLayer.scala 133:59]
  assign _GEN_315 = vld ? $signed(_T_2506) : $signed(cummulativeSums_14); // @[DenseLayer.scala 132:18]
  assign _GEN_316 = rst ? $signed(16'sh0) : $signed(_GEN_315); // @[DenseLayer.scala 135:18]
  assign _GEN_317 = _T_2438 ? $signed(MultiplyAccumulate_14_io_sum) : $signed(_GEN_316); // @[DenseLayer.scala 138:24]
  assign _T_2509 = $signed(cummulativeSums_15) + $signed(MultiplyAccumulate_15_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2510 = _T_2509[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2511 = $signed(_T_2510); // @[DenseLayer.scala 133:59]
  assign _GEN_318 = vld ? $signed(_T_2511) : $signed(cummulativeSums_15); // @[DenseLayer.scala 132:18]
  assign _GEN_319 = rst ? $signed(16'sh0) : $signed(_GEN_318); // @[DenseLayer.scala 135:18]
  assign _GEN_320 = _T_2438 ? $signed(MultiplyAccumulate_15_io_sum) : $signed(_GEN_319); // @[DenseLayer.scala 138:24]
  assign _T_2514 = $signed(cummulativeSums_16) + $signed(MultiplyAccumulate_16_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2515 = _T_2514[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2516 = $signed(_T_2515); // @[DenseLayer.scala 133:59]
  assign _GEN_321 = vld ? $signed(_T_2516) : $signed(cummulativeSums_16); // @[DenseLayer.scala 132:18]
  assign _GEN_322 = rst ? $signed(16'sh0) : $signed(_GEN_321); // @[DenseLayer.scala 135:18]
  assign _GEN_323 = _T_2438 ? $signed(MultiplyAccumulate_16_io_sum) : $signed(_GEN_322); // @[DenseLayer.scala 138:24]
  assign _T_2519 = $signed(cummulativeSums_17) + $signed(MultiplyAccumulate_17_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2520 = _T_2519[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2521 = $signed(_T_2520); // @[DenseLayer.scala 133:59]
  assign _GEN_324 = vld ? $signed(_T_2521) : $signed(cummulativeSums_17); // @[DenseLayer.scala 132:18]
  assign _GEN_325 = rst ? $signed(16'sh0) : $signed(_GEN_324); // @[DenseLayer.scala 135:18]
  assign _GEN_326 = _T_2438 ? $signed(MultiplyAccumulate_17_io_sum) : $signed(_GEN_325); // @[DenseLayer.scala 138:24]
  assign _T_2524 = $signed(cummulativeSums_18) + $signed(MultiplyAccumulate_18_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2525 = _T_2524[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2526 = $signed(_T_2525); // @[DenseLayer.scala 133:59]
  assign _GEN_327 = vld ? $signed(_T_2526) : $signed(cummulativeSums_18); // @[DenseLayer.scala 132:18]
  assign _GEN_328 = rst ? $signed(16'sh0) : $signed(_GEN_327); // @[DenseLayer.scala 135:18]
  assign _GEN_329 = _T_2438 ? $signed(MultiplyAccumulate_18_io_sum) : $signed(_GEN_328); // @[DenseLayer.scala 138:24]
  assign _T_2529 = $signed(cummulativeSums_19) + $signed(MultiplyAccumulate_19_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2530 = _T_2529[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2531 = $signed(_T_2530); // @[DenseLayer.scala 133:59]
  assign _GEN_330 = vld ? $signed(_T_2531) : $signed(cummulativeSums_19); // @[DenseLayer.scala 132:18]
  assign _GEN_331 = rst ? $signed(16'sh0) : $signed(_GEN_330); // @[DenseLayer.scala 135:18]
  assign _GEN_332 = _T_2438 ? $signed(MultiplyAccumulate_19_io_sum) : $signed(_GEN_331); // @[DenseLayer.scala 138:24]
  assign _T_2534 = $signed(cummulativeSums_20) + $signed(MultiplyAccumulate_20_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2535 = _T_2534[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2536 = $signed(_T_2535); // @[DenseLayer.scala 133:59]
  assign _GEN_333 = vld ? $signed(_T_2536) : $signed(cummulativeSums_20); // @[DenseLayer.scala 132:18]
  assign _GEN_334 = rst ? $signed(16'sh0) : $signed(_GEN_333); // @[DenseLayer.scala 135:18]
  assign _GEN_335 = _T_2438 ? $signed(MultiplyAccumulate_20_io_sum) : $signed(_GEN_334); // @[DenseLayer.scala 138:24]
  assign _T_2539 = $signed(cummulativeSums_21) + $signed(MultiplyAccumulate_21_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2540 = _T_2539[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2541 = $signed(_T_2540); // @[DenseLayer.scala 133:59]
  assign _GEN_336 = vld ? $signed(_T_2541) : $signed(cummulativeSums_21); // @[DenseLayer.scala 132:18]
  assign _GEN_337 = rst ? $signed(16'sh0) : $signed(_GEN_336); // @[DenseLayer.scala 135:18]
  assign _GEN_338 = _T_2438 ? $signed(MultiplyAccumulate_21_io_sum) : $signed(_GEN_337); // @[DenseLayer.scala 138:24]
  assign _T_2544 = $signed(cummulativeSums_22) + $signed(MultiplyAccumulate_22_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2545 = _T_2544[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2546 = $signed(_T_2545); // @[DenseLayer.scala 133:59]
  assign _GEN_339 = vld ? $signed(_T_2546) : $signed(cummulativeSums_22); // @[DenseLayer.scala 132:18]
  assign _GEN_340 = rst ? $signed(16'sh0) : $signed(_GEN_339); // @[DenseLayer.scala 135:18]
  assign _GEN_341 = _T_2438 ? $signed(MultiplyAccumulate_22_io_sum) : $signed(_GEN_340); // @[DenseLayer.scala 138:24]
  assign _T_2549 = $signed(cummulativeSums_23) + $signed(MultiplyAccumulate_23_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2550 = _T_2549[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2551 = $signed(_T_2550); // @[DenseLayer.scala 133:59]
  assign _GEN_342 = vld ? $signed(_T_2551) : $signed(cummulativeSums_23); // @[DenseLayer.scala 132:18]
  assign _GEN_343 = rst ? $signed(16'sh0) : $signed(_GEN_342); // @[DenseLayer.scala 135:18]
  assign _GEN_344 = _T_2438 ? $signed(MultiplyAccumulate_23_io_sum) : $signed(_GEN_343); // @[DenseLayer.scala 138:24]
  assign _T_2554 = $signed(cummulativeSums_24) + $signed(MultiplyAccumulate_24_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2555 = _T_2554[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2556 = $signed(_T_2555); // @[DenseLayer.scala 133:59]
  assign _GEN_345 = vld ? $signed(_T_2556) : $signed(cummulativeSums_24); // @[DenseLayer.scala 132:18]
  assign _GEN_346 = rst ? $signed(16'sh0) : $signed(_GEN_345); // @[DenseLayer.scala 135:18]
  assign _GEN_347 = _T_2438 ? $signed(MultiplyAccumulate_24_io_sum) : $signed(_GEN_346); // @[DenseLayer.scala 138:24]
  assign _T_2559 = $signed(cummulativeSums_25) + $signed(MultiplyAccumulate_25_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2560 = _T_2559[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2561 = $signed(_T_2560); // @[DenseLayer.scala 133:59]
  assign _GEN_348 = vld ? $signed(_T_2561) : $signed(cummulativeSums_25); // @[DenseLayer.scala 132:18]
  assign _GEN_349 = rst ? $signed(16'sh0) : $signed(_GEN_348); // @[DenseLayer.scala 135:18]
  assign _GEN_350 = _T_2438 ? $signed(MultiplyAccumulate_25_io_sum) : $signed(_GEN_349); // @[DenseLayer.scala 138:24]
  assign _T_2564 = $signed(cummulativeSums_26) + $signed(MultiplyAccumulate_26_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2565 = _T_2564[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2566 = $signed(_T_2565); // @[DenseLayer.scala 133:59]
  assign _GEN_351 = vld ? $signed(_T_2566) : $signed(cummulativeSums_26); // @[DenseLayer.scala 132:18]
  assign _GEN_352 = rst ? $signed(16'sh0) : $signed(_GEN_351); // @[DenseLayer.scala 135:18]
  assign _GEN_353 = _T_2438 ? $signed(MultiplyAccumulate_26_io_sum) : $signed(_GEN_352); // @[DenseLayer.scala 138:24]
  assign _T_2569 = $signed(cummulativeSums_27) + $signed(MultiplyAccumulate_27_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2570 = _T_2569[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2571 = $signed(_T_2570); // @[DenseLayer.scala 133:59]
  assign _GEN_354 = vld ? $signed(_T_2571) : $signed(cummulativeSums_27); // @[DenseLayer.scala 132:18]
  assign _GEN_355 = rst ? $signed(16'sh0) : $signed(_GEN_354); // @[DenseLayer.scala 135:18]
  assign _GEN_356 = _T_2438 ? $signed(MultiplyAccumulate_27_io_sum) : $signed(_GEN_355); // @[DenseLayer.scala 138:24]
  assign _T_2574 = $signed(cummulativeSums_28) + $signed(MultiplyAccumulate_28_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2575 = _T_2574[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2576 = $signed(_T_2575); // @[DenseLayer.scala 133:59]
  assign _GEN_357 = vld ? $signed(_T_2576) : $signed(cummulativeSums_28); // @[DenseLayer.scala 132:18]
  assign _GEN_358 = rst ? $signed(16'sh0) : $signed(_GEN_357); // @[DenseLayer.scala 135:18]
  assign _GEN_359 = _T_2438 ? $signed(MultiplyAccumulate_28_io_sum) : $signed(_GEN_358); // @[DenseLayer.scala 138:24]
  assign _T_2579 = $signed(cummulativeSums_29) + $signed(MultiplyAccumulate_29_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2580 = _T_2579[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2581 = $signed(_T_2580); // @[DenseLayer.scala 133:59]
  assign _GEN_360 = vld ? $signed(_T_2581) : $signed(cummulativeSums_29); // @[DenseLayer.scala 132:18]
  assign _GEN_361 = rst ? $signed(16'sh0) : $signed(_GEN_360); // @[DenseLayer.scala 135:18]
  assign _GEN_362 = _T_2438 ? $signed(MultiplyAccumulate_29_io_sum) : $signed(_GEN_361); // @[DenseLayer.scala 138:24]
  assign _T_2584 = $signed(cummulativeSums_30) + $signed(MultiplyAccumulate_30_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2585 = _T_2584[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2586 = $signed(_T_2585); // @[DenseLayer.scala 133:59]
  assign _GEN_363 = vld ? $signed(_T_2586) : $signed(cummulativeSums_30); // @[DenseLayer.scala 132:18]
  assign _GEN_364 = rst ? $signed(16'sh0) : $signed(_GEN_363); // @[DenseLayer.scala 135:18]
  assign _GEN_365 = _T_2438 ? $signed(MultiplyAccumulate_30_io_sum) : $signed(_GEN_364); // @[DenseLayer.scala 138:24]
  assign _T_2589 = $signed(cummulativeSums_31) + $signed(MultiplyAccumulate_31_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2590 = _T_2589[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2591 = $signed(_T_2590); // @[DenseLayer.scala 133:59]
  assign _GEN_366 = vld ? $signed(_T_2591) : $signed(cummulativeSums_31); // @[DenseLayer.scala 132:18]
  assign _GEN_367 = rst ? $signed(16'sh0) : $signed(_GEN_366); // @[DenseLayer.scala 135:18]
  assign _GEN_368 = _T_2438 ? $signed(MultiplyAccumulate_31_io_sum) : $signed(_GEN_367); // @[DenseLayer.scala 138:24]
  assign _T_2594 = $signed(cummulativeSums_32) + $signed(MultiplyAccumulate_32_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2595 = _T_2594[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2596 = $signed(_T_2595); // @[DenseLayer.scala 133:59]
  assign _GEN_369 = vld ? $signed(_T_2596) : $signed(cummulativeSums_32); // @[DenseLayer.scala 132:18]
  assign _GEN_370 = rst ? $signed(16'sh0) : $signed(_GEN_369); // @[DenseLayer.scala 135:18]
  assign _GEN_371 = _T_2438 ? $signed(MultiplyAccumulate_32_io_sum) : $signed(_GEN_370); // @[DenseLayer.scala 138:24]
  assign _T_2599 = $signed(cummulativeSums_33) + $signed(MultiplyAccumulate_33_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2600 = _T_2599[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2601 = $signed(_T_2600); // @[DenseLayer.scala 133:59]
  assign _GEN_372 = vld ? $signed(_T_2601) : $signed(cummulativeSums_33); // @[DenseLayer.scala 132:18]
  assign _GEN_373 = rst ? $signed(16'sh0) : $signed(_GEN_372); // @[DenseLayer.scala 135:18]
  assign _GEN_374 = _T_2438 ? $signed(MultiplyAccumulate_33_io_sum) : $signed(_GEN_373); // @[DenseLayer.scala 138:24]
  assign _T_2604 = $signed(cummulativeSums_34) + $signed(MultiplyAccumulate_34_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2605 = _T_2604[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2606 = $signed(_T_2605); // @[DenseLayer.scala 133:59]
  assign _GEN_375 = vld ? $signed(_T_2606) : $signed(cummulativeSums_34); // @[DenseLayer.scala 132:18]
  assign _GEN_376 = rst ? $signed(16'sh0) : $signed(_GEN_375); // @[DenseLayer.scala 135:18]
  assign _GEN_377 = _T_2438 ? $signed(MultiplyAccumulate_34_io_sum) : $signed(_GEN_376); // @[DenseLayer.scala 138:24]
  assign _T_2609 = $signed(cummulativeSums_35) + $signed(MultiplyAccumulate_35_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2610 = _T_2609[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2611 = $signed(_T_2610); // @[DenseLayer.scala 133:59]
  assign _GEN_378 = vld ? $signed(_T_2611) : $signed(cummulativeSums_35); // @[DenseLayer.scala 132:18]
  assign _GEN_379 = rst ? $signed(16'sh0) : $signed(_GEN_378); // @[DenseLayer.scala 135:18]
  assign _GEN_380 = _T_2438 ? $signed(MultiplyAccumulate_35_io_sum) : $signed(_GEN_379); // @[DenseLayer.scala 138:24]
  assign _T_2614 = $signed(cummulativeSums_36) + $signed(MultiplyAccumulate_36_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2615 = _T_2614[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2616 = $signed(_T_2615); // @[DenseLayer.scala 133:59]
  assign _GEN_381 = vld ? $signed(_T_2616) : $signed(cummulativeSums_36); // @[DenseLayer.scala 132:18]
  assign _GEN_382 = rst ? $signed(16'sh0) : $signed(_GEN_381); // @[DenseLayer.scala 135:18]
  assign _GEN_383 = _T_2438 ? $signed(MultiplyAccumulate_36_io_sum) : $signed(_GEN_382); // @[DenseLayer.scala 138:24]
  assign _T_2619 = $signed(cummulativeSums_37) + $signed(MultiplyAccumulate_37_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2620 = _T_2619[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2621 = $signed(_T_2620); // @[DenseLayer.scala 133:59]
  assign _GEN_384 = vld ? $signed(_T_2621) : $signed(cummulativeSums_37); // @[DenseLayer.scala 132:18]
  assign _GEN_385 = rst ? $signed(16'sh0) : $signed(_GEN_384); // @[DenseLayer.scala 135:18]
  assign _GEN_386 = _T_2438 ? $signed(MultiplyAccumulate_37_io_sum) : $signed(_GEN_385); // @[DenseLayer.scala 138:24]
  assign _T_2624 = $signed(cummulativeSums_38) + $signed(MultiplyAccumulate_38_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2625 = _T_2624[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2626 = $signed(_T_2625); // @[DenseLayer.scala 133:59]
  assign _GEN_387 = vld ? $signed(_T_2626) : $signed(cummulativeSums_38); // @[DenseLayer.scala 132:18]
  assign _GEN_388 = rst ? $signed(16'sh0) : $signed(_GEN_387); // @[DenseLayer.scala 135:18]
  assign _GEN_389 = _T_2438 ? $signed(MultiplyAccumulate_38_io_sum) : $signed(_GEN_388); // @[DenseLayer.scala 138:24]
  assign _T_2629 = $signed(cummulativeSums_39) + $signed(MultiplyAccumulate_39_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2630 = _T_2629[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2631 = $signed(_T_2630); // @[DenseLayer.scala 133:59]
  assign _GEN_390 = vld ? $signed(_T_2631) : $signed(cummulativeSums_39); // @[DenseLayer.scala 132:18]
  assign _GEN_391 = rst ? $signed(16'sh0) : $signed(_GEN_390); // @[DenseLayer.scala 135:18]
  assign _GEN_392 = _T_2438 ? $signed(MultiplyAccumulate_39_io_sum) : $signed(_GEN_391); // @[DenseLayer.scala 138:24]
  assign _T_2634 = $signed(cummulativeSums_40) + $signed(MultiplyAccumulate_40_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2635 = _T_2634[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2636 = $signed(_T_2635); // @[DenseLayer.scala 133:59]
  assign _GEN_393 = vld ? $signed(_T_2636) : $signed(cummulativeSums_40); // @[DenseLayer.scala 132:18]
  assign _GEN_394 = rst ? $signed(16'sh0) : $signed(_GEN_393); // @[DenseLayer.scala 135:18]
  assign _GEN_395 = _T_2438 ? $signed(MultiplyAccumulate_40_io_sum) : $signed(_GEN_394); // @[DenseLayer.scala 138:24]
  assign _T_2639 = $signed(cummulativeSums_41) + $signed(MultiplyAccumulate_41_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2640 = _T_2639[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2641 = $signed(_T_2640); // @[DenseLayer.scala 133:59]
  assign _GEN_396 = vld ? $signed(_T_2641) : $signed(cummulativeSums_41); // @[DenseLayer.scala 132:18]
  assign _GEN_397 = rst ? $signed(16'sh0) : $signed(_GEN_396); // @[DenseLayer.scala 135:18]
  assign _GEN_398 = _T_2438 ? $signed(MultiplyAccumulate_41_io_sum) : $signed(_GEN_397); // @[DenseLayer.scala 138:24]
  assign _T_2644 = $signed(cummulativeSums_42) + $signed(MultiplyAccumulate_42_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2645 = _T_2644[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2646 = $signed(_T_2645); // @[DenseLayer.scala 133:59]
  assign _GEN_399 = vld ? $signed(_T_2646) : $signed(cummulativeSums_42); // @[DenseLayer.scala 132:18]
  assign _GEN_400 = rst ? $signed(16'sh0) : $signed(_GEN_399); // @[DenseLayer.scala 135:18]
  assign _GEN_401 = _T_2438 ? $signed(MultiplyAccumulate_42_io_sum) : $signed(_GEN_400); // @[DenseLayer.scala 138:24]
  assign _T_2649 = $signed(cummulativeSums_43) + $signed(MultiplyAccumulate_43_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2650 = _T_2649[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2651 = $signed(_T_2650); // @[DenseLayer.scala 133:59]
  assign _GEN_402 = vld ? $signed(_T_2651) : $signed(cummulativeSums_43); // @[DenseLayer.scala 132:18]
  assign _GEN_403 = rst ? $signed(16'sh0) : $signed(_GEN_402); // @[DenseLayer.scala 135:18]
  assign _GEN_404 = _T_2438 ? $signed(MultiplyAccumulate_43_io_sum) : $signed(_GEN_403); // @[DenseLayer.scala 138:24]
  assign _T_2654 = $signed(cummulativeSums_44) + $signed(MultiplyAccumulate_44_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2655 = _T_2654[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2656 = $signed(_T_2655); // @[DenseLayer.scala 133:59]
  assign _GEN_405 = vld ? $signed(_T_2656) : $signed(cummulativeSums_44); // @[DenseLayer.scala 132:18]
  assign _GEN_406 = rst ? $signed(16'sh0) : $signed(_GEN_405); // @[DenseLayer.scala 135:18]
  assign _GEN_407 = _T_2438 ? $signed(MultiplyAccumulate_44_io_sum) : $signed(_GEN_406); // @[DenseLayer.scala 138:24]
  assign _T_2659 = $signed(cummulativeSums_45) + $signed(MultiplyAccumulate_45_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2660 = _T_2659[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2661 = $signed(_T_2660); // @[DenseLayer.scala 133:59]
  assign _GEN_408 = vld ? $signed(_T_2661) : $signed(cummulativeSums_45); // @[DenseLayer.scala 132:18]
  assign _GEN_409 = rst ? $signed(16'sh0) : $signed(_GEN_408); // @[DenseLayer.scala 135:18]
  assign _GEN_410 = _T_2438 ? $signed(MultiplyAccumulate_45_io_sum) : $signed(_GEN_409); // @[DenseLayer.scala 138:24]
  assign _T_2664 = $signed(cummulativeSums_46) + $signed(MultiplyAccumulate_46_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2665 = _T_2664[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2666 = $signed(_T_2665); // @[DenseLayer.scala 133:59]
  assign _GEN_411 = vld ? $signed(_T_2666) : $signed(cummulativeSums_46); // @[DenseLayer.scala 132:18]
  assign _GEN_412 = rst ? $signed(16'sh0) : $signed(_GEN_411); // @[DenseLayer.scala 135:18]
  assign _GEN_413 = _T_2438 ? $signed(MultiplyAccumulate_46_io_sum) : $signed(_GEN_412); // @[DenseLayer.scala 138:24]
  assign _T_2669 = $signed(cummulativeSums_47) + $signed(MultiplyAccumulate_47_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2670 = _T_2669[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2671 = $signed(_T_2670); // @[DenseLayer.scala 133:59]
  assign _GEN_414 = vld ? $signed(_T_2671) : $signed(cummulativeSums_47); // @[DenseLayer.scala 132:18]
  assign _GEN_415 = rst ? $signed(16'sh0) : $signed(_GEN_414); // @[DenseLayer.scala 135:18]
  assign _GEN_416 = _T_2438 ? $signed(MultiplyAccumulate_47_io_sum) : $signed(_GEN_415); // @[DenseLayer.scala 138:24]
  assign _T_2674 = $signed(cummulativeSums_48) + $signed(MultiplyAccumulate_48_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2675 = _T_2674[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2676 = $signed(_T_2675); // @[DenseLayer.scala 133:59]
  assign _GEN_417 = vld ? $signed(_T_2676) : $signed(cummulativeSums_48); // @[DenseLayer.scala 132:18]
  assign _GEN_418 = rst ? $signed(16'sh0) : $signed(_GEN_417); // @[DenseLayer.scala 135:18]
  assign _GEN_419 = _T_2438 ? $signed(MultiplyAccumulate_48_io_sum) : $signed(_GEN_418); // @[DenseLayer.scala 138:24]
  assign _T_2679 = $signed(cummulativeSums_49) + $signed(MultiplyAccumulate_49_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2680 = _T_2679[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2681 = $signed(_T_2680); // @[DenseLayer.scala 133:59]
  assign _GEN_420 = vld ? $signed(_T_2681) : $signed(cummulativeSums_49); // @[DenseLayer.scala 132:18]
  assign _GEN_421 = rst ? $signed(16'sh0) : $signed(_GEN_420); // @[DenseLayer.scala 135:18]
  assign _GEN_422 = _T_2438 ? $signed(MultiplyAccumulate_49_io_sum) : $signed(_GEN_421); // @[DenseLayer.scala 138:24]
  assign _T_2684 = $signed(cummulativeSums_50) + $signed(MultiplyAccumulate_50_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2685 = _T_2684[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2686 = $signed(_T_2685); // @[DenseLayer.scala 133:59]
  assign _GEN_423 = vld ? $signed(_T_2686) : $signed(cummulativeSums_50); // @[DenseLayer.scala 132:18]
  assign _GEN_424 = rst ? $signed(16'sh0) : $signed(_GEN_423); // @[DenseLayer.scala 135:18]
  assign _GEN_425 = _T_2438 ? $signed(MultiplyAccumulate_50_io_sum) : $signed(_GEN_424); // @[DenseLayer.scala 138:24]
  assign _T_2689 = $signed(cummulativeSums_51) + $signed(MultiplyAccumulate_51_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2690 = _T_2689[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2691 = $signed(_T_2690); // @[DenseLayer.scala 133:59]
  assign _GEN_426 = vld ? $signed(_T_2691) : $signed(cummulativeSums_51); // @[DenseLayer.scala 132:18]
  assign _GEN_427 = rst ? $signed(16'sh0) : $signed(_GEN_426); // @[DenseLayer.scala 135:18]
  assign _GEN_428 = _T_2438 ? $signed(MultiplyAccumulate_51_io_sum) : $signed(_GEN_427); // @[DenseLayer.scala 138:24]
  assign _T_2694 = $signed(cummulativeSums_52) + $signed(MultiplyAccumulate_52_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2695 = _T_2694[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2696 = $signed(_T_2695); // @[DenseLayer.scala 133:59]
  assign _GEN_429 = vld ? $signed(_T_2696) : $signed(cummulativeSums_52); // @[DenseLayer.scala 132:18]
  assign _GEN_430 = rst ? $signed(16'sh0) : $signed(_GEN_429); // @[DenseLayer.scala 135:18]
  assign _GEN_431 = _T_2438 ? $signed(MultiplyAccumulate_52_io_sum) : $signed(_GEN_430); // @[DenseLayer.scala 138:24]
  assign _T_2699 = $signed(cummulativeSums_53) + $signed(MultiplyAccumulate_53_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2700 = _T_2699[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2701 = $signed(_T_2700); // @[DenseLayer.scala 133:59]
  assign _GEN_432 = vld ? $signed(_T_2701) : $signed(cummulativeSums_53); // @[DenseLayer.scala 132:18]
  assign _GEN_433 = rst ? $signed(16'sh0) : $signed(_GEN_432); // @[DenseLayer.scala 135:18]
  assign _GEN_434 = _T_2438 ? $signed(MultiplyAccumulate_53_io_sum) : $signed(_GEN_433); // @[DenseLayer.scala 138:24]
  assign _T_2704 = $signed(cummulativeSums_54) + $signed(MultiplyAccumulate_54_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2705 = _T_2704[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2706 = $signed(_T_2705); // @[DenseLayer.scala 133:59]
  assign _GEN_435 = vld ? $signed(_T_2706) : $signed(cummulativeSums_54); // @[DenseLayer.scala 132:18]
  assign _GEN_436 = rst ? $signed(16'sh0) : $signed(_GEN_435); // @[DenseLayer.scala 135:18]
  assign _GEN_437 = _T_2438 ? $signed(MultiplyAccumulate_54_io_sum) : $signed(_GEN_436); // @[DenseLayer.scala 138:24]
  assign _T_2709 = $signed(cummulativeSums_55) + $signed(MultiplyAccumulate_55_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2710 = _T_2709[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2711 = $signed(_T_2710); // @[DenseLayer.scala 133:59]
  assign _GEN_438 = vld ? $signed(_T_2711) : $signed(cummulativeSums_55); // @[DenseLayer.scala 132:18]
  assign _GEN_439 = rst ? $signed(16'sh0) : $signed(_GEN_438); // @[DenseLayer.scala 135:18]
  assign _GEN_440 = _T_2438 ? $signed(MultiplyAccumulate_55_io_sum) : $signed(_GEN_439); // @[DenseLayer.scala 138:24]
  assign _T_2714 = $signed(cummulativeSums_56) + $signed(MultiplyAccumulate_56_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2715 = _T_2714[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2716 = $signed(_T_2715); // @[DenseLayer.scala 133:59]
  assign _GEN_441 = vld ? $signed(_T_2716) : $signed(cummulativeSums_56); // @[DenseLayer.scala 132:18]
  assign _GEN_442 = rst ? $signed(16'sh0) : $signed(_GEN_441); // @[DenseLayer.scala 135:18]
  assign _GEN_443 = _T_2438 ? $signed(MultiplyAccumulate_56_io_sum) : $signed(_GEN_442); // @[DenseLayer.scala 138:24]
  assign _T_2719 = $signed(cummulativeSums_57) + $signed(MultiplyAccumulate_57_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2720 = _T_2719[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2721 = $signed(_T_2720); // @[DenseLayer.scala 133:59]
  assign _GEN_444 = vld ? $signed(_T_2721) : $signed(cummulativeSums_57); // @[DenseLayer.scala 132:18]
  assign _GEN_445 = rst ? $signed(16'sh0) : $signed(_GEN_444); // @[DenseLayer.scala 135:18]
  assign _GEN_446 = _T_2438 ? $signed(MultiplyAccumulate_57_io_sum) : $signed(_GEN_445); // @[DenseLayer.scala 138:24]
  assign _T_2724 = $signed(cummulativeSums_58) + $signed(MultiplyAccumulate_58_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2725 = _T_2724[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2726 = $signed(_T_2725); // @[DenseLayer.scala 133:59]
  assign _GEN_447 = vld ? $signed(_T_2726) : $signed(cummulativeSums_58); // @[DenseLayer.scala 132:18]
  assign _GEN_448 = rst ? $signed(16'sh0) : $signed(_GEN_447); // @[DenseLayer.scala 135:18]
  assign _GEN_449 = _T_2438 ? $signed(MultiplyAccumulate_58_io_sum) : $signed(_GEN_448); // @[DenseLayer.scala 138:24]
  assign _T_2729 = $signed(cummulativeSums_59) + $signed(MultiplyAccumulate_59_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2730 = _T_2729[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2731 = $signed(_T_2730); // @[DenseLayer.scala 133:59]
  assign _GEN_450 = vld ? $signed(_T_2731) : $signed(cummulativeSums_59); // @[DenseLayer.scala 132:18]
  assign _GEN_451 = rst ? $signed(16'sh0) : $signed(_GEN_450); // @[DenseLayer.scala 135:18]
  assign _GEN_452 = _T_2438 ? $signed(MultiplyAccumulate_59_io_sum) : $signed(_GEN_451); // @[DenseLayer.scala 138:24]
  assign _T_2734 = $signed(cummulativeSums_60) + $signed(MultiplyAccumulate_60_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2735 = _T_2734[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2736 = $signed(_T_2735); // @[DenseLayer.scala 133:59]
  assign _GEN_453 = vld ? $signed(_T_2736) : $signed(cummulativeSums_60); // @[DenseLayer.scala 132:18]
  assign _GEN_454 = rst ? $signed(16'sh0) : $signed(_GEN_453); // @[DenseLayer.scala 135:18]
  assign _GEN_455 = _T_2438 ? $signed(MultiplyAccumulate_60_io_sum) : $signed(_GEN_454); // @[DenseLayer.scala 138:24]
  assign _T_2739 = $signed(cummulativeSums_61) + $signed(MultiplyAccumulate_61_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2740 = _T_2739[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2741 = $signed(_T_2740); // @[DenseLayer.scala 133:59]
  assign _GEN_456 = vld ? $signed(_T_2741) : $signed(cummulativeSums_61); // @[DenseLayer.scala 132:18]
  assign _GEN_457 = rst ? $signed(16'sh0) : $signed(_GEN_456); // @[DenseLayer.scala 135:18]
  assign _GEN_458 = _T_2438 ? $signed(MultiplyAccumulate_61_io_sum) : $signed(_GEN_457); // @[DenseLayer.scala 138:24]
  assign _T_2744 = $signed(cummulativeSums_62) + $signed(MultiplyAccumulate_62_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2745 = _T_2744[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2746 = $signed(_T_2745); // @[DenseLayer.scala 133:59]
  assign _GEN_459 = vld ? $signed(_T_2746) : $signed(cummulativeSums_62); // @[DenseLayer.scala 132:18]
  assign _GEN_460 = rst ? $signed(16'sh0) : $signed(_GEN_459); // @[DenseLayer.scala 135:18]
  assign _GEN_461 = _T_2438 ? $signed(MultiplyAccumulate_62_io_sum) : $signed(_GEN_460); // @[DenseLayer.scala 138:24]
  assign _T_2749 = $signed(cummulativeSums_63) + $signed(MultiplyAccumulate_63_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2750 = _T_2749[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2751 = $signed(_T_2750); // @[DenseLayer.scala 133:59]
  assign _GEN_462 = vld ? $signed(_T_2751) : $signed(cummulativeSums_63); // @[DenseLayer.scala 132:18]
  assign _GEN_463 = rst ? $signed(16'sh0) : $signed(_GEN_462); // @[DenseLayer.scala 135:18]
  assign _GEN_464 = _T_2438 ? $signed(MultiplyAccumulate_63_io_sum) : $signed(_GEN_463); // @[DenseLayer.scala 138:24]
  assign _T_2754 = $signed(cummulativeSums_64) + $signed(MultiplyAccumulate_64_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2755 = _T_2754[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2756 = $signed(_T_2755); // @[DenseLayer.scala 133:59]
  assign _GEN_465 = vld ? $signed(_T_2756) : $signed(cummulativeSums_64); // @[DenseLayer.scala 132:18]
  assign _GEN_466 = rst ? $signed(16'sh0) : $signed(_GEN_465); // @[DenseLayer.scala 135:18]
  assign _GEN_467 = _T_2438 ? $signed(MultiplyAccumulate_64_io_sum) : $signed(_GEN_466); // @[DenseLayer.scala 138:24]
  assign _T_2759 = $signed(cummulativeSums_65) + $signed(MultiplyAccumulate_65_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2760 = _T_2759[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2761 = $signed(_T_2760); // @[DenseLayer.scala 133:59]
  assign _GEN_468 = vld ? $signed(_T_2761) : $signed(cummulativeSums_65); // @[DenseLayer.scala 132:18]
  assign _GEN_469 = rst ? $signed(16'sh0) : $signed(_GEN_468); // @[DenseLayer.scala 135:18]
  assign _GEN_470 = _T_2438 ? $signed(MultiplyAccumulate_65_io_sum) : $signed(_GEN_469); // @[DenseLayer.scala 138:24]
  assign _T_2764 = $signed(cummulativeSums_66) + $signed(MultiplyAccumulate_66_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2765 = _T_2764[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2766 = $signed(_T_2765); // @[DenseLayer.scala 133:59]
  assign _GEN_471 = vld ? $signed(_T_2766) : $signed(cummulativeSums_66); // @[DenseLayer.scala 132:18]
  assign _GEN_472 = rst ? $signed(16'sh0) : $signed(_GEN_471); // @[DenseLayer.scala 135:18]
  assign _GEN_473 = _T_2438 ? $signed(MultiplyAccumulate_66_io_sum) : $signed(_GEN_472); // @[DenseLayer.scala 138:24]
  assign _T_2769 = $signed(cummulativeSums_67) + $signed(MultiplyAccumulate_67_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2770 = _T_2769[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2771 = $signed(_T_2770); // @[DenseLayer.scala 133:59]
  assign _GEN_474 = vld ? $signed(_T_2771) : $signed(cummulativeSums_67); // @[DenseLayer.scala 132:18]
  assign _GEN_475 = rst ? $signed(16'sh0) : $signed(_GEN_474); // @[DenseLayer.scala 135:18]
  assign _GEN_476 = _T_2438 ? $signed(MultiplyAccumulate_67_io_sum) : $signed(_GEN_475); // @[DenseLayer.scala 138:24]
  assign _T_2774 = $signed(cummulativeSums_68) + $signed(MultiplyAccumulate_68_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2775 = _T_2774[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2776 = $signed(_T_2775); // @[DenseLayer.scala 133:59]
  assign _GEN_477 = vld ? $signed(_T_2776) : $signed(cummulativeSums_68); // @[DenseLayer.scala 132:18]
  assign _GEN_478 = rst ? $signed(16'sh0) : $signed(_GEN_477); // @[DenseLayer.scala 135:18]
  assign _GEN_479 = _T_2438 ? $signed(MultiplyAccumulate_68_io_sum) : $signed(_GEN_478); // @[DenseLayer.scala 138:24]
  assign _T_2779 = $signed(cummulativeSums_69) + $signed(MultiplyAccumulate_69_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2780 = _T_2779[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2781 = $signed(_T_2780); // @[DenseLayer.scala 133:59]
  assign _GEN_480 = vld ? $signed(_T_2781) : $signed(cummulativeSums_69); // @[DenseLayer.scala 132:18]
  assign _GEN_481 = rst ? $signed(16'sh0) : $signed(_GEN_480); // @[DenseLayer.scala 135:18]
  assign _GEN_482 = _T_2438 ? $signed(MultiplyAccumulate_69_io_sum) : $signed(_GEN_481); // @[DenseLayer.scala 138:24]
  assign _T_2784 = $signed(cummulativeSums_70) + $signed(MultiplyAccumulate_70_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2785 = _T_2784[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2786 = $signed(_T_2785); // @[DenseLayer.scala 133:59]
  assign _GEN_483 = vld ? $signed(_T_2786) : $signed(cummulativeSums_70); // @[DenseLayer.scala 132:18]
  assign _GEN_484 = rst ? $signed(16'sh0) : $signed(_GEN_483); // @[DenseLayer.scala 135:18]
  assign _GEN_485 = _T_2438 ? $signed(MultiplyAccumulate_70_io_sum) : $signed(_GEN_484); // @[DenseLayer.scala 138:24]
  assign _T_2789 = $signed(cummulativeSums_71) + $signed(MultiplyAccumulate_71_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2790 = _T_2789[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2791 = $signed(_T_2790); // @[DenseLayer.scala 133:59]
  assign _GEN_486 = vld ? $signed(_T_2791) : $signed(cummulativeSums_71); // @[DenseLayer.scala 132:18]
  assign _GEN_487 = rst ? $signed(16'sh0) : $signed(_GEN_486); // @[DenseLayer.scala 135:18]
  assign _GEN_488 = _T_2438 ? $signed(MultiplyAccumulate_71_io_sum) : $signed(_GEN_487); // @[DenseLayer.scala 138:24]
  assign _T_2794 = $signed(cummulativeSums_72) + $signed(MultiplyAccumulate_72_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2795 = _T_2794[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2796 = $signed(_T_2795); // @[DenseLayer.scala 133:59]
  assign _GEN_489 = vld ? $signed(_T_2796) : $signed(cummulativeSums_72); // @[DenseLayer.scala 132:18]
  assign _GEN_490 = rst ? $signed(16'sh0) : $signed(_GEN_489); // @[DenseLayer.scala 135:18]
  assign _GEN_491 = _T_2438 ? $signed(MultiplyAccumulate_72_io_sum) : $signed(_GEN_490); // @[DenseLayer.scala 138:24]
  assign _T_2799 = $signed(cummulativeSums_73) + $signed(MultiplyAccumulate_73_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2800 = _T_2799[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2801 = $signed(_T_2800); // @[DenseLayer.scala 133:59]
  assign _GEN_492 = vld ? $signed(_T_2801) : $signed(cummulativeSums_73); // @[DenseLayer.scala 132:18]
  assign _GEN_493 = rst ? $signed(16'sh0) : $signed(_GEN_492); // @[DenseLayer.scala 135:18]
  assign _GEN_494 = _T_2438 ? $signed(MultiplyAccumulate_73_io_sum) : $signed(_GEN_493); // @[DenseLayer.scala 138:24]
  assign _T_2804 = $signed(cummulativeSums_74) + $signed(MultiplyAccumulate_74_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2805 = _T_2804[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2806 = $signed(_T_2805); // @[DenseLayer.scala 133:59]
  assign _GEN_495 = vld ? $signed(_T_2806) : $signed(cummulativeSums_74); // @[DenseLayer.scala 132:18]
  assign _GEN_496 = rst ? $signed(16'sh0) : $signed(_GEN_495); // @[DenseLayer.scala 135:18]
  assign _GEN_497 = _T_2438 ? $signed(MultiplyAccumulate_74_io_sum) : $signed(_GEN_496); // @[DenseLayer.scala 138:24]
  assign _T_2809 = $signed(cummulativeSums_75) + $signed(MultiplyAccumulate_75_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2810 = _T_2809[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2811 = $signed(_T_2810); // @[DenseLayer.scala 133:59]
  assign _GEN_498 = vld ? $signed(_T_2811) : $signed(cummulativeSums_75); // @[DenseLayer.scala 132:18]
  assign _GEN_499 = rst ? $signed(16'sh0) : $signed(_GEN_498); // @[DenseLayer.scala 135:18]
  assign _GEN_500 = _T_2438 ? $signed(MultiplyAccumulate_75_io_sum) : $signed(_GEN_499); // @[DenseLayer.scala 138:24]
  assign _T_2814 = $signed(cummulativeSums_76) + $signed(MultiplyAccumulate_76_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2815 = _T_2814[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2816 = $signed(_T_2815); // @[DenseLayer.scala 133:59]
  assign _GEN_501 = vld ? $signed(_T_2816) : $signed(cummulativeSums_76); // @[DenseLayer.scala 132:18]
  assign _GEN_502 = rst ? $signed(16'sh0) : $signed(_GEN_501); // @[DenseLayer.scala 135:18]
  assign _GEN_503 = _T_2438 ? $signed(MultiplyAccumulate_76_io_sum) : $signed(_GEN_502); // @[DenseLayer.scala 138:24]
  assign _T_2819 = $signed(cummulativeSums_77) + $signed(MultiplyAccumulate_77_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2820 = _T_2819[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2821 = $signed(_T_2820); // @[DenseLayer.scala 133:59]
  assign _GEN_504 = vld ? $signed(_T_2821) : $signed(cummulativeSums_77); // @[DenseLayer.scala 132:18]
  assign _GEN_505 = rst ? $signed(16'sh0) : $signed(_GEN_504); // @[DenseLayer.scala 135:18]
  assign _GEN_506 = _T_2438 ? $signed(MultiplyAccumulate_77_io_sum) : $signed(_GEN_505); // @[DenseLayer.scala 138:24]
  assign _T_2824 = $signed(cummulativeSums_78) + $signed(MultiplyAccumulate_78_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2825 = _T_2824[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2826 = $signed(_T_2825); // @[DenseLayer.scala 133:59]
  assign _GEN_507 = vld ? $signed(_T_2826) : $signed(cummulativeSums_78); // @[DenseLayer.scala 132:18]
  assign _GEN_508 = rst ? $signed(16'sh0) : $signed(_GEN_507); // @[DenseLayer.scala 135:18]
  assign _GEN_509 = _T_2438 ? $signed(MultiplyAccumulate_78_io_sum) : $signed(_GEN_508); // @[DenseLayer.scala 138:24]
  assign _T_2829 = $signed(cummulativeSums_79) + $signed(MultiplyAccumulate_79_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2830 = _T_2829[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2831 = $signed(_T_2830); // @[DenseLayer.scala 133:59]
  assign _GEN_510 = vld ? $signed(_T_2831) : $signed(cummulativeSums_79); // @[DenseLayer.scala 132:18]
  assign _GEN_511 = rst ? $signed(16'sh0) : $signed(_GEN_510); // @[DenseLayer.scala 135:18]
  assign _GEN_512 = _T_2438 ? $signed(MultiplyAccumulate_79_io_sum) : $signed(_GEN_511); // @[DenseLayer.scala 138:24]
  assign _T_2834 = $signed(cummulativeSums_80) + $signed(MultiplyAccumulate_80_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2835 = _T_2834[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2836 = $signed(_T_2835); // @[DenseLayer.scala 133:59]
  assign _GEN_513 = vld ? $signed(_T_2836) : $signed(cummulativeSums_80); // @[DenseLayer.scala 132:18]
  assign _GEN_514 = rst ? $signed(16'sh0) : $signed(_GEN_513); // @[DenseLayer.scala 135:18]
  assign _GEN_515 = _T_2438 ? $signed(MultiplyAccumulate_80_io_sum) : $signed(_GEN_514); // @[DenseLayer.scala 138:24]
  assign _T_2839 = $signed(cummulativeSums_81) + $signed(MultiplyAccumulate_81_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2840 = _T_2839[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2841 = $signed(_T_2840); // @[DenseLayer.scala 133:59]
  assign _GEN_516 = vld ? $signed(_T_2841) : $signed(cummulativeSums_81); // @[DenseLayer.scala 132:18]
  assign _GEN_517 = rst ? $signed(16'sh0) : $signed(_GEN_516); // @[DenseLayer.scala 135:18]
  assign _GEN_518 = _T_2438 ? $signed(MultiplyAccumulate_81_io_sum) : $signed(_GEN_517); // @[DenseLayer.scala 138:24]
  assign _T_2844 = $signed(cummulativeSums_82) + $signed(MultiplyAccumulate_82_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2845 = _T_2844[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2846 = $signed(_T_2845); // @[DenseLayer.scala 133:59]
  assign _GEN_519 = vld ? $signed(_T_2846) : $signed(cummulativeSums_82); // @[DenseLayer.scala 132:18]
  assign _GEN_520 = rst ? $signed(16'sh0) : $signed(_GEN_519); // @[DenseLayer.scala 135:18]
  assign _GEN_521 = _T_2438 ? $signed(MultiplyAccumulate_82_io_sum) : $signed(_GEN_520); // @[DenseLayer.scala 138:24]
  assign _T_2849 = $signed(cummulativeSums_83) + $signed(MultiplyAccumulate_83_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2850 = _T_2849[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2851 = $signed(_T_2850); // @[DenseLayer.scala 133:59]
  assign _GEN_522 = vld ? $signed(_T_2851) : $signed(cummulativeSums_83); // @[DenseLayer.scala 132:18]
  assign _GEN_523 = rst ? $signed(16'sh0) : $signed(_GEN_522); // @[DenseLayer.scala 135:18]
  assign _GEN_524 = _T_2438 ? $signed(MultiplyAccumulate_83_io_sum) : $signed(_GEN_523); // @[DenseLayer.scala 138:24]
  assign _T_2854 = $signed(cummulativeSums_84) + $signed(MultiplyAccumulate_84_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2855 = _T_2854[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2856 = $signed(_T_2855); // @[DenseLayer.scala 133:59]
  assign _GEN_525 = vld ? $signed(_T_2856) : $signed(cummulativeSums_84); // @[DenseLayer.scala 132:18]
  assign _GEN_526 = rst ? $signed(16'sh0) : $signed(_GEN_525); // @[DenseLayer.scala 135:18]
  assign _GEN_527 = _T_2438 ? $signed(MultiplyAccumulate_84_io_sum) : $signed(_GEN_526); // @[DenseLayer.scala 138:24]
  assign _T_2859 = $signed(cummulativeSums_85) + $signed(MultiplyAccumulate_85_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2860 = _T_2859[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2861 = $signed(_T_2860); // @[DenseLayer.scala 133:59]
  assign _GEN_528 = vld ? $signed(_T_2861) : $signed(cummulativeSums_85); // @[DenseLayer.scala 132:18]
  assign _GEN_529 = rst ? $signed(16'sh0) : $signed(_GEN_528); // @[DenseLayer.scala 135:18]
  assign _GEN_530 = _T_2438 ? $signed(MultiplyAccumulate_85_io_sum) : $signed(_GEN_529); // @[DenseLayer.scala 138:24]
  assign _T_2864 = $signed(cummulativeSums_86) + $signed(MultiplyAccumulate_86_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2865 = _T_2864[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2866 = $signed(_T_2865); // @[DenseLayer.scala 133:59]
  assign _GEN_531 = vld ? $signed(_T_2866) : $signed(cummulativeSums_86); // @[DenseLayer.scala 132:18]
  assign _GEN_532 = rst ? $signed(16'sh0) : $signed(_GEN_531); // @[DenseLayer.scala 135:18]
  assign _GEN_533 = _T_2438 ? $signed(MultiplyAccumulate_86_io_sum) : $signed(_GEN_532); // @[DenseLayer.scala 138:24]
  assign _T_2869 = $signed(cummulativeSums_87) + $signed(MultiplyAccumulate_87_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2870 = _T_2869[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2871 = $signed(_T_2870); // @[DenseLayer.scala 133:59]
  assign _GEN_534 = vld ? $signed(_T_2871) : $signed(cummulativeSums_87); // @[DenseLayer.scala 132:18]
  assign _GEN_535 = rst ? $signed(16'sh0) : $signed(_GEN_534); // @[DenseLayer.scala 135:18]
  assign _GEN_536 = _T_2438 ? $signed(MultiplyAccumulate_87_io_sum) : $signed(_GEN_535); // @[DenseLayer.scala 138:24]
  assign _T_2874 = $signed(cummulativeSums_88) + $signed(MultiplyAccumulate_88_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2875 = _T_2874[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2876 = $signed(_T_2875); // @[DenseLayer.scala 133:59]
  assign _GEN_537 = vld ? $signed(_T_2876) : $signed(cummulativeSums_88); // @[DenseLayer.scala 132:18]
  assign _GEN_538 = rst ? $signed(16'sh0) : $signed(_GEN_537); // @[DenseLayer.scala 135:18]
  assign _GEN_539 = _T_2438 ? $signed(MultiplyAccumulate_88_io_sum) : $signed(_GEN_538); // @[DenseLayer.scala 138:24]
  assign _T_2879 = $signed(cummulativeSums_89) + $signed(MultiplyAccumulate_89_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2880 = _T_2879[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2881 = $signed(_T_2880); // @[DenseLayer.scala 133:59]
  assign _GEN_540 = vld ? $signed(_T_2881) : $signed(cummulativeSums_89); // @[DenseLayer.scala 132:18]
  assign _GEN_541 = rst ? $signed(16'sh0) : $signed(_GEN_540); // @[DenseLayer.scala 135:18]
  assign _GEN_542 = _T_2438 ? $signed(MultiplyAccumulate_89_io_sum) : $signed(_GEN_541); // @[DenseLayer.scala 138:24]
  assign _T_2884 = $signed(cummulativeSums_90) + $signed(MultiplyAccumulate_90_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2885 = _T_2884[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2886 = $signed(_T_2885); // @[DenseLayer.scala 133:59]
  assign _GEN_543 = vld ? $signed(_T_2886) : $signed(cummulativeSums_90); // @[DenseLayer.scala 132:18]
  assign _GEN_544 = rst ? $signed(16'sh0) : $signed(_GEN_543); // @[DenseLayer.scala 135:18]
  assign _GEN_545 = _T_2438 ? $signed(MultiplyAccumulate_90_io_sum) : $signed(_GEN_544); // @[DenseLayer.scala 138:24]
  assign _T_2889 = $signed(cummulativeSums_91) + $signed(MultiplyAccumulate_91_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2890 = _T_2889[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2891 = $signed(_T_2890); // @[DenseLayer.scala 133:59]
  assign _GEN_546 = vld ? $signed(_T_2891) : $signed(cummulativeSums_91); // @[DenseLayer.scala 132:18]
  assign _GEN_547 = rst ? $signed(16'sh0) : $signed(_GEN_546); // @[DenseLayer.scala 135:18]
  assign _GEN_548 = _T_2438 ? $signed(MultiplyAccumulate_91_io_sum) : $signed(_GEN_547); // @[DenseLayer.scala 138:24]
  assign _T_2894 = $signed(cummulativeSums_92) + $signed(MultiplyAccumulate_92_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2895 = _T_2894[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2896 = $signed(_T_2895); // @[DenseLayer.scala 133:59]
  assign _GEN_549 = vld ? $signed(_T_2896) : $signed(cummulativeSums_92); // @[DenseLayer.scala 132:18]
  assign _GEN_550 = rst ? $signed(16'sh0) : $signed(_GEN_549); // @[DenseLayer.scala 135:18]
  assign _GEN_551 = _T_2438 ? $signed(MultiplyAccumulate_92_io_sum) : $signed(_GEN_550); // @[DenseLayer.scala 138:24]
  assign _T_2899 = $signed(cummulativeSums_93) + $signed(MultiplyAccumulate_93_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2900 = _T_2899[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2901 = $signed(_T_2900); // @[DenseLayer.scala 133:59]
  assign _GEN_552 = vld ? $signed(_T_2901) : $signed(cummulativeSums_93); // @[DenseLayer.scala 132:18]
  assign _GEN_553 = rst ? $signed(16'sh0) : $signed(_GEN_552); // @[DenseLayer.scala 135:18]
  assign _GEN_554 = _T_2438 ? $signed(MultiplyAccumulate_93_io_sum) : $signed(_GEN_553); // @[DenseLayer.scala 138:24]
  assign _T_2904 = $signed(cummulativeSums_94) + $signed(MultiplyAccumulate_94_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2905 = _T_2904[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2906 = $signed(_T_2905); // @[DenseLayer.scala 133:59]
  assign _GEN_555 = vld ? $signed(_T_2906) : $signed(cummulativeSums_94); // @[DenseLayer.scala 132:18]
  assign _GEN_556 = rst ? $signed(16'sh0) : $signed(_GEN_555); // @[DenseLayer.scala 135:18]
  assign _GEN_557 = _T_2438 ? $signed(MultiplyAccumulate_94_io_sum) : $signed(_GEN_556); // @[DenseLayer.scala 138:24]
  assign _T_2909 = $signed(cummulativeSums_95) + $signed(MultiplyAccumulate_95_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2910 = _T_2909[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2911 = $signed(_T_2910); // @[DenseLayer.scala 133:59]
  assign _GEN_558 = vld ? $signed(_T_2911) : $signed(cummulativeSums_95); // @[DenseLayer.scala 132:18]
  assign _GEN_559 = rst ? $signed(16'sh0) : $signed(_GEN_558); // @[DenseLayer.scala 135:18]
  assign _GEN_560 = _T_2438 ? $signed(MultiplyAccumulate_95_io_sum) : $signed(_GEN_559); // @[DenseLayer.scala 138:24]
  assign _T_2914 = $signed(cummulativeSums_96) + $signed(MultiplyAccumulate_96_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2915 = _T_2914[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2916 = $signed(_T_2915); // @[DenseLayer.scala 133:59]
  assign _GEN_561 = vld ? $signed(_T_2916) : $signed(cummulativeSums_96); // @[DenseLayer.scala 132:18]
  assign _GEN_562 = rst ? $signed(16'sh0) : $signed(_GEN_561); // @[DenseLayer.scala 135:18]
  assign _GEN_563 = _T_2438 ? $signed(MultiplyAccumulate_96_io_sum) : $signed(_GEN_562); // @[DenseLayer.scala 138:24]
  assign _T_2919 = $signed(cummulativeSums_97) + $signed(MultiplyAccumulate_97_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2920 = _T_2919[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2921 = $signed(_T_2920); // @[DenseLayer.scala 133:59]
  assign _GEN_564 = vld ? $signed(_T_2921) : $signed(cummulativeSums_97); // @[DenseLayer.scala 132:18]
  assign _GEN_565 = rst ? $signed(16'sh0) : $signed(_GEN_564); // @[DenseLayer.scala 135:18]
  assign _GEN_566 = _T_2438 ? $signed(MultiplyAccumulate_97_io_sum) : $signed(_GEN_565); // @[DenseLayer.scala 138:24]
  assign _T_2924 = $signed(cummulativeSums_98) + $signed(MultiplyAccumulate_98_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2925 = _T_2924[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2926 = $signed(_T_2925); // @[DenseLayer.scala 133:59]
  assign _GEN_567 = vld ? $signed(_T_2926) : $signed(cummulativeSums_98); // @[DenseLayer.scala 132:18]
  assign _GEN_568 = rst ? $signed(16'sh0) : $signed(_GEN_567); // @[DenseLayer.scala 135:18]
  assign _GEN_569 = _T_2438 ? $signed(MultiplyAccumulate_98_io_sum) : $signed(_GEN_568); // @[DenseLayer.scala 138:24]
  assign _T_2929 = $signed(cummulativeSums_99) + $signed(MultiplyAccumulate_99_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2930 = _T_2929[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2931 = $signed(_T_2930); // @[DenseLayer.scala 133:59]
  assign _GEN_570 = vld ? $signed(_T_2931) : $signed(cummulativeSums_99); // @[DenseLayer.scala 132:18]
  assign _GEN_571 = rst ? $signed(16'sh0) : $signed(_GEN_570); // @[DenseLayer.scala 135:18]
  assign _GEN_572 = _T_2438 ? $signed(MultiplyAccumulate_99_io_sum) : $signed(_GEN_571); // @[DenseLayer.scala 138:24]
  assign _T_2934 = $signed(cummulativeSums_100) + $signed(MultiplyAccumulate_100_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2935 = _T_2934[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2936 = $signed(_T_2935); // @[DenseLayer.scala 133:59]
  assign _GEN_573 = vld ? $signed(_T_2936) : $signed(cummulativeSums_100); // @[DenseLayer.scala 132:18]
  assign _GEN_574 = rst ? $signed(16'sh0) : $signed(_GEN_573); // @[DenseLayer.scala 135:18]
  assign _GEN_575 = _T_2438 ? $signed(MultiplyAccumulate_100_io_sum) : $signed(_GEN_574); // @[DenseLayer.scala 138:24]
  assign _T_2939 = $signed(cummulativeSums_101) + $signed(MultiplyAccumulate_101_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2940 = _T_2939[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2941 = $signed(_T_2940); // @[DenseLayer.scala 133:59]
  assign _GEN_576 = vld ? $signed(_T_2941) : $signed(cummulativeSums_101); // @[DenseLayer.scala 132:18]
  assign _GEN_577 = rst ? $signed(16'sh0) : $signed(_GEN_576); // @[DenseLayer.scala 135:18]
  assign _GEN_578 = _T_2438 ? $signed(MultiplyAccumulate_101_io_sum) : $signed(_GEN_577); // @[DenseLayer.scala 138:24]
  assign _T_2944 = $signed(cummulativeSums_102) + $signed(MultiplyAccumulate_102_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2945 = _T_2944[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2946 = $signed(_T_2945); // @[DenseLayer.scala 133:59]
  assign _GEN_579 = vld ? $signed(_T_2946) : $signed(cummulativeSums_102); // @[DenseLayer.scala 132:18]
  assign _GEN_580 = rst ? $signed(16'sh0) : $signed(_GEN_579); // @[DenseLayer.scala 135:18]
  assign _GEN_581 = _T_2438 ? $signed(MultiplyAccumulate_102_io_sum) : $signed(_GEN_580); // @[DenseLayer.scala 138:24]
  assign _T_2949 = $signed(cummulativeSums_103) + $signed(MultiplyAccumulate_103_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2950 = _T_2949[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2951 = $signed(_T_2950); // @[DenseLayer.scala 133:59]
  assign _GEN_582 = vld ? $signed(_T_2951) : $signed(cummulativeSums_103); // @[DenseLayer.scala 132:18]
  assign _GEN_583 = rst ? $signed(16'sh0) : $signed(_GEN_582); // @[DenseLayer.scala 135:18]
  assign _GEN_584 = _T_2438 ? $signed(MultiplyAccumulate_103_io_sum) : $signed(_GEN_583); // @[DenseLayer.scala 138:24]
  assign _T_2954 = $signed(cummulativeSums_104) + $signed(MultiplyAccumulate_104_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2955 = _T_2954[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2956 = $signed(_T_2955); // @[DenseLayer.scala 133:59]
  assign _GEN_585 = vld ? $signed(_T_2956) : $signed(cummulativeSums_104); // @[DenseLayer.scala 132:18]
  assign _GEN_586 = rst ? $signed(16'sh0) : $signed(_GEN_585); // @[DenseLayer.scala 135:18]
  assign _GEN_587 = _T_2438 ? $signed(MultiplyAccumulate_104_io_sum) : $signed(_GEN_586); // @[DenseLayer.scala 138:24]
  assign _T_2959 = $signed(cummulativeSums_105) + $signed(MultiplyAccumulate_105_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2960 = _T_2959[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2961 = $signed(_T_2960); // @[DenseLayer.scala 133:59]
  assign _GEN_588 = vld ? $signed(_T_2961) : $signed(cummulativeSums_105); // @[DenseLayer.scala 132:18]
  assign _GEN_589 = rst ? $signed(16'sh0) : $signed(_GEN_588); // @[DenseLayer.scala 135:18]
  assign _GEN_590 = _T_2438 ? $signed(MultiplyAccumulate_105_io_sum) : $signed(_GEN_589); // @[DenseLayer.scala 138:24]
  assign _T_2964 = $signed(cummulativeSums_106) + $signed(MultiplyAccumulate_106_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2965 = _T_2964[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2966 = $signed(_T_2965); // @[DenseLayer.scala 133:59]
  assign _GEN_591 = vld ? $signed(_T_2966) : $signed(cummulativeSums_106); // @[DenseLayer.scala 132:18]
  assign _GEN_592 = rst ? $signed(16'sh0) : $signed(_GEN_591); // @[DenseLayer.scala 135:18]
  assign _GEN_593 = _T_2438 ? $signed(MultiplyAccumulate_106_io_sum) : $signed(_GEN_592); // @[DenseLayer.scala 138:24]
  assign _T_2969 = $signed(cummulativeSums_107) + $signed(MultiplyAccumulate_107_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2970 = _T_2969[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2971 = $signed(_T_2970); // @[DenseLayer.scala 133:59]
  assign _GEN_594 = vld ? $signed(_T_2971) : $signed(cummulativeSums_107); // @[DenseLayer.scala 132:18]
  assign _GEN_595 = rst ? $signed(16'sh0) : $signed(_GEN_594); // @[DenseLayer.scala 135:18]
  assign _GEN_596 = _T_2438 ? $signed(MultiplyAccumulate_107_io_sum) : $signed(_GEN_595); // @[DenseLayer.scala 138:24]
  assign _T_2974 = $signed(cummulativeSums_108) + $signed(MultiplyAccumulate_108_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2975 = _T_2974[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2976 = $signed(_T_2975); // @[DenseLayer.scala 133:59]
  assign _GEN_597 = vld ? $signed(_T_2976) : $signed(cummulativeSums_108); // @[DenseLayer.scala 132:18]
  assign _GEN_598 = rst ? $signed(16'sh0) : $signed(_GEN_597); // @[DenseLayer.scala 135:18]
  assign _GEN_599 = _T_2438 ? $signed(MultiplyAccumulate_108_io_sum) : $signed(_GEN_598); // @[DenseLayer.scala 138:24]
  assign _T_2979 = $signed(cummulativeSums_109) + $signed(MultiplyAccumulate_109_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2980 = _T_2979[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2981 = $signed(_T_2980); // @[DenseLayer.scala 133:59]
  assign _GEN_600 = vld ? $signed(_T_2981) : $signed(cummulativeSums_109); // @[DenseLayer.scala 132:18]
  assign _GEN_601 = rst ? $signed(16'sh0) : $signed(_GEN_600); // @[DenseLayer.scala 135:18]
  assign _GEN_602 = _T_2438 ? $signed(MultiplyAccumulate_109_io_sum) : $signed(_GEN_601); // @[DenseLayer.scala 138:24]
  assign _T_2984 = $signed(cummulativeSums_110) + $signed(MultiplyAccumulate_110_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2985 = _T_2984[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2986 = $signed(_T_2985); // @[DenseLayer.scala 133:59]
  assign _GEN_603 = vld ? $signed(_T_2986) : $signed(cummulativeSums_110); // @[DenseLayer.scala 132:18]
  assign _GEN_604 = rst ? $signed(16'sh0) : $signed(_GEN_603); // @[DenseLayer.scala 135:18]
  assign _GEN_605 = _T_2438 ? $signed(MultiplyAccumulate_110_io_sum) : $signed(_GEN_604); // @[DenseLayer.scala 138:24]
  assign _T_2989 = $signed(cummulativeSums_111) + $signed(MultiplyAccumulate_111_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2990 = _T_2989[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2991 = $signed(_T_2990); // @[DenseLayer.scala 133:59]
  assign _GEN_606 = vld ? $signed(_T_2991) : $signed(cummulativeSums_111); // @[DenseLayer.scala 132:18]
  assign _GEN_607 = rst ? $signed(16'sh0) : $signed(_GEN_606); // @[DenseLayer.scala 135:18]
  assign _GEN_608 = _T_2438 ? $signed(MultiplyAccumulate_111_io_sum) : $signed(_GEN_607); // @[DenseLayer.scala 138:24]
  assign _T_2994 = $signed(cummulativeSums_112) + $signed(MultiplyAccumulate_112_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_2995 = _T_2994[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_2996 = $signed(_T_2995); // @[DenseLayer.scala 133:59]
  assign _GEN_609 = vld ? $signed(_T_2996) : $signed(cummulativeSums_112); // @[DenseLayer.scala 132:18]
  assign _GEN_610 = rst ? $signed(16'sh0) : $signed(_GEN_609); // @[DenseLayer.scala 135:18]
  assign _GEN_611 = _T_2438 ? $signed(MultiplyAccumulate_112_io_sum) : $signed(_GEN_610); // @[DenseLayer.scala 138:24]
  assign _T_2999 = $signed(cummulativeSums_113) + $signed(MultiplyAccumulate_113_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_3000 = _T_2999[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_3001 = $signed(_T_3000); // @[DenseLayer.scala 133:59]
  assign _GEN_612 = vld ? $signed(_T_3001) : $signed(cummulativeSums_113); // @[DenseLayer.scala 132:18]
  assign _GEN_613 = rst ? $signed(16'sh0) : $signed(_GEN_612); // @[DenseLayer.scala 135:18]
  assign _GEN_614 = _T_2438 ? $signed(MultiplyAccumulate_113_io_sum) : $signed(_GEN_613); // @[DenseLayer.scala 138:24]
  assign _T_3004 = $signed(cummulativeSums_114) + $signed(MultiplyAccumulate_114_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_3005 = _T_3004[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_3006 = $signed(_T_3005); // @[DenseLayer.scala 133:59]
  assign _GEN_615 = vld ? $signed(_T_3006) : $signed(cummulativeSums_114); // @[DenseLayer.scala 132:18]
  assign _GEN_616 = rst ? $signed(16'sh0) : $signed(_GEN_615); // @[DenseLayer.scala 135:18]
  assign _GEN_617 = _T_2438 ? $signed(MultiplyAccumulate_114_io_sum) : $signed(_GEN_616); // @[DenseLayer.scala 138:24]
  assign _T_3009 = $signed(cummulativeSums_115) + $signed(MultiplyAccumulate_115_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_3010 = _T_3009[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_3011 = $signed(_T_3010); // @[DenseLayer.scala 133:59]
  assign _GEN_618 = vld ? $signed(_T_3011) : $signed(cummulativeSums_115); // @[DenseLayer.scala 132:18]
  assign _GEN_619 = rst ? $signed(16'sh0) : $signed(_GEN_618); // @[DenseLayer.scala 135:18]
  assign _GEN_620 = _T_2438 ? $signed(MultiplyAccumulate_115_io_sum) : $signed(_GEN_619); // @[DenseLayer.scala 138:24]
  assign _T_3014 = $signed(cummulativeSums_116) + $signed(MultiplyAccumulate_116_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_3015 = _T_3014[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_3016 = $signed(_T_3015); // @[DenseLayer.scala 133:59]
  assign _GEN_621 = vld ? $signed(_T_3016) : $signed(cummulativeSums_116); // @[DenseLayer.scala 132:18]
  assign _GEN_622 = rst ? $signed(16'sh0) : $signed(_GEN_621); // @[DenseLayer.scala 135:18]
  assign _GEN_623 = _T_2438 ? $signed(MultiplyAccumulate_116_io_sum) : $signed(_GEN_622); // @[DenseLayer.scala 138:24]
  assign _T_3019 = $signed(cummulativeSums_117) + $signed(MultiplyAccumulate_117_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_3020 = _T_3019[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_3021 = $signed(_T_3020); // @[DenseLayer.scala 133:59]
  assign _GEN_624 = vld ? $signed(_T_3021) : $signed(cummulativeSums_117); // @[DenseLayer.scala 132:18]
  assign _GEN_625 = rst ? $signed(16'sh0) : $signed(_GEN_624); // @[DenseLayer.scala 135:18]
  assign _GEN_626 = _T_2438 ? $signed(MultiplyAccumulate_117_io_sum) : $signed(_GEN_625); // @[DenseLayer.scala 138:24]
  assign _T_3024 = $signed(cummulativeSums_118) + $signed(MultiplyAccumulate_118_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_3025 = _T_3024[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_3026 = $signed(_T_3025); // @[DenseLayer.scala 133:59]
  assign _GEN_627 = vld ? $signed(_T_3026) : $signed(cummulativeSums_118); // @[DenseLayer.scala 132:18]
  assign _GEN_628 = rst ? $signed(16'sh0) : $signed(_GEN_627); // @[DenseLayer.scala 135:18]
  assign _GEN_629 = _T_2438 ? $signed(MultiplyAccumulate_118_io_sum) : $signed(_GEN_628); // @[DenseLayer.scala 138:24]
  assign _T_3029 = $signed(cummulativeSums_119) + $signed(MultiplyAccumulate_119_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_3030 = _T_3029[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_3031 = $signed(_T_3030); // @[DenseLayer.scala 133:59]
  assign _GEN_630 = vld ? $signed(_T_3031) : $signed(cummulativeSums_119); // @[DenseLayer.scala 132:18]
  assign _GEN_631 = rst ? $signed(16'sh0) : $signed(_GEN_630); // @[DenseLayer.scala 135:18]
  assign _GEN_632 = _T_2438 ? $signed(MultiplyAccumulate_119_io_sum) : $signed(_GEN_631); // @[DenseLayer.scala 138:24]
  assign _T_3034 = $signed(cummulativeSums_120) + $signed(MultiplyAccumulate_120_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_3035 = _T_3034[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_3036 = $signed(_T_3035); // @[DenseLayer.scala 133:59]
  assign _GEN_633 = vld ? $signed(_T_3036) : $signed(cummulativeSums_120); // @[DenseLayer.scala 132:18]
  assign _GEN_634 = rst ? $signed(16'sh0) : $signed(_GEN_633); // @[DenseLayer.scala 135:18]
  assign _GEN_635 = _T_2438 ? $signed(MultiplyAccumulate_120_io_sum) : $signed(_GEN_634); // @[DenseLayer.scala 138:24]
  assign _T_3039 = $signed(cummulativeSums_121) + $signed(MultiplyAccumulate_121_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_3040 = _T_3039[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_3041 = $signed(_T_3040); // @[DenseLayer.scala 133:59]
  assign _GEN_636 = vld ? $signed(_T_3041) : $signed(cummulativeSums_121); // @[DenseLayer.scala 132:18]
  assign _GEN_637 = rst ? $signed(16'sh0) : $signed(_GEN_636); // @[DenseLayer.scala 135:18]
  assign _GEN_638 = _T_2438 ? $signed(MultiplyAccumulate_121_io_sum) : $signed(_GEN_637); // @[DenseLayer.scala 138:24]
  assign _T_3044 = $signed(cummulativeSums_122) + $signed(MultiplyAccumulate_122_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_3045 = _T_3044[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_3046 = $signed(_T_3045); // @[DenseLayer.scala 133:59]
  assign _GEN_639 = vld ? $signed(_T_3046) : $signed(cummulativeSums_122); // @[DenseLayer.scala 132:18]
  assign _GEN_640 = rst ? $signed(16'sh0) : $signed(_GEN_639); // @[DenseLayer.scala 135:18]
  assign _GEN_641 = _T_2438 ? $signed(MultiplyAccumulate_122_io_sum) : $signed(_GEN_640); // @[DenseLayer.scala 138:24]
  assign _T_3049 = $signed(cummulativeSums_123) + $signed(MultiplyAccumulate_123_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_3050 = _T_3049[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_3051 = $signed(_T_3050); // @[DenseLayer.scala 133:59]
  assign _GEN_642 = vld ? $signed(_T_3051) : $signed(cummulativeSums_123); // @[DenseLayer.scala 132:18]
  assign _GEN_643 = rst ? $signed(16'sh0) : $signed(_GEN_642); // @[DenseLayer.scala 135:18]
  assign _GEN_644 = _T_2438 ? $signed(MultiplyAccumulate_123_io_sum) : $signed(_GEN_643); // @[DenseLayer.scala 138:24]
  assign _T_3054 = $signed(cummulativeSums_124) + $signed(MultiplyAccumulate_124_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_3055 = _T_3054[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_3056 = $signed(_T_3055); // @[DenseLayer.scala 133:59]
  assign _GEN_645 = vld ? $signed(_T_3056) : $signed(cummulativeSums_124); // @[DenseLayer.scala 132:18]
  assign _GEN_646 = rst ? $signed(16'sh0) : $signed(_GEN_645); // @[DenseLayer.scala 135:18]
  assign _GEN_647 = _T_2438 ? $signed(MultiplyAccumulate_124_io_sum) : $signed(_GEN_646); // @[DenseLayer.scala 138:24]
  assign _T_3059 = $signed(cummulativeSums_125) + $signed(MultiplyAccumulate_125_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_3060 = _T_3059[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_3061 = $signed(_T_3060); // @[DenseLayer.scala 133:59]
  assign _GEN_648 = vld ? $signed(_T_3061) : $signed(cummulativeSums_125); // @[DenseLayer.scala 132:18]
  assign _GEN_649 = rst ? $signed(16'sh0) : $signed(_GEN_648); // @[DenseLayer.scala 135:18]
  assign _GEN_650 = _T_2438 ? $signed(MultiplyAccumulate_125_io_sum) : $signed(_GEN_649); // @[DenseLayer.scala 138:24]
  assign _T_3064 = $signed(cummulativeSums_126) + $signed(MultiplyAccumulate_126_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_3065 = _T_3064[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_3066 = $signed(_T_3065); // @[DenseLayer.scala 133:59]
  assign _GEN_651 = vld ? $signed(_T_3066) : $signed(cummulativeSums_126); // @[DenseLayer.scala 132:18]
  assign _GEN_652 = rst ? $signed(16'sh0) : $signed(_GEN_651); // @[DenseLayer.scala 135:18]
  assign _GEN_653 = _T_2438 ? $signed(MultiplyAccumulate_126_io_sum) : $signed(_GEN_652); // @[DenseLayer.scala 138:24]
  assign _T_3069 = $signed(cummulativeSums_127) + $signed(MultiplyAccumulate_127_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_3070 = _T_3069[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_3071 = $signed(_T_3070); // @[DenseLayer.scala 133:59]
  assign _GEN_654 = vld ? $signed(_T_3071) : $signed(cummulativeSums_127); // @[DenseLayer.scala 132:18]
  assign _GEN_655 = rst ? $signed(16'sh0) : $signed(_GEN_654); // @[DenseLayer.scala 135:18]
  assign _GEN_656 = _T_2438 ? $signed(MultiplyAccumulate_127_io_sum) : $signed(_GEN_655); // @[DenseLayer.scala 138:24]
  assign io_dataOut_valid = _T_2418;
  assign io_dataOut_bits_0 = cummulativeSums_0;
  assign io_dataOut_bits_1 = cummulativeSums_1;
  assign io_dataOut_bits_2 = cummulativeSums_2;
  assign io_dataOut_bits_3 = cummulativeSums_3;
  assign io_dataOut_bits_4 = cummulativeSums_4;
  assign io_dataOut_bits_5 = cummulativeSums_5;
  assign io_dataOut_bits_6 = cummulativeSums_6;
  assign io_dataOut_bits_7 = cummulativeSums_7;
  assign io_dataOut_bits_8 = cummulativeSums_8;
  assign io_dataOut_bits_9 = cummulativeSums_9;
  assign io_dataOut_bits_10 = cummulativeSums_10;
  assign io_dataOut_bits_11 = cummulativeSums_11;
  assign io_dataOut_bits_12 = cummulativeSums_12;
  assign io_dataOut_bits_13 = cummulativeSums_13;
  assign io_dataOut_bits_14 = cummulativeSums_14;
  assign io_dataOut_bits_15 = cummulativeSums_15;
  assign io_dataOut_bits_16 = cummulativeSums_16;
  assign io_dataOut_bits_17 = cummulativeSums_17;
  assign io_dataOut_bits_18 = cummulativeSums_18;
  assign io_dataOut_bits_19 = cummulativeSums_19;
  assign io_dataOut_bits_20 = cummulativeSums_20;
  assign io_dataOut_bits_21 = cummulativeSums_21;
  assign io_dataOut_bits_22 = cummulativeSums_22;
  assign io_dataOut_bits_23 = cummulativeSums_23;
  assign io_dataOut_bits_24 = cummulativeSums_24;
  assign io_dataOut_bits_25 = cummulativeSums_25;
  assign io_dataOut_bits_26 = cummulativeSums_26;
  assign io_dataOut_bits_27 = cummulativeSums_27;
  assign io_dataOut_bits_28 = cummulativeSums_28;
  assign io_dataOut_bits_29 = cummulativeSums_29;
  assign io_dataOut_bits_30 = cummulativeSums_30;
  assign io_dataOut_bits_31 = cummulativeSums_31;
  assign io_dataOut_bits_32 = cummulativeSums_32;
  assign io_dataOut_bits_33 = cummulativeSums_33;
  assign io_dataOut_bits_34 = cummulativeSums_34;
  assign io_dataOut_bits_35 = cummulativeSums_35;
  assign io_dataOut_bits_36 = cummulativeSums_36;
  assign io_dataOut_bits_37 = cummulativeSums_37;
  assign io_dataOut_bits_38 = cummulativeSums_38;
  assign io_dataOut_bits_39 = cummulativeSums_39;
  assign io_dataOut_bits_40 = cummulativeSums_40;
  assign io_dataOut_bits_41 = cummulativeSums_41;
  assign io_dataOut_bits_42 = cummulativeSums_42;
  assign io_dataOut_bits_43 = cummulativeSums_43;
  assign io_dataOut_bits_44 = cummulativeSums_44;
  assign io_dataOut_bits_45 = cummulativeSums_45;
  assign io_dataOut_bits_46 = cummulativeSums_46;
  assign io_dataOut_bits_47 = cummulativeSums_47;
  assign io_dataOut_bits_48 = cummulativeSums_48;
  assign io_dataOut_bits_49 = cummulativeSums_49;
  assign io_dataOut_bits_50 = cummulativeSums_50;
  assign io_dataOut_bits_51 = cummulativeSums_51;
  assign io_dataOut_bits_52 = cummulativeSums_52;
  assign io_dataOut_bits_53 = cummulativeSums_53;
  assign io_dataOut_bits_54 = cummulativeSums_54;
  assign io_dataOut_bits_55 = cummulativeSums_55;
  assign io_dataOut_bits_56 = cummulativeSums_56;
  assign io_dataOut_bits_57 = cummulativeSums_57;
  assign io_dataOut_bits_58 = cummulativeSums_58;
  assign io_dataOut_bits_59 = cummulativeSums_59;
  assign io_dataOut_bits_60 = cummulativeSums_60;
  assign io_dataOut_bits_61 = cummulativeSums_61;
  assign io_dataOut_bits_62 = cummulativeSums_62;
  assign io_dataOut_bits_63 = cummulativeSums_63;
  assign io_dataOut_bits_64 = cummulativeSums_64;
  assign io_dataOut_bits_65 = cummulativeSums_65;
  assign io_dataOut_bits_66 = cummulativeSums_66;
  assign io_dataOut_bits_67 = cummulativeSums_67;
  assign io_dataOut_bits_68 = cummulativeSums_68;
  assign io_dataOut_bits_69 = cummulativeSums_69;
  assign io_dataOut_bits_70 = cummulativeSums_70;
  assign io_dataOut_bits_71 = cummulativeSums_71;
  assign io_dataOut_bits_72 = cummulativeSums_72;
  assign io_dataOut_bits_73 = cummulativeSums_73;
  assign io_dataOut_bits_74 = cummulativeSums_74;
  assign io_dataOut_bits_75 = cummulativeSums_75;
  assign io_dataOut_bits_76 = cummulativeSums_76;
  assign io_dataOut_bits_77 = cummulativeSums_77;
  assign io_dataOut_bits_78 = cummulativeSums_78;
  assign io_dataOut_bits_79 = cummulativeSums_79;
  assign io_dataOut_bits_80 = cummulativeSums_80;
  assign io_dataOut_bits_81 = cummulativeSums_81;
  assign io_dataOut_bits_82 = cummulativeSums_82;
  assign io_dataOut_bits_83 = cummulativeSums_83;
  assign io_dataOut_bits_84 = cummulativeSums_84;
  assign io_dataOut_bits_85 = cummulativeSums_85;
  assign io_dataOut_bits_86 = cummulativeSums_86;
  assign io_dataOut_bits_87 = cummulativeSums_87;
  assign io_dataOut_bits_88 = cummulativeSums_88;
  assign io_dataOut_bits_89 = cummulativeSums_89;
  assign io_dataOut_bits_90 = cummulativeSums_90;
  assign io_dataOut_bits_91 = cummulativeSums_91;
  assign io_dataOut_bits_92 = cummulativeSums_92;
  assign io_dataOut_bits_93 = cummulativeSums_93;
  assign io_dataOut_bits_94 = cummulativeSums_94;
  assign io_dataOut_bits_95 = cummulativeSums_95;
  assign io_dataOut_bits_96 = cummulativeSums_96;
  assign io_dataOut_bits_97 = cummulativeSums_97;
  assign io_dataOut_bits_98 = cummulativeSums_98;
  assign io_dataOut_bits_99 = cummulativeSums_99;
  assign io_dataOut_bits_100 = cummulativeSums_100;
  assign io_dataOut_bits_101 = cummulativeSums_101;
  assign io_dataOut_bits_102 = cummulativeSums_102;
  assign io_dataOut_bits_103 = cummulativeSums_103;
  assign io_dataOut_bits_104 = cummulativeSums_104;
  assign io_dataOut_bits_105 = cummulativeSums_105;
  assign io_dataOut_bits_106 = cummulativeSums_106;
  assign io_dataOut_bits_107 = cummulativeSums_107;
  assign io_dataOut_bits_108 = cummulativeSums_108;
  assign io_dataOut_bits_109 = cummulativeSums_109;
  assign io_dataOut_bits_110 = cummulativeSums_110;
  assign io_dataOut_bits_111 = cummulativeSums_111;
  assign io_dataOut_bits_112 = cummulativeSums_112;
  assign io_dataOut_bits_113 = cummulativeSums_113;
  assign io_dataOut_bits_114 = cummulativeSums_114;
  assign io_dataOut_bits_115 = cummulativeSums_115;
  assign io_dataOut_bits_116 = cummulativeSums_116;
  assign io_dataOut_bits_117 = cummulativeSums_117;
  assign io_dataOut_bits_118 = cummulativeSums_118;
  assign io_dataOut_bits_119 = cummulativeSums_119;
  assign io_dataOut_bits_120 = cummulativeSums_120;
  assign io_dataOut_bits_121 = cummulativeSums_121;
  assign io_dataOut_bits_122 = cummulativeSums_122;
  assign io_dataOut_bits_123 = cummulativeSums_123;
  assign io_dataOut_bits_124 = cummulativeSums_124;
  assign io_dataOut_bits_125 = cummulativeSums_125;
  assign io_dataOut_bits_126 = cummulativeSums_126;
  assign io_dataOut_bits_127 = cummulativeSums_127;
  assign weightsRAM_readAddr = _T_293;
  assign weightsRAM_clock = clock;
  assign FanoutAWS_clock = clock;
  assign FanoutAWS_io_in = currActs_0;
  assign FanoutAWS_1_clock = clock;
  assign FanoutAWS_1_io_in = currActs_1;
  assign FanoutAWS_2_clock = clock;
  assign FanoutAWS_2_io_in = currActs_2;
  assign FanoutAWS_3_clock = clock;
  assign FanoutAWS_3_io_in = currActs_3;
  assign MultiplyAccumulate_clock = clock;
  assign MultiplyAccumulate_io_activations_0 = FanoutAWS_io_out_0;
  assign MultiplyAccumulate_io_activations_1 = FanoutAWS_1_io_out_0;
  assign MultiplyAccumulate_io_activations_2 = FanoutAWS_2_io_out_0;
  assign MultiplyAccumulate_io_activations_3 = FanoutAWS_3_io_out_0;
  assign MultiplyAccumulate_io_weights = delayWeights_0;
  assign MultiplyAccumulate_1_clock = clock;
  assign MultiplyAccumulate_1_io_activations_0 = FanoutAWS_io_out_1;
  assign MultiplyAccumulate_1_io_activations_1 = FanoutAWS_1_io_out_1;
  assign MultiplyAccumulate_1_io_activations_2 = FanoutAWS_2_io_out_1;
  assign MultiplyAccumulate_1_io_activations_3 = FanoutAWS_3_io_out_1;
  assign MultiplyAccumulate_1_io_weights = delayWeights_1;
  assign MultiplyAccumulate_2_clock = clock;
  assign MultiplyAccumulate_2_io_activations_0 = FanoutAWS_io_out_2;
  assign MultiplyAccumulate_2_io_activations_1 = FanoutAWS_1_io_out_2;
  assign MultiplyAccumulate_2_io_activations_2 = FanoutAWS_2_io_out_2;
  assign MultiplyAccumulate_2_io_activations_3 = FanoutAWS_3_io_out_2;
  assign MultiplyAccumulate_2_io_weights = delayWeights_2;
  assign MultiplyAccumulate_3_clock = clock;
  assign MultiplyAccumulate_3_io_activations_0 = FanoutAWS_io_out_3;
  assign MultiplyAccumulate_3_io_activations_1 = FanoutAWS_1_io_out_3;
  assign MultiplyAccumulate_3_io_activations_2 = FanoutAWS_2_io_out_3;
  assign MultiplyAccumulate_3_io_activations_3 = FanoutAWS_3_io_out_3;
  assign MultiplyAccumulate_3_io_weights = delayWeights_3;
  assign MultiplyAccumulate_4_clock = clock;
  assign MultiplyAccumulate_4_io_activations_0 = FanoutAWS_io_out_4;
  assign MultiplyAccumulate_4_io_activations_1 = FanoutAWS_1_io_out_4;
  assign MultiplyAccumulate_4_io_activations_2 = FanoutAWS_2_io_out_4;
  assign MultiplyAccumulate_4_io_activations_3 = FanoutAWS_3_io_out_4;
  assign MultiplyAccumulate_4_io_weights = delayWeights_4;
  assign MultiplyAccumulate_5_clock = clock;
  assign MultiplyAccumulate_5_io_activations_0 = FanoutAWS_io_out_5;
  assign MultiplyAccumulate_5_io_activations_1 = FanoutAWS_1_io_out_5;
  assign MultiplyAccumulate_5_io_activations_2 = FanoutAWS_2_io_out_5;
  assign MultiplyAccumulate_5_io_activations_3 = FanoutAWS_3_io_out_5;
  assign MultiplyAccumulate_5_io_weights = delayWeights_5;
  assign MultiplyAccumulate_6_clock = clock;
  assign MultiplyAccumulate_6_io_activations_0 = FanoutAWS_io_out_6;
  assign MultiplyAccumulate_6_io_activations_1 = FanoutAWS_1_io_out_6;
  assign MultiplyAccumulate_6_io_activations_2 = FanoutAWS_2_io_out_6;
  assign MultiplyAccumulate_6_io_activations_3 = FanoutAWS_3_io_out_6;
  assign MultiplyAccumulate_6_io_weights = delayWeights_6;
  assign MultiplyAccumulate_7_clock = clock;
  assign MultiplyAccumulate_7_io_activations_0 = FanoutAWS_io_out_7;
  assign MultiplyAccumulate_7_io_activations_1 = FanoutAWS_1_io_out_7;
  assign MultiplyAccumulate_7_io_activations_2 = FanoutAWS_2_io_out_7;
  assign MultiplyAccumulate_7_io_activations_3 = FanoutAWS_3_io_out_7;
  assign MultiplyAccumulate_7_io_weights = delayWeights_7;
  assign MultiplyAccumulate_8_clock = clock;
  assign MultiplyAccumulate_8_io_activations_0 = FanoutAWS_io_out_8;
  assign MultiplyAccumulate_8_io_activations_1 = FanoutAWS_1_io_out_8;
  assign MultiplyAccumulate_8_io_activations_2 = FanoutAWS_2_io_out_8;
  assign MultiplyAccumulate_8_io_activations_3 = FanoutAWS_3_io_out_8;
  assign MultiplyAccumulate_8_io_weights = delayWeights_8;
  assign MultiplyAccumulate_9_clock = clock;
  assign MultiplyAccumulate_9_io_activations_0 = FanoutAWS_io_out_9;
  assign MultiplyAccumulate_9_io_activations_1 = FanoutAWS_1_io_out_9;
  assign MultiplyAccumulate_9_io_activations_2 = FanoutAWS_2_io_out_9;
  assign MultiplyAccumulate_9_io_activations_3 = FanoutAWS_3_io_out_9;
  assign MultiplyAccumulate_9_io_weights = delayWeights_9;
  assign MultiplyAccumulate_10_clock = clock;
  assign MultiplyAccumulate_10_io_activations_0 = FanoutAWS_io_out_10;
  assign MultiplyAccumulate_10_io_activations_1 = FanoutAWS_1_io_out_10;
  assign MultiplyAccumulate_10_io_activations_2 = FanoutAWS_2_io_out_10;
  assign MultiplyAccumulate_10_io_activations_3 = FanoutAWS_3_io_out_10;
  assign MultiplyAccumulate_10_io_weights = delayWeights_10;
  assign MultiplyAccumulate_11_clock = clock;
  assign MultiplyAccumulate_11_io_activations_0 = FanoutAWS_io_out_11;
  assign MultiplyAccumulate_11_io_activations_1 = FanoutAWS_1_io_out_11;
  assign MultiplyAccumulate_11_io_activations_2 = FanoutAWS_2_io_out_11;
  assign MultiplyAccumulate_11_io_activations_3 = FanoutAWS_3_io_out_11;
  assign MultiplyAccumulate_11_io_weights = delayWeights_11;
  assign MultiplyAccumulate_12_clock = clock;
  assign MultiplyAccumulate_12_io_activations_0 = FanoutAWS_io_out_12;
  assign MultiplyAccumulate_12_io_activations_1 = FanoutAWS_1_io_out_12;
  assign MultiplyAccumulate_12_io_activations_2 = FanoutAWS_2_io_out_12;
  assign MultiplyAccumulate_12_io_activations_3 = FanoutAWS_3_io_out_12;
  assign MultiplyAccumulate_12_io_weights = delayWeights_12;
  assign MultiplyAccumulate_13_clock = clock;
  assign MultiplyAccumulate_13_io_activations_0 = FanoutAWS_io_out_13;
  assign MultiplyAccumulate_13_io_activations_1 = FanoutAWS_1_io_out_13;
  assign MultiplyAccumulate_13_io_activations_2 = FanoutAWS_2_io_out_13;
  assign MultiplyAccumulate_13_io_activations_3 = FanoutAWS_3_io_out_13;
  assign MultiplyAccumulate_13_io_weights = delayWeights_13;
  assign MultiplyAccumulate_14_clock = clock;
  assign MultiplyAccumulate_14_io_activations_0 = FanoutAWS_io_out_14;
  assign MultiplyAccumulate_14_io_activations_1 = FanoutAWS_1_io_out_14;
  assign MultiplyAccumulate_14_io_activations_2 = FanoutAWS_2_io_out_14;
  assign MultiplyAccumulate_14_io_activations_3 = FanoutAWS_3_io_out_14;
  assign MultiplyAccumulate_14_io_weights = delayWeights_14;
  assign MultiplyAccumulate_15_clock = clock;
  assign MultiplyAccumulate_15_io_activations_0 = FanoutAWS_io_out_15;
  assign MultiplyAccumulate_15_io_activations_1 = FanoutAWS_1_io_out_15;
  assign MultiplyAccumulate_15_io_activations_2 = FanoutAWS_2_io_out_15;
  assign MultiplyAccumulate_15_io_activations_3 = FanoutAWS_3_io_out_15;
  assign MultiplyAccumulate_15_io_weights = delayWeights_15;
  assign MultiplyAccumulate_16_clock = clock;
  assign MultiplyAccumulate_16_io_activations_0 = FanoutAWS_io_out_16;
  assign MultiplyAccumulate_16_io_activations_1 = FanoutAWS_1_io_out_16;
  assign MultiplyAccumulate_16_io_activations_2 = FanoutAWS_2_io_out_16;
  assign MultiplyAccumulate_16_io_activations_3 = FanoutAWS_3_io_out_16;
  assign MultiplyAccumulate_16_io_weights = delayWeights_16;
  assign MultiplyAccumulate_17_clock = clock;
  assign MultiplyAccumulate_17_io_activations_0 = FanoutAWS_io_out_17;
  assign MultiplyAccumulate_17_io_activations_1 = FanoutAWS_1_io_out_17;
  assign MultiplyAccumulate_17_io_activations_2 = FanoutAWS_2_io_out_17;
  assign MultiplyAccumulate_17_io_activations_3 = FanoutAWS_3_io_out_17;
  assign MultiplyAccumulate_17_io_weights = delayWeights_17;
  assign MultiplyAccumulate_18_clock = clock;
  assign MultiplyAccumulate_18_io_activations_0 = FanoutAWS_io_out_18;
  assign MultiplyAccumulate_18_io_activations_1 = FanoutAWS_1_io_out_18;
  assign MultiplyAccumulate_18_io_activations_2 = FanoutAWS_2_io_out_18;
  assign MultiplyAccumulate_18_io_activations_3 = FanoutAWS_3_io_out_18;
  assign MultiplyAccumulate_18_io_weights = delayWeights_18;
  assign MultiplyAccumulate_19_clock = clock;
  assign MultiplyAccumulate_19_io_activations_0 = FanoutAWS_io_out_19;
  assign MultiplyAccumulate_19_io_activations_1 = FanoutAWS_1_io_out_19;
  assign MultiplyAccumulate_19_io_activations_2 = FanoutAWS_2_io_out_19;
  assign MultiplyAccumulate_19_io_activations_3 = FanoutAWS_3_io_out_19;
  assign MultiplyAccumulate_19_io_weights = delayWeights_19;
  assign MultiplyAccumulate_20_clock = clock;
  assign MultiplyAccumulate_20_io_activations_0 = FanoutAWS_io_out_20;
  assign MultiplyAccumulate_20_io_activations_1 = FanoutAWS_1_io_out_20;
  assign MultiplyAccumulate_20_io_activations_2 = FanoutAWS_2_io_out_20;
  assign MultiplyAccumulate_20_io_activations_3 = FanoutAWS_3_io_out_20;
  assign MultiplyAccumulate_20_io_weights = delayWeights_20;
  assign MultiplyAccumulate_21_clock = clock;
  assign MultiplyAccumulate_21_io_activations_0 = FanoutAWS_io_out_21;
  assign MultiplyAccumulate_21_io_activations_1 = FanoutAWS_1_io_out_21;
  assign MultiplyAccumulate_21_io_activations_2 = FanoutAWS_2_io_out_21;
  assign MultiplyAccumulate_21_io_activations_3 = FanoutAWS_3_io_out_21;
  assign MultiplyAccumulate_21_io_weights = delayWeights_21;
  assign MultiplyAccumulate_22_clock = clock;
  assign MultiplyAccumulate_22_io_activations_0 = FanoutAWS_io_out_22;
  assign MultiplyAccumulate_22_io_activations_1 = FanoutAWS_1_io_out_22;
  assign MultiplyAccumulate_22_io_activations_2 = FanoutAWS_2_io_out_22;
  assign MultiplyAccumulate_22_io_activations_3 = FanoutAWS_3_io_out_22;
  assign MultiplyAccumulate_22_io_weights = delayWeights_22;
  assign MultiplyAccumulate_23_clock = clock;
  assign MultiplyAccumulate_23_io_activations_0 = FanoutAWS_io_out_23;
  assign MultiplyAccumulate_23_io_activations_1 = FanoutAWS_1_io_out_23;
  assign MultiplyAccumulate_23_io_activations_2 = FanoutAWS_2_io_out_23;
  assign MultiplyAccumulate_23_io_activations_3 = FanoutAWS_3_io_out_23;
  assign MultiplyAccumulate_23_io_weights = delayWeights_23;
  assign MultiplyAccumulate_24_clock = clock;
  assign MultiplyAccumulate_24_io_activations_0 = FanoutAWS_io_out_24;
  assign MultiplyAccumulate_24_io_activations_1 = FanoutAWS_1_io_out_24;
  assign MultiplyAccumulate_24_io_activations_2 = FanoutAWS_2_io_out_24;
  assign MultiplyAccumulate_24_io_activations_3 = FanoutAWS_3_io_out_24;
  assign MultiplyAccumulate_24_io_weights = delayWeights_24;
  assign MultiplyAccumulate_25_clock = clock;
  assign MultiplyAccumulate_25_io_activations_0 = FanoutAWS_io_out_25;
  assign MultiplyAccumulate_25_io_activations_1 = FanoutAWS_1_io_out_25;
  assign MultiplyAccumulate_25_io_activations_2 = FanoutAWS_2_io_out_25;
  assign MultiplyAccumulate_25_io_activations_3 = FanoutAWS_3_io_out_25;
  assign MultiplyAccumulate_25_io_weights = delayWeights_25;
  assign MultiplyAccumulate_26_clock = clock;
  assign MultiplyAccumulate_26_io_activations_0 = FanoutAWS_io_out_26;
  assign MultiplyAccumulate_26_io_activations_1 = FanoutAWS_1_io_out_26;
  assign MultiplyAccumulate_26_io_activations_2 = FanoutAWS_2_io_out_26;
  assign MultiplyAccumulate_26_io_activations_3 = FanoutAWS_3_io_out_26;
  assign MultiplyAccumulate_26_io_weights = delayWeights_26;
  assign MultiplyAccumulate_27_clock = clock;
  assign MultiplyAccumulate_27_io_activations_0 = FanoutAWS_io_out_27;
  assign MultiplyAccumulate_27_io_activations_1 = FanoutAWS_1_io_out_27;
  assign MultiplyAccumulate_27_io_activations_2 = FanoutAWS_2_io_out_27;
  assign MultiplyAccumulate_27_io_activations_3 = FanoutAWS_3_io_out_27;
  assign MultiplyAccumulate_27_io_weights = delayWeights_27;
  assign MultiplyAccumulate_28_clock = clock;
  assign MultiplyAccumulate_28_io_activations_0 = FanoutAWS_io_out_28;
  assign MultiplyAccumulate_28_io_activations_1 = FanoutAWS_1_io_out_28;
  assign MultiplyAccumulate_28_io_activations_2 = FanoutAWS_2_io_out_28;
  assign MultiplyAccumulate_28_io_activations_3 = FanoutAWS_3_io_out_28;
  assign MultiplyAccumulate_28_io_weights = delayWeights_28;
  assign MultiplyAccumulate_29_clock = clock;
  assign MultiplyAccumulate_29_io_activations_0 = FanoutAWS_io_out_29;
  assign MultiplyAccumulate_29_io_activations_1 = FanoutAWS_1_io_out_29;
  assign MultiplyAccumulate_29_io_activations_2 = FanoutAWS_2_io_out_29;
  assign MultiplyAccumulate_29_io_activations_3 = FanoutAWS_3_io_out_29;
  assign MultiplyAccumulate_29_io_weights = delayWeights_29;
  assign MultiplyAccumulate_30_clock = clock;
  assign MultiplyAccumulate_30_io_activations_0 = FanoutAWS_io_out_30;
  assign MultiplyAccumulate_30_io_activations_1 = FanoutAWS_1_io_out_30;
  assign MultiplyAccumulate_30_io_activations_2 = FanoutAWS_2_io_out_30;
  assign MultiplyAccumulate_30_io_activations_3 = FanoutAWS_3_io_out_30;
  assign MultiplyAccumulate_30_io_weights = delayWeights_30;
  assign MultiplyAccumulate_31_clock = clock;
  assign MultiplyAccumulate_31_io_activations_0 = FanoutAWS_io_out_31;
  assign MultiplyAccumulate_31_io_activations_1 = FanoutAWS_1_io_out_31;
  assign MultiplyAccumulate_31_io_activations_2 = FanoutAWS_2_io_out_31;
  assign MultiplyAccumulate_31_io_activations_3 = FanoutAWS_3_io_out_31;
  assign MultiplyAccumulate_31_io_weights = delayWeights_31;
  assign MultiplyAccumulate_32_clock = clock;
  assign MultiplyAccumulate_32_io_activations_0 = FanoutAWS_io_out_32;
  assign MultiplyAccumulate_32_io_activations_1 = FanoutAWS_1_io_out_32;
  assign MultiplyAccumulate_32_io_activations_2 = FanoutAWS_2_io_out_32;
  assign MultiplyAccumulate_32_io_activations_3 = FanoutAWS_3_io_out_32;
  assign MultiplyAccumulate_32_io_weights = delayWeights_32;
  assign MultiplyAccumulate_33_clock = clock;
  assign MultiplyAccumulate_33_io_activations_0 = FanoutAWS_io_out_33;
  assign MultiplyAccumulate_33_io_activations_1 = FanoutAWS_1_io_out_33;
  assign MultiplyAccumulate_33_io_activations_2 = FanoutAWS_2_io_out_33;
  assign MultiplyAccumulate_33_io_activations_3 = FanoutAWS_3_io_out_33;
  assign MultiplyAccumulate_33_io_weights = delayWeights_33;
  assign MultiplyAccumulate_34_clock = clock;
  assign MultiplyAccumulate_34_io_activations_0 = FanoutAWS_io_out_34;
  assign MultiplyAccumulate_34_io_activations_1 = FanoutAWS_1_io_out_34;
  assign MultiplyAccumulate_34_io_activations_2 = FanoutAWS_2_io_out_34;
  assign MultiplyAccumulate_34_io_activations_3 = FanoutAWS_3_io_out_34;
  assign MultiplyAccumulate_34_io_weights = delayWeights_34;
  assign MultiplyAccumulate_35_clock = clock;
  assign MultiplyAccumulate_35_io_activations_0 = FanoutAWS_io_out_35;
  assign MultiplyAccumulate_35_io_activations_1 = FanoutAWS_1_io_out_35;
  assign MultiplyAccumulate_35_io_activations_2 = FanoutAWS_2_io_out_35;
  assign MultiplyAccumulate_35_io_activations_3 = FanoutAWS_3_io_out_35;
  assign MultiplyAccumulate_35_io_weights = delayWeights_35;
  assign MultiplyAccumulate_36_clock = clock;
  assign MultiplyAccumulate_36_io_activations_0 = FanoutAWS_io_out_36;
  assign MultiplyAccumulate_36_io_activations_1 = FanoutAWS_1_io_out_36;
  assign MultiplyAccumulate_36_io_activations_2 = FanoutAWS_2_io_out_36;
  assign MultiplyAccumulate_36_io_activations_3 = FanoutAWS_3_io_out_36;
  assign MultiplyAccumulate_36_io_weights = delayWeights_36;
  assign MultiplyAccumulate_37_clock = clock;
  assign MultiplyAccumulate_37_io_activations_0 = FanoutAWS_io_out_37;
  assign MultiplyAccumulate_37_io_activations_1 = FanoutAWS_1_io_out_37;
  assign MultiplyAccumulate_37_io_activations_2 = FanoutAWS_2_io_out_37;
  assign MultiplyAccumulate_37_io_activations_3 = FanoutAWS_3_io_out_37;
  assign MultiplyAccumulate_37_io_weights = delayWeights_37;
  assign MultiplyAccumulate_38_clock = clock;
  assign MultiplyAccumulate_38_io_activations_0 = FanoutAWS_io_out_38;
  assign MultiplyAccumulate_38_io_activations_1 = FanoutAWS_1_io_out_38;
  assign MultiplyAccumulate_38_io_activations_2 = FanoutAWS_2_io_out_38;
  assign MultiplyAccumulate_38_io_activations_3 = FanoutAWS_3_io_out_38;
  assign MultiplyAccumulate_38_io_weights = delayWeights_38;
  assign MultiplyAccumulate_39_clock = clock;
  assign MultiplyAccumulate_39_io_activations_0 = FanoutAWS_io_out_39;
  assign MultiplyAccumulate_39_io_activations_1 = FanoutAWS_1_io_out_39;
  assign MultiplyAccumulate_39_io_activations_2 = FanoutAWS_2_io_out_39;
  assign MultiplyAccumulate_39_io_activations_3 = FanoutAWS_3_io_out_39;
  assign MultiplyAccumulate_39_io_weights = delayWeights_39;
  assign MultiplyAccumulate_40_clock = clock;
  assign MultiplyAccumulate_40_io_activations_0 = FanoutAWS_io_out_40;
  assign MultiplyAccumulate_40_io_activations_1 = FanoutAWS_1_io_out_40;
  assign MultiplyAccumulate_40_io_activations_2 = FanoutAWS_2_io_out_40;
  assign MultiplyAccumulate_40_io_activations_3 = FanoutAWS_3_io_out_40;
  assign MultiplyAccumulate_40_io_weights = delayWeights_40;
  assign MultiplyAccumulate_41_clock = clock;
  assign MultiplyAccumulate_41_io_activations_0 = FanoutAWS_io_out_41;
  assign MultiplyAccumulate_41_io_activations_1 = FanoutAWS_1_io_out_41;
  assign MultiplyAccumulate_41_io_activations_2 = FanoutAWS_2_io_out_41;
  assign MultiplyAccumulate_41_io_activations_3 = FanoutAWS_3_io_out_41;
  assign MultiplyAccumulate_41_io_weights = delayWeights_41;
  assign MultiplyAccumulate_42_clock = clock;
  assign MultiplyAccumulate_42_io_activations_0 = FanoutAWS_io_out_42;
  assign MultiplyAccumulate_42_io_activations_1 = FanoutAWS_1_io_out_42;
  assign MultiplyAccumulate_42_io_activations_2 = FanoutAWS_2_io_out_42;
  assign MultiplyAccumulate_42_io_activations_3 = FanoutAWS_3_io_out_42;
  assign MultiplyAccumulate_42_io_weights = delayWeights_42;
  assign MultiplyAccumulate_43_clock = clock;
  assign MultiplyAccumulate_43_io_activations_0 = FanoutAWS_io_out_43;
  assign MultiplyAccumulate_43_io_activations_1 = FanoutAWS_1_io_out_43;
  assign MultiplyAccumulate_43_io_activations_2 = FanoutAWS_2_io_out_43;
  assign MultiplyAccumulate_43_io_activations_3 = FanoutAWS_3_io_out_43;
  assign MultiplyAccumulate_43_io_weights = delayWeights_43;
  assign MultiplyAccumulate_44_clock = clock;
  assign MultiplyAccumulate_44_io_activations_0 = FanoutAWS_io_out_44;
  assign MultiplyAccumulate_44_io_activations_1 = FanoutAWS_1_io_out_44;
  assign MultiplyAccumulate_44_io_activations_2 = FanoutAWS_2_io_out_44;
  assign MultiplyAccumulate_44_io_activations_3 = FanoutAWS_3_io_out_44;
  assign MultiplyAccumulate_44_io_weights = delayWeights_44;
  assign MultiplyAccumulate_45_clock = clock;
  assign MultiplyAccumulate_45_io_activations_0 = FanoutAWS_io_out_45;
  assign MultiplyAccumulate_45_io_activations_1 = FanoutAWS_1_io_out_45;
  assign MultiplyAccumulate_45_io_activations_2 = FanoutAWS_2_io_out_45;
  assign MultiplyAccumulate_45_io_activations_3 = FanoutAWS_3_io_out_45;
  assign MultiplyAccumulate_45_io_weights = delayWeights_45;
  assign MultiplyAccumulate_46_clock = clock;
  assign MultiplyAccumulate_46_io_activations_0 = FanoutAWS_io_out_46;
  assign MultiplyAccumulate_46_io_activations_1 = FanoutAWS_1_io_out_46;
  assign MultiplyAccumulate_46_io_activations_2 = FanoutAWS_2_io_out_46;
  assign MultiplyAccumulate_46_io_activations_3 = FanoutAWS_3_io_out_46;
  assign MultiplyAccumulate_46_io_weights = delayWeights_46;
  assign MultiplyAccumulate_47_clock = clock;
  assign MultiplyAccumulate_47_io_activations_0 = FanoutAWS_io_out_47;
  assign MultiplyAccumulate_47_io_activations_1 = FanoutAWS_1_io_out_47;
  assign MultiplyAccumulate_47_io_activations_2 = FanoutAWS_2_io_out_47;
  assign MultiplyAccumulate_47_io_activations_3 = FanoutAWS_3_io_out_47;
  assign MultiplyAccumulate_47_io_weights = delayWeights_47;
  assign MultiplyAccumulate_48_clock = clock;
  assign MultiplyAccumulate_48_io_activations_0 = FanoutAWS_io_out_48;
  assign MultiplyAccumulate_48_io_activations_1 = FanoutAWS_1_io_out_48;
  assign MultiplyAccumulate_48_io_activations_2 = FanoutAWS_2_io_out_48;
  assign MultiplyAccumulate_48_io_activations_3 = FanoutAWS_3_io_out_48;
  assign MultiplyAccumulate_48_io_weights = delayWeights_48;
  assign MultiplyAccumulate_49_clock = clock;
  assign MultiplyAccumulate_49_io_activations_0 = FanoutAWS_io_out_49;
  assign MultiplyAccumulate_49_io_activations_1 = FanoutAWS_1_io_out_49;
  assign MultiplyAccumulate_49_io_activations_2 = FanoutAWS_2_io_out_49;
  assign MultiplyAccumulate_49_io_activations_3 = FanoutAWS_3_io_out_49;
  assign MultiplyAccumulate_49_io_weights = delayWeights_49;
  assign MultiplyAccumulate_50_clock = clock;
  assign MultiplyAccumulate_50_io_activations_0 = FanoutAWS_io_out_50;
  assign MultiplyAccumulate_50_io_activations_1 = FanoutAWS_1_io_out_50;
  assign MultiplyAccumulate_50_io_activations_2 = FanoutAWS_2_io_out_50;
  assign MultiplyAccumulate_50_io_activations_3 = FanoutAWS_3_io_out_50;
  assign MultiplyAccumulate_50_io_weights = delayWeights_50;
  assign MultiplyAccumulate_51_clock = clock;
  assign MultiplyAccumulate_51_io_activations_0 = FanoutAWS_io_out_51;
  assign MultiplyAccumulate_51_io_activations_1 = FanoutAWS_1_io_out_51;
  assign MultiplyAccumulate_51_io_activations_2 = FanoutAWS_2_io_out_51;
  assign MultiplyAccumulate_51_io_activations_3 = FanoutAWS_3_io_out_51;
  assign MultiplyAccumulate_51_io_weights = delayWeights_51;
  assign MultiplyAccumulate_52_clock = clock;
  assign MultiplyAccumulate_52_io_activations_0 = FanoutAWS_io_out_52;
  assign MultiplyAccumulate_52_io_activations_1 = FanoutAWS_1_io_out_52;
  assign MultiplyAccumulate_52_io_activations_2 = FanoutAWS_2_io_out_52;
  assign MultiplyAccumulate_52_io_activations_3 = FanoutAWS_3_io_out_52;
  assign MultiplyAccumulate_52_io_weights = delayWeights_52;
  assign MultiplyAccumulate_53_clock = clock;
  assign MultiplyAccumulate_53_io_activations_0 = FanoutAWS_io_out_53;
  assign MultiplyAccumulate_53_io_activations_1 = FanoutAWS_1_io_out_53;
  assign MultiplyAccumulate_53_io_activations_2 = FanoutAWS_2_io_out_53;
  assign MultiplyAccumulate_53_io_activations_3 = FanoutAWS_3_io_out_53;
  assign MultiplyAccumulate_53_io_weights = delayWeights_53;
  assign MultiplyAccumulate_54_clock = clock;
  assign MultiplyAccumulate_54_io_activations_0 = FanoutAWS_io_out_54;
  assign MultiplyAccumulate_54_io_activations_1 = FanoutAWS_1_io_out_54;
  assign MultiplyAccumulate_54_io_activations_2 = FanoutAWS_2_io_out_54;
  assign MultiplyAccumulate_54_io_activations_3 = FanoutAWS_3_io_out_54;
  assign MultiplyAccumulate_54_io_weights = delayWeights_54;
  assign MultiplyAccumulate_55_clock = clock;
  assign MultiplyAccumulate_55_io_activations_0 = FanoutAWS_io_out_55;
  assign MultiplyAccumulate_55_io_activations_1 = FanoutAWS_1_io_out_55;
  assign MultiplyAccumulate_55_io_activations_2 = FanoutAWS_2_io_out_55;
  assign MultiplyAccumulate_55_io_activations_3 = FanoutAWS_3_io_out_55;
  assign MultiplyAccumulate_55_io_weights = delayWeights_55;
  assign MultiplyAccumulate_56_clock = clock;
  assign MultiplyAccumulate_56_io_activations_0 = FanoutAWS_io_out_56;
  assign MultiplyAccumulate_56_io_activations_1 = FanoutAWS_1_io_out_56;
  assign MultiplyAccumulate_56_io_activations_2 = FanoutAWS_2_io_out_56;
  assign MultiplyAccumulate_56_io_activations_3 = FanoutAWS_3_io_out_56;
  assign MultiplyAccumulate_56_io_weights = delayWeights_56;
  assign MultiplyAccumulate_57_clock = clock;
  assign MultiplyAccumulate_57_io_activations_0 = FanoutAWS_io_out_57;
  assign MultiplyAccumulate_57_io_activations_1 = FanoutAWS_1_io_out_57;
  assign MultiplyAccumulate_57_io_activations_2 = FanoutAWS_2_io_out_57;
  assign MultiplyAccumulate_57_io_activations_3 = FanoutAWS_3_io_out_57;
  assign MultiplyAccumulate_57_io_weights = delayWeights_57;
  assign MultiplyAccumulate_58_clock = clock;
  assign MultiplyAccumulate_58_io_activations_0 = FanoutAWS_io_out_58;
  assign MultiplyAccumulate_58_io_activations_1 = FanoutAWS_1_io_out_58;
  assign MultiplyAccumulate_58_io_activations_2 = FanoutAWS_2_io_out_58;
  assign MultiplyAccumulate_58_io_activations_3 = FanoutAWS_3_io_out_58;
  assign MultiplyAccumulate_58_io_weights = delayWeights_58;
  assign MultiplyAccumulate_59_clock = clock;
  assign MultiplyAccumulate_59_io_activations_0 = FanoutAWS_io_out_59;
  assign MultiplyAccumulate_59_io_activations_1 = FanoutAWS_1_io_out_59;
  assign MultiplyAccumulate_59_io_activations_2 = FanoutAWS_2_io_out_59;
  assign MultiplyAccumulate_59_io_activations_3 = FanoutAWS_3_io_out_59;
  assign MultiplyAccumulate_59_io_weights = delayWeights_59;
  assign MultiplyAccumulate_60_clock = clock;
  assign MultiplyAccumulate_60_io_activations_0 = FanoutAWS_io_out_60;
  assign MultiplyAccumulate_60_io_activations_1 = FanoutAWS_1_io_out_60;
  assign MultiplyAccumulate_60_io_activations_2 = FanoutAWS_2_io_out_60;
  assign MultiplyAccumulate_60_io_activations_3 = FanoutAWS_3_io_out_60;
  assign MultiplyAccumulate_60_io_weights = delayWeights_60;
  assign MultiplyAccumulate_61_clock = clock;
  assign MultiplyAccumulate_61_io_activations_0 = FanoutAWS_io_out_61;
  assign MultiplyAccumulate_61_io_activations_1 = FanoutAWS_1_io_out_61;
  assign MultiplyAccumulate_61_io_activations_2 = FanoutAWS_2_io_out_61;
  assign MultiplyAccumulate_61_io_activations_3 = FanoutAWS_3_io_out_61;
  assign MultiplyAccumulate_61_io_weights = delayWeights_61;
  assign MultiplyAccumulate_62_clock = clock;
  assign MultiplyAccumulate_62_io_activations_0 = FanoutAWS_io_out_62;
  assign MultiplyAccumulate_62_io_activations_1 = FanoutAWS_1_io_out_62;
  assign MultiplyAccumulate_62_io_activations_2 = FanoutAWS_2_io_out_62;
  assign MultiplyAccumulate_62_io_activations_3 = FanoutAWS_3_io_out_62;
  assign MultiplyAccumulate_62_io_weights = delayWeights_62;
  assign MultiplyAccumulate_63_clock = clock;
  assign MultiplyAccumulate_63_io_activations_0 = FanoutAWS_io_out_63;
  assign MultiplyAccumulate_63_io_activations_1 = FanoutAWS_1_io_out_63;
  assign MultiplyAccumulate_63_io_activations_2 = FanoutAWS_2_io_out_63;
  assign MultiplyAccumulate_63_io_activations_3 = FanoutAWS_3_io_out_63;
  assign MultiplyAccumulate_63_io_weights = delayWeights_63;
  assign MultiplyAccumulate_64_clock = clock;
  assign MultiplyAccumulate_64_io_activations_0 = FanoutAWS_io_out_64;
  assign MultiplyAccumulate_64_io_activations_1 = FanoutAWS_1_io_out_64;
  assign MultiplyAccumulate_64_io_activations_2 = FanoutAWS_2_io_out_64;
  assign MultiplyAccumulate_64_io_activations_3 = FanoutAWS_3_io_out_64;
  assign MultiplyAccumulate_64_io_weights = delayWeights_64;
  assign MultiplyAccumulate_65_clock = clock;
  assign MultiplyAccumulate_65_io_activations_0 = FanoutAWS_io_out_65;
  assign MultiplyAccumulate_65_io_activations_1 = FanoutAWS_1_io_out_65;
  assign MultiplyAccumulate_65_io_activations_2 = FanoutAWS_2_io_out_65;
  assign MultiplyAccumulate_65_io_activations_3 = FanoutAWS_3_io_out_65;
  assign MultiplyAccumulate_65_io_weights = delayWeights_65;
  assign MultiplyAccumulate_66_clock = clock;
  assign MultiplyAccumulate_66_io_activations_0 = FanoutAWS_io_out_66;
  assign MultiplyAccumulate_66_io_activations_1 = FanoutAWS_1_io_out_66;
  assign MultiplyAccumulate_66_io_activations_2 = FanoutAWS_2_io_out_66;
  assign MultiplyAccumulate_66_io_activations_3 = FanoutAWS_3_io_out_66;
  assign MultiplyAccumulate_66_io_weights = delayWeights_66;
  assign MultiplyAccumulate_67_clock = clock;
  assign MultiplyAccumulate_67_io_activations_0 = FanoutAWS_io_out_67;
  assign MultiplyAccumulate_67_io_activations_1 = FanoutAWS_1_io_out_67;
  assign MultiplyAccumulate_67_io_activations_2 = FanoutAWS_2_io_out_67;
  assign MultiplyAccumulate_67_io_activations_3 = FanoutAWS_3_io_out_67;
  assign MultiplyAccumulate_67_io_weights = delayWeights_67;
  assign MultiplyAccumulate_68_clock = clock;
  assign MultiplyAccumulate_68_io_activations_0 = FanoutAWS_io_out_68;
  assign MultiplyAccumulate_68_io_activations_1 = FanoutAWS_1_io_out_68;
  assign MultiplyAccumulate_68_io_activations_2 = FanoutAWS_2_io_out_68;
  assign MultiplyAccumulate_68_io_activations_3 = FanoutAWS_3_io_out_68;
  assign MultiplyAccumulate_68_io_weights = delayWeights_68;
  assign MultiplyAccumulate_69_clock = clock;
  assign MultiplyAccumulate_69_io_activations_0 = FanoutAWS_io_out_69;
  assign MultiplyAccumulate_69_io_activations_1 = FanoutAWS_1_io_out_69;
  assign MultiplyAccumulate_69_io_activations_2 = FanoutAWS_2_io_out_69;
  assign MultiplyAccumulate_69_io_activations_3 = FanoutAWS_3_io_out_69;
  assign MultiplyAccumulate_69_io_weights = delayWeights_69;
  assign MultiplyAccumulate_70_clock = clock;
  assign MultiplyAccumulate_70_io_activations_0 = FanoutAWS_io_out_70;
  assign MultiplyAccumulate_70_io_activations_1 = FanoutAWS_1_io_out_70;
  assign MultiplyAccumulate_70_io_activations_2 = FanoutAWS_2_io_out_70;
  assign MultiplyAccumulate_70_io_activations_3 = FanoutAWS_3_io_out_70;
  assign MultiplyAccumulate_70_io_weights = delayWeights_70;
  assign MultiplyAccumulate_71_clock = clock;
  assign MultiplyAccumulate_71_io_activations_0 = FanoutAWS_io_out_71;
  assign MultiplyAccumulate_71_io_activations_1 = FanoutAWS_1_io_out_71;
  assign MultiplyAccumulate_71_io_activations_2 = FanoutAWS_2_io_out_71;
  assign MultiplyAccumulate_71_io_activations_3 = FanoutAWS_3_io_out_71;
  assign MultiplyAccumulate_71_io_weights = delayWeights_71;
  assign MultiplyAccumulate_72_clock = clock;
  assign MultiplyAccumulate_72_io_activations_0 = FanoutAWS_io_out_72;
  assign MultiplyAccumulate_72_io_activations_1 = FanoutAWS_1_io_out_72;
  assign MultiplyAccumulate_72_io_activations_2 = FanoutAWS_2_io_out_72;
  assign MultiplyAccumulate_72_io_activations_3 = FanoutAWS_3_io_out_72;
  assign MultiplyAccumulate_72_io_weights = delayWeights_72;
  assign MultiplyAccumulate_73_clock = clock;
  assign MultiplyAccumulate_73_io_activations_0 = FanoutAWS_io_out_73;
  assign MultiplyAccumulate_73_io_activations_1 = FanoutAWS_1_io_out_73;
  assign MultiplyAccumulate_73_io_activations_2 = FanoutAWS_2_io_out_73;
  assign MultiplyAccumulate_73_io_activations_3 = FanoutAWS_3_io_out_73;
  assign MultiplyAccumulate_73_io_weights = delayWeights_73;
  assign MultiplyAccumulate_74_clock = clock;
  assign MultiplyAccumulate_74_io_activations_0 = FanoutAWS_io_out_74;
  assign MultiplyAccumulate_74_io_activations_1 = FanoutAWS_1_io_out_74;
  assign MultiplyAccumulate_74_io_activations_2 = FanoutAWS_2_io_out_74;
  assign MultiplyAccumulate_74_io_activations_3 = FanoutAWS_3_io_out_74;
  assign MultiplyAccumulate_74_io_weights = delayWeights_74;
  assign MultiplyAccumulate_75_clock = clock;
  assign MultiplyAccumulate_75_io_activations_0 = FanoutAWS_io_out_75;
  assign MultiplyAccumulate_75_io_activations_1 = FanoutAWS_1_io_out_75;
  assign MultiplyAccumulate_75_io_activations_2 = FanoutAWS_2_io_out_75;
  assign MultiplyAccumulate_75_io_activations_3 = FanoutAWS_3_io_out_75;
  assign MultiplyAccumulate_75_io_weights = delayWeights_75;
  assign MultiplyAccumulate_76_clock = clock;
  assign MultiplyAccumulate_76_io_activations_0 = FanoutAWS_io_out_76;
  assign MultiplyAccumulate_76_io_activations_1 = FanoutAWS_1_io_out_76;
  assign MultiplyAccumulate_76_io_activations_2 = FanoutAWS_2_io_out_76;
  assign MultiplyAccumulate_76_io_activations_3 = FanoutAWS_3_io_out_76;
  assign MultiplyAccumulate_76_io_weights = delayWeights_76;
  assign MultiplyAccumulate_77_clock = clock;
  assign MultiplyAccumulate_77_io_activations_0 = FanoutAWS_io_out_77;
  assign MultiplyAccumulate_77_io_activations_1 = FanoutAWS_1_io_out_77;
  assign MultiplyAccumulate_77_io_activations_2 = FanoutAWS_2_io_out_77;
  assign MultiplyAccumulate_77_io_activations_3 = FanoutAWS_3_io_out_77;
  assign MultiplyAccumulate_77_io_weights = delayWeights_77;
  assign MultiplyAccumulate_78_clock = clock;
  assign MultiplyAccumulate_78_io_activations_0 = FanoutAWS_io_out_78;
  assign MultiplyAccumulate_78_io_activations_1 = FanoutAWS_1_io_out_78;
  assign MultiplyAccumulate_78_io_activations_2 = FanoutAWS_2_io_out_78;
  assign MultiplyAccumulate_78_io_activations_3 = FanoutAWS_3_io_out_78;
  assign MultiplyAccumulate_78_io_weights = delayWeights_78;
  assign MultiplyAccumulate_79_clock = clock;
  assign MultiplyAccumulate_79_io_activations_0 = FanoutAWS_io_out_79;
  assign MultiplyAccumulate_79_io_activations_1 = FanoutAWS_1_io_out_79;
  assign MultiplyAccumulate_79_io_activations_2 = FanoutAWS_2_io_out_79;
  assign MultiplyAccumulate_79_io_activations_3 = FanoutAWS_3_io_out_79;
  assign MultiplyAccumulate_79_io_weights = delayWeights_79;
  assign MultiplyAccumulate_80_clock = clock;
  assign MultiplyAccumulate_80_io_activations_0 = FanoutAWS_io_out_80;
  assign MultiplyAccumulate_80_io_activations_1 = FanoutAWS_1_io_out_80;
  assign MultiplyAccumulate_80_io_activations_2 = FanoutAWS_2_io_out_80;
  assign MultiplyAccumulate_80_io_activations_3 = FanoutAWS_3_io_out_80;
  assign MultiplyAccumulate_80_io_weights = delayWeights_80;
  assign MultiplyAccumulate_81_clock = clock;
  assign MultiplyAccumulate_81_io_activations_0 = FanoutAWS_io_out_81;
  assign MultiplyAccumulate_81_io_activations_1 = FanoutAWS_1_io_out_81;
  assign MultiplyAccumulate_81_io_activations_2 = FanoutAWS_2_io_out_81;
  assign MultiplyAccumulate_81_io_activations_3 = FanoutAWS_3_io_out_81;
  assign MultiplyAccumulate_81_io_weights = delayWeights_81;
  assign MultiplyAccumulate_82_clock = clock;
  assign MultiplyAccumulate_82_io_activations_0 = FanoutAWS_io_out_82;
  assign MultiplyAccumulate_82_io_activations_1 = FanoutAWS_1_io_out_82;
  assign MultiplyAccumulate_82_io_activations_2 = FanoutAWS_2_io_out_82;
  assign MultiplyAccumulate_82_io_activations_3 = FanoutAWS_3_io_out_82;
  assign MultiplyAccumulate_82_io_weights = delayWeights_82;
  assign MultiplyAccumulate_83_clock = clock;
  assign MultiplyAccumulate_83_io_activations_0 = FanoutAWS_io_out_83;
  assign MultiplyAccumulate_83_io_activations_1 = FanoutAWS_1_io_out_83;
  assign MultiplyAccumulate_83_io_activations_2 = FanoutAWS_2_io_out_83;
  assign MultiplyAccumulate_83_io_activations_3 = FanoutAWS_3_io_out_83;
  assign MultiplyAccumulate_83_io_weights = delayWeights_83;
  assign MultiplyAccumulate_84_clock = clock;
  assign MultiplyAccumulate_84_io_activations_0 = FanoutAWS_io_out_84;
  assign MultiplyAccumulate_84_io_activations_1 = FanoutAWS_1_io_out_84;
  assign MultiplyAccumulate_84_io_activations_2 = FanoutAWS_2_io_out_84;
  assign MultiplyAccumulate_84_io_activations_3 = FanoutAWS_3_io_out_84;
  assign MultiplyAccumulate_84_io_weights = delayWeights_84;
  assign MultiplyAccumulate_85_clock = clock;
  assign MultiplyAccumulate_85_io_activations_0 = FanoutAWS_io_out_85;
  assign MultiplyAccumulate_85_io_activations_1 = FanoutAWS_1_io_out_85;
  assign MultiplyAccumulate_85_io_activations_2 = FanoutAWS_2_io_out_85;
  assign MultiplyAccumulate_85_io_activations_3 = FanoutAWS_3_io_out_85;
  assign MultiplyAccumulate_85_io_weights = delayWeights_85;
  assign MultiplyAccumulate_86_clock = clock;
  assign MultiplyAccumulate_86_io_activations_0 = FanoutAWS_io_out_86;
  assign MultiplyAccumulate_86_io_activations_1 = FanoutAWS_1_io_out_86;
  assign MultiplyAccumulate_86_io_activations_2 = FanoutAWS_2_io_out_86;
  assign MultiplyAccumulate_86_io_activations_3 = FanoutAWS_3_io_out_86;
  assign MultiplyAccumulate_86_io_weights = delayWeights_86;
  assign MultiplyAccumulate_87_clock = clock;
  assign MultiplyAccumulate_87_io_activations_0 = FanoutAWS_io_out_87;
  assign MultiplyAccumulate_87_io_activations_1 = FanoutAWS_1_io_out_87;
  assign MultiplyAccumulate_87_io_activations_2 = FanoutAWS_2_io_out_87;
  assign MultiplyAccumulate_87_io_activations_3 = FanoutAWS_3_io_out_87;
  assign MultiplyAccumulate_87_io_weights = delayWeights_87;
  assign MultiplyAccumulate_88_clock = clock;
  assign MultiplyAccumulate_88_io_activations_0 = FanoutAWS_io_out_88;
  assign MultiplyAccumulate_88_io_activations_1 = FanoutAWS_1_io_out_88;
  assign MultiplyAccumulate_88_io_activations_2 = FanoutAWS_2_io_out_88;
  assign MultiplyAccumulate_88_io_activations_3 = FanoutAWS_3_io_out_88;
  assign MultiplyAccumulate_88_io_weights = delayWeights_88;
  assign MultiplyAccumulate_89_clock = clock;
  assign MultiplyAccumulate_89_io_activations_0 = FanoutAWS_io_out_89;
  assign MultiplyAccumulate_89_io_activations_1 = FanoutAWS_1_io_out_89;
  assign MultiplyAccumulate_89_io_activations_2 = FanoutAWS_2_io_out_89;
  assign MultiplyAccumulate_89_io_activations_3 = FanoutAWS_3_io_out_89;
  assign MultiplyAccumulate_89_io_weights = delayWeights_89;
  assign MultiplyAccumulate_90_clock = clock;
  assign MultiplyAccumulate_90_io_activations_0 = FanoutAWS_io_out_90;
  assign MultiplyAccumulate_90_io_activations_1 = FanoutAWS_1_io_out_90;
  assign MultiplyAccumulate_90_io_activations_2 = FanoutAWS_2_io_out_90;
  assign MultiplyAccumulate_90_io_activations_3 = FanoutAWS_3_io_out_90;
  assign MultiplyAccumulate_90_io_weights = delayWeights_90;
  assign MultiplyAccumulate_91_clock = clock;
  assign MultiplyAccumulate_91_io_activations_0 = FanoutAWS_io_out_91;
  assign MultiplyAccumulate_91_io_activations_1 = FanoutAWS_1_io_out_91;
  assign MultiplyAccumulate_91_io_activations_2 = FanoutAWS_2_io_out_91;
  assign MultiplyAccumulate_91_io_activations_3 = FanoutAWS_3_io_out_91;
  assign MultiplyAccumulate_91_io_weights = delayWeights_91;
  assign MultiplyAccumulate_92_clock = clock;
  assign MultiplyAccumulate_92_io_activations_0 = FanoutAWS_io_out_92;
  assign MultiplyAccumulate_92_io_activations_1 = FanoutAWS_1_io_out_92;
  assign MultiplyAccumulate_92_io_activations_2 = FanoutAWS_2_io_out_92;
  assign MultiplyAccumulate_92_io_activations_3 = FanoutAWS_3_io_out_92;
  assign MultiplyAccumulate_92_io_weights = delayWeights_92;
  assign MultiplyAccumulate_93_clock = clock;
  assign MultiplyAccumulate_93_io_activations_0 = FanoutAWS_io_out_93;
  assign MultiplyAccumulate_93_io_activations_1 = FanoutAWS_1_io_out_93;
  assign MultiplyAccumulate_93_io_activations_2 = FanoutAWS_2_io_out_93;
  assign MultiplyAccumulate_93_io_activations_3 = FanoutAWS_3_io_out_93;
  assign MultiplyAccumulate_93_io_weights = delayWeights_93;
  assign MultiplyAccumulate_94_clock = clock;
  assign MultiplyAccumulate_94_io_activations_0 = FanoutAWS_io_out_94;
  assign MultiplyAccumulate_94_io_activations_1 = FanoutAWS_1_io_out_94;
  assign MultiplyAccumulate_94_io_activations_2 = FanoutAWS_2_io_out_94;
  assign MultiplyAccumulate_94_io_activations_3 = FanoutAWS_3_io_out_94;
  assign MultiplyAccumulate_94_io_weights = delayWeights_94;
  assign MultiplyAccumulate_95_clock = clock;
  assign MultiplyAccumulate_95_io_activations_0 = FanoutAWS_io_out_95;
  assign MultiplyAccumulate_95_io_activations_1 = FanoutAWS_1_io_out_95;
  assign MultiplyAccumulate_95_io_activations_2 = FanoutAWS_2_io_out_95;
  assign MultiplyAccumulate_95_io_activations_3 = FanoutAWS_3_io_out_95;
  assign MultiplyAccumulate_95_io_weights = delayWeights_95;
  assign MultiplyAccumulate_96_clock = clock;
  assign MultiplyAccumulate_96_io_activations_0 = FanoutAWS_io_out_96;
  assign MultiplyAccumulate_96_io_activations_1 = FanoutAWS_1_io_out_96;
  assign MultiplyAccumulate_96_io_activations_2 = FanoutAWS_2_io_out_96;
  assign MultiplyAccumulate_96_io_activations_3 = FanoutAWS_3_io_out_96;
  assign MultiplyAccumulate_96_io_weights = delayWeights_96;
  assign MultiplyAccumulate_97_clock = clock;
  assign MultiplyAccumulate_97_io_activations_0 = FanoutAWS_io_out_97;
  assign MultiplyAccumulate_97_io_activations_1 = FanoutAWS_1_io_out_97;
  assign MultiplyAccumulate_97_io_activations_2 = FanoutAWS_2_io_out_97;
  assign MultiplyAccumulate_97_io_activations_3 = FanoutAWS_3_io_out_97;
  assign MultiplyAccumulate_97_io_weights = delayWeights_97;
  assign MultiplyAccumulate_98_clock = clock;
  assign MultiplyAccumulate_98_io_activations_0 = FanoutAWS_io_out_98;
  assign MultiplyAccumulate_98_io_activations_1 = FanoutAWS_1_io_out_98;
  assign MultiplyAccumulate_98_io_activations_2 = FanoutAWS_2_io_out_98;
  assign MultiplyAccumulate_98_io_activations_3 = FanoutAWS_3_io_out_98;
  assign MultiplyAccumulate_98_io_weights = delayWeights_98;
  assign MultiplyAccumulate_99_clock = clock;
  assign MultiplyAccumulate_99_io_activations_0 = FanoutAWS_io_out_99;
  assign MultiplyAccumulate_99_io_activations_1 = FanoutAWS_1_io_out_99;
  assign MultiplyAccumulate_99_io_activations_2 = FanoutAWS_2_io_out_99;
  assign MultiplyAccumulate_99_io_activations_3 = FanoutAWS_3_io_out_99;
  assign MultiplyAccumulate_99_io_weights = delayWeights_99;
  assign MultiplyAccumulate_100_clock = clock;
  assign MultiplyAccumulate_100_io_activations_0 = FanoutAWS_io_out_100;
  assign MultiplyAccumulate_100_io_activations_1 = FanoutAWS_1_io_out_100;
  assign MultiplyAccumulate_100_io_activations_2 = FanoutAWS_2_io_out_100;
  assign MultiplyAccumulate_100_io_activations_3 = FanoutAWS_3_io_out_100;
  assign MultiplyAccumulate_100_io_weights = delayWeights_100;
  assign MultiplyAccumulate_101_clock = clock;
  assign MultiplyAccumulate_101_io_activations_0 = FanoutAWS_io_out_101;
  assign MultiplyAccumulate_101_io_activations_1 = FanoutAWS_1_io_out_101;
  assign MultiplyAccumulate_101_io_activations_2 = FanoutAWS_2_io_out_101;
  assign MultiplyAccumulate_101_io_activations_3 = FanoutAWS_3_io_out_101;
  assign MultiplyAccumulate_101_io_weights = delayWeights_101;
  assign MultiplyAccumulate_102_clock = clock;
  assign MultiplyAccumulate_102_io_activations_0 = FanoutAWS_io_out_102;
  assign MultiplyAccumulate_102_io_activations_1 = FanoutAWS_1_io_out_102;
  assign MultiplyAccumulate_102_io_activations_2 = FanoutAWS_2_io_out_102;
  assign MultiplyAccumulate_102_io_activations_3 = FanoutAWS_3_io_out_102;
  assign MultiplyAccumulate_102_io_weights = delayWeights_102;
  assign MultiplyAccumulate_103_clock = clock;
  assign MultiplyAccumulate_103_io_activations_0 = FanoutAWS_io_out_103;
  assign MultiplyAccumulate_103_io_activations_1 = FanoutAWS_1_io_out_103;
  assign MultiplyAccumulate_103_io_activations_2 = FanoutAWS_2_io_out_103;
  assign MultiplyAccumulate_103_io_activations_3 = FanoutAWS_3_io_out_103;
  assign MultiplyAccumulate_103_io_weights = delayWeights_103;
  assign MultiplyAccumulate_104_clock = clock;
  assign MultiplyAccumulate_104_io_activations_0 = FanoutAWS_io_out_104;
  assign MultiplyAccumulate_104_io_activations_1 = FanoutAWS_1_io_out_104;
  assign MultiplyAccumulate_104_io_activations_2 = FanoutAWS_2_io_out_104;
  assign MultiplyAccumulate_104_io_activations_3 = FanoutAWS_3_io_out_104;
  assign MultiplyAccumulate_104_io_weights = delayWeights_104;
  assign MultiplyAccumulate_105_clock = clock;
  assign MultiplyAccumulate_105_io_activations_0 = FanoutAWS_io_out_105;
  assign MultiplyAccumulate_105_io_activations_1 = FanoutAWS_1_io_out_105;
  assign MultiplyAccumulate_105_io_activations_2 = FanoutAWS_2_io_out_105;
  assign MultiplyAccumulate_105_io_activations_3 = FanoutAWS_3_io_out_105;
  assign MultiplyAccumulate_105_io_weights = delayWeights_105;
  assign MultiplyAccumulate_106_clock = clock;
  assign MultiplyAccumulate_106_io_activations_0 = FanoutAWS_io_out_106;
  assign MultiplyAccumulate_106_io_activations_1 = FanoutAWS_1_io_out_106;
  assign MultiplyAccumulate_106_io_activations_2 = FanoutAWS_2_io_out_106;
  assign MultiplyAccumulate_106_io_activations_3 = FanoutAWS_3_io_out_106;
  assign MultiplyAccumulate_106_io_weights = delayWeights_106;
  assign MultiplyAccumulate_107_clock = clock;
  assign MultiplyAccumulate_107_io_activations_0 = FanoutAWS_io_out_107;
  assign MultiplyAccumulate_107_io_activations_1 = FanoutAWS_1_io_out_107;
  assign MultiplyAccumulate_107_io_activations_2 = FanoutAWS_2_io_out_107;
  assign MultiplyAccumulate_107_io_activations_3 = FanoutAWS_3_io_out_107;
  assign MultiplyAccumulate_107_io_weights = delayWeights_107;
  assign MultiplyAccumulate_108_clock = clock;
  assign MultiplyAccumulate_108_io_activations_0 = FanoutAWS_io_out_108;
  assign MultiplyAccumulate_108_io_activations_1 = FanoutAWS_1_io_out_108;
  assign MultiplyAccumulate_108_io_activations_2 = FanoutAWS_2_io_out_108;
  assign MultiplyAccumulate_108_io_activations_3 = FanoutAWS_3_io_out_108;
  assign MultiplyAccumulate_108_io_weights = delayWeights_108;
  assign MultiplyAccumulate_109_clock = clock;
  assign MultiplyAccumulate_109_io_activations_0 = FanoutAWS_io_out_109;
  assign MultiplyAccumulate_109_io_activations_1 = FanoutAWS_1_io_out_109;
  assign MultiplyAccumulate_109_io_activations_2 = FanoutAWS_2_io_out_109;
  assign MultiplyAccumulate_109_io_activations_3 = FanoutAWS_3_io_out_109;
  assign MultiplyAccumulate_109_io_weights = delayWeights_109;
  assign MultiplyAccumulate_110_clock = clock;
  assign MultiplyAccumulate_110_io_activations_0 = FanoutAWS_io_out_110;
  assign MultiplyAccumulate_110_io_activations_1 = FanoutAWS_1_io_out_110;
  assign MultiplyAccumulate_110_io_activations_2 = FanoutAWS_2_io_out_110;
  assign MultiplyAccumulate_110_io_activations_3 = FanoutAWS_3_io_out_110;
  assign MultiplyAccumulate_110_io_weights = delayWeights_110;
  assign MultiplyAccumulate_111_clock = clock;
  assign MultiplyAccumulate_111_io_activations_0 = FanoutAWS_io_out_111;
  assign MultiplyAccumulate_111_io_activations_1 = FanoutAWS_1_io_out_111;
  assign MultiplyAccumulate_111_io_activations_2 = FanoutAWS_2_io_out_111;
  assign MultiplyAccumulate_111_io_activations_3 = FanoutAWS_3_io_out_111;
  assign MultiplyAccumulate_111_io_weights = delayWeights_111;
  assign MultiplyAccumulate_112_clock = clock;
  assign MultiplyAccumulate_112_io_activations_0 = FanoutAWS_io_out_112;
  assign MultiplyAccumulate_112_io_activations_1 = FanoutAWS_1_io_out_112;
  assign MultiplyAccumulate_112_io_activations_2 = FanoutAWS_2_io_out_112;
  assign MultiplyAccumulate_112_io_activations_3 = FanoutAWS_3_io_out_112;
  assign MultiplyAccumulate_112_io_weights = delayWeights_112;
  assign MultiplyAccumulate_113_clock = clock;
  assign MultiplyAccumulate_113_io_activations_0 = FanoutAWS_io_out_113;
  assign MultiplyAccumulate_113_io_activations_1 = FanoutAWS_1_io_out_113;
  assign MultiplyAccumulate_113_io_activations_2 = FanoutAWS_2_io_out_113;
  assign MultiplyAccumulate_113_io_activations_3 = FanoutAWS_3_io_out_113;
  assign MultiplyAccumulate_113_io_weights = delayWeights_113;
  assign MultiplyAccumulate_114_clock = clock;
  assign MultiplyAccumulate_114_io_activations_0 = FanoutAWS_io_out_114;
  assign MultiplyAccumulate_114_io_activations_1 = FanoutAWS_1_io_out_114;
  assign MultiplyAccumulate_114_io_activations_2 = FanoutAWS_2_io_out_114;
  assign MultiplyAccumulate_114_io_activations_3 = FanoutAWS_3_io_out_114;
  assign MultiplyAccumulate_114_io_weights = delayWeights_114;
  assign MultiplyAccumulate_115_clock = clock;
  assign MultiplyAccumulate_115_io_activations_0 = FanoutAWS_io_out_115;
  assign MultiplyAccumulate_115_io_activations_1 = FanoutAWS_1_io_out_115;
  assign MultiplyAccumulate_115_io_activations_2 = FanoutAWS_2_io_out_115;
  assign MultiplyAccumulate_115_io_activations_3 = FanoutAWS_3_io_out_115;
  assign MultiplyAccumulate_115_io_weights = delayWeights_115;
  assign MultiplyAccumulate_116_clock = clock;
  assign MultiplyAccumulate_116_io_activations_0 = FanoutAWS_io_out_116;
  assign MultiplyAccumulate_116_io_activations_1 = FanoutAWS_1_io_out_116;
  assign MultiplyAccumulate_116_io_activations_2 = FanoutAWS_2_io_out_116;
  assign MultiplyAccumulate_116_io_activations_3 = FanoutAWS_3_io_out_116;
  assign MultiplyAccumulate_116_io_weights = delayWeights_116;
  assign MultiplyAccumulate_117_clock = clock;
  assign MultiplyAccumulate_117_io_activations_0 = FanoutAWS_io_out_117;
  assign MultiplyAccumulate_117_io_activations_1 = FanoutAWS_1_io_out_117;
  assign MultiplyAccumulate_117_io_activations_2 = FanoutAWS_2_io_out_117;
  assign MultiplyAccumulate_117_io_activations_3 = FanoutAWS_3_io_out_117;
  assign MultiplyAccumulate_117_io_weights = delayWeights_117;
  assign MultiplyAccumulate_118_clock = clock;
  assign MultiplyAccumulate_118_io_activations_0 = FanoutAWS_io_out_118;
  assign MultiplyAccumulate_118_io_activations_1 = FanoutAWS_1_io_out_118;
  assign MultiplyAccumulate_118_io_activations_2 = FanoutAWS_2_io_out_118;
  assign MultiplyAccumulate_118_io_activations_3 = FanoutAWS_3_io_out_118;
  assign MultiplyAccumulate_118_io_weights = delayWeights_118;
  assign MultiplyAccumulate_119_clock = clock;
  assign MultiplyAccumulate_119_io_activations_0 = FanoutAWS_io_out_119;
  assign MultiplyAccumulate_119_io_activations_1 = FanoutAWS_1_io_out_119;
  assign MultiplyAccumulate_119_io_activations_2 = FanoutAWS_2_io_out_119;
  assign MultiplyAccumulate_119_io_activations_3 = FanoutAWS_3_io_out_119;
  assign MultiplyAccumulate_119_io_weights = delayWeights_119;
  assign MultiplyAccumulate_120_clock = clock;
  assign MultiplyAccumulate_120_io_activations_0 = FanoutAWS_io_out_120;
  assign MultiplyAccumulate_120_io_activations_1 = FanoutAWS_1_io_out_120;
  assign MultiplyAccumulate_120_io_activations_2 = FanoutAWS_2_io_out_120;
  assign MultiplyAccumulate_120_io_activations_3 = FanoutAWS_3_io_out_120;
  assign MultiplyAccumulate_120_io_weights = delayWeights_120;
  assign MultiplyAccumulate_121_clock = clock;
  assign MultiplyAccumulate_121_io_activations_0 = FanoutAWS_io_out_121;
  assign MultiplyAccumulate_121_io_activations_1 = FanoutAWS_1_io_out_121;
  assign MultiplyAccumulate_121_io_activations_2 = FanoutAWS_2_io_out_121;
  assign MultiplyAccumulate_121_io_activations_3 = FanoutAWS_3_io_out_121;
  assign MultiplyAccumulate_121_io_weights = delayWeights_121;
  assign MultiplyAccumulate_122_clock = clock;
  assign MultiplyAccumulate_122_io_activations_0 = FanoutAWS_io_out_122;
  assign MultiplyAccumulate_122_io_activations_1 = FanoutAWS_1_io_out_122;
  assign MultiplyAccumulate_122_io_activations_2 = FanoutAWS_2_io_out_122;
  assign MultiplyAccumulate_122_io_activations_3 = FanoutAWS_3_io_out_122;
  assign MultiplyAccumulate_122_io_weights = delayWeights_122;
  assign MultiplyAccumulate_123_clock = clock;
  assign MultiplyAccumulate_123_io_activations_0 = FanoutAWS_io_out_123;
  assign MultiplyAccumulate_123_io_activations_1 = FanoutAWS_1_io_out_123;
  assign MultiplyAccumulate_123_io_activations_2 = FanoutAWS_2_io_out_123;
  assign MultiplyAccumulate_123_io_activations_3 = FanoutAWS_3_io_out_123;
  assign MultiplyAccumulate_123_io_weights = delayWeights_123;
  assign MultiplyAccumulate_124_clock = clock;
  assign MultiplyAccumulate_124_io_activations_0 = FanoutAWS_io_out_124;
  assign MultiplyAccumulate_124_io_activations_1 = FanoutAWS_1_io_out_124;
  assign MultiplyAccumulate_124_io_activations_2 = FanoutAWS_2_io_out_124;
  assign MultiplyAccumulate_124_io_activations_3 = FanoutAWS_3_io_out_124;
  assign MultiplyAccumulate_124_io_weights = delayWeights_124;
  assign MultiplyAccumulate_125_clock = clock;
  assign MultiplyAccumulate_125_io_activations_0 = FanoutAWS_io_out_125;
  assign MultiplyAccumulate_125_io_activations_1 = FanoutAWS_1_io_out_125;
  assign MultiplyAccumulate_125_io_activations_2 = FanoutAWS_2_io_out_125;
  assign MultiplyAccumulate_125_io_activations_3 = FanoutAWS_3_io_out_125;
  assign MultiplyAccumulate_125_io_weights = delayWeights_125;
  assign MultiplyAccumulate_126_clock = clock;
  assign MultiplyAccumulate_126_io_activations_0 = FanoutAWS_io_out_126;
  assign MultiplyAccumulate_126_io_activations_1 = FanoutAWS_1_io_out_126;
  assign MultiplyAccumulate_126_io_activations_2 = FanoutAWS_2_io_out_126;
  assign MultiplyAccumulate_126_io_activations_3 = FanoutAWS_3_io_out_126;
  assign MultiplyAccumulate_126_io_weights = delayWeights_126;
  assign MultiplyAccumulate_127_clock = clock;
  assign MultiplyAccumulate_127_io_activations_0 = FanoutAWS_io_out_127;
  assign MultiplyAccumulate_127_io_activations_1 = FanoutAWS_1_io_out_127;
  assign MultiplyAccumulate_127_io_activations_2 = FanoutAWS_2_io_out_127;
  assign MultiplyAccumulate_127_io_activations_3 = FanoutAWS_3_io_out_127;
  assign MultiplyAccumulate_127_io_weights = delayWeights_127;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  cntr = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_293 = _RAND_1[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  currActs_0 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  currActs_1 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  currActs_2 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  currActs_3 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  _T_711_0 = _RAND_6[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  _T_711_1 = _RAND_7[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  _T_711_2 = _RAND_8[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  _T_711_3 = _RAND_9[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  _T_711_4 = _RAND_10[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  _T_711_5 = _RAND_11[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  _T_711_6 = _RAND_12[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  _T_711_7 = _RAND_13[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  _T_711_8 = _RAND_14[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  _T_711_9 = _RAND_15[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  _T_711_10 = _RAND_16[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  _T_711_11 = _RAND_17[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  _T_711_12 = _RAND_18[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  _T_711_13 = _RAND_19[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  _T_711_14 = _RAND_20[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  _T_711_15 = _RAND_21[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  _T_711_16 = _RAND_22[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  _T_711_17 = _RAND_23[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  _T_711_18 = _RAND_24[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  _T_711_19 = _RAND_25[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  _T_711_20 = _RAND_26[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  _T_711_21 = _RAND_27[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  _T_711_22 = _RAND_28[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  _T_711_23 = _RAND_29[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  _T_711_24 = _RAND_30[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  _T_711_25 = _RAND_31[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  _T_711_26 = _RAND_32[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{$random}};
  _T_711_27 = _RAND_33[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{$random}};
  _T_711_28 = _RAND_34[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{$random}};
  _T_711_29 = _RAND_35[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{$random}};
  _T_711_30 = _RAND_36[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{$random}};
  _T_711_31 = _RAND_37[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{$random}};
  _T_711_32 = _RAND_38[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{$random}};
  _T_711_33 = _RAND_39[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{$random}};
  _T_711_34 = _RAND_40[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{$random}};
  _T_711_35 = _RAND_41[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{$random}};
  _T_711_36 = _RAND_42[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{$random}};
  _T_711_37 = _RAND_43[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{$random}};
  _T_711_38 = _RAND_44[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{$random}};
  _T_711_39 = _RAND_45[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{$random}};
  _T_711_40 = _RAND_46[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{$random}};
  _T_711_41 = _RAND_47[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{$random}};
  _T_711_42 = _RAND_48[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{$random}};
  _T_711_43 = _RAND_49[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{$random}};
  _T_711_44 = _RAND_50[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{$random}};
  _T_711_45 = _RAND_51[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{$random}};
  _T_711_46 = _RAND_52[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{$random}};
  _T_711_47 = _RAND_53[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{$random}};
  _T_711_48 = _RAND_54[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{$random}};
  _T_711_49 = _RAND_55[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{$random}};
  _T_711_50 = _RAND_56[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{$random}};
  _T_711_51 = _RAND_57[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{$random}};
  _T_711_52 = _RAND_58[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{$random}};
  _T_711_53 = _RAND_59[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{$random}};
  _T_711_54 = _RAND_60[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{$random}};
  _T_711_55 = _RAND_61[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{$random}};
  _T_711_56 = _RAND_62[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{$random}};
  _T_711_57 = _RAND_63[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{$random}};
  _T_711_58 = _RAND_64[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{$random}};
  _T_711_59 = _RAND_65[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{$random}};
  _T_711_60 = _RAND_66[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{$random}};
  _T_711_61 = _RAND_67[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{$random}};
  _T_711_62 = _RAND_68[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{$random}};
  _T_711_63 = _RAND_69[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{$random}};
  _T_711_64 = _RAND_70[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{$random}};
  _T_711_65 = _RAND_71[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{$random}};
  _T_711_66 = _RAND_72[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{$random}};
  _T_711_67 = _RAND_73[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{$random}};
  _T_711_68 = _RAND_74[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{$random}};
  _T_711_69 = _RAND_75[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{$random}};
  _T_711_70 = _RAND_76[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{$random}};
  _T_711_71 = _RAND_77[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{$random}};
  _T_711_72 = _RAND_78[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{$random}};
  _T_711_73 = _RAND_79[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{$random}};
  _T_711_74 = _RAND_80[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{$random}};
  _T_711_75 = _RAND_81[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{$random}};
  _T_711_76 = _RAND_82[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{$random}};
  _T_711_77 = _RAND_83[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{$random}};
  _T_711_78 = _RAND_84[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{$random}};
  _T_711_79 = _RAND_85[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{$random}};
  _T_711_80 = _RAND_86[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{$random}};
  _T_711_81 = _RAND_87[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{$random}};
  _T_711_82 = _RAND_88[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{$random}};
  _T_711_83 = _RAND_89[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{$random}};
  _T_711_84 = _RAND_90[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{$random}};
  _T_711_85 = _RAND_91[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{$random}};
  _T_711_86 = _RAND_92[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{$random}};
  _T_711_87 = _RAND_93[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{$random}};
  _T_711_88 = _RAND_94[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{$random}};
  _T_711_89 = _RAND_95[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{$random}};
  _T_711_90 = _RAND_96[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{$random}};
  _T_711_91 = _RAND_97[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{$random}};
  _T_711_92 = _RAND_98[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{$random}};
  _T_711_93 = _RAND_99[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{$random}};
  _T_711_94 = _RAND_100[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{$random}};
  _T_711_95 = _RAND_101[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{$random}};
  _T_711_96 = _RAND_102[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{$random}};
  _T_711_97 = _RAND_103[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{$random}};
  _T_711_98 = _RAND_104[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{$random}};
  _T_711_99 = _RAND_105[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{$random}};
  _T_711_100 = _RAND_106[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{$random}};
  _T_711_101 = _RAND_107[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{$random}};
  _T_711_102 = _RAND_108[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{$random}};
  _T_711_103 = _RAND_109[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{$random}};
  _T_711_104 = _RAND_110[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{$random}};
  _T_711_105 = _RAND_111[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{$random}};
  _T_711_106 = _RAND_112[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{$random}};
  _T_711_107 = _RAND_113[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{$random}};
  _T_711_108 = _RAND_114[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{$random}};
  _T_711_109 = _RAND_115[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{$random}};
  _T_711_110 = _RAND_116[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{$random}};
  _T_711_111 = _RAND_117[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{$random}};
  _T_711_112 = _RAND_118[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{$random}};
  _T_711_113 = _RAND_119[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{$random}};
  _T_711_114 = _RAND_120[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{$random}};
  _T_711_115 = _RAND_121[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{$random}};
  _T_711_116 = _RAND_122[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{$random}};
  _T_711_117 = _RAND_123[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{$random}};
  _T_711_118 = _RAND_124[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{$random}};
  _T_711_119 = _RAND_125[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{$random}};
  _T_711_120 = _RAND_126[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{$random}};
  _T_711_121 = _RAND_127[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{$random}};
  _T_711_122 = _RAND_128[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{$random}};
  _T_711_123 = _RAND_129[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{$random}};
  _T_711_124 = _RAND_130[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{$random}};
  _T_711_125 = _RAND_131[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{$random}};
  _T_711_126 = _RAND_132[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{$random}};
  _T_711_127 = _RAND_133[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{$random}};
  delayWeights_0 = _RAND_134[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{$random}};
  delayWeights_1 = _RAND_135[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{$random}};
  delayWeights_2 = _RAND_136[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{$random}};
  delayWeights_3 = _RAND_137[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{$random}};
  delayWeights_4 = _RAND_138[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{$random}};
  delayWeights_5 = _RAND_139[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{$random}};
  delayWeights_6 = _RAND_140[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{$random}};
  delayWeights_7 = _RAND_141[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{$random}};
  delayWeights_8 = _RAND_142[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{$random}};
  delayWeights_9 = _RAND_143[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{$random}};
  delayWeights_10 = _RAND_144[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{$random}};
  delayWeights_11 = _RAND_145[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{$random}};
  delayWeights_12 = _RAND_146[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{$random}};
  delayWeights_13 = _RAND_147[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{$random}};
  delayWeights_14 = _RAND_148[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{$random}};
  delayWeights_15 = _RAND_149[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{$random}};
  delayWeights_16 = _RAND_150[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{$random}};
  delayWeights_17 = _RAND_151[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{$random}};
  delayWeights_18 = _RAND_152[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{$random}};
  delayWeights_19 = _RAND_153[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{$random}};
  delayWeights_20 = _RAND_154[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{$random}};
  delayWeights_21 = _RAND_155[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{$random}};
  delayWeights_22 = _RAND_156[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{$random}};
  delayWeights_23 = _RAND_157[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{$random}};
  delayWeights_24 = _RAND_158[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{$random}};
  delayWeights_25 = _RAND_159[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{$random}};
  delayWeights_26 = _RAND_160[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{$random}};
  delayWeights_27 = _RAND_161[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{$random}};
  delayWeights_28 = _RAND_162[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{$random}};
  delayWeights_29 = _RAND_163[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{$random}};
  delayWeights_30 = _RAND_164[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{$random}};
  delayWeights_31 = _RAND_165[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{$random}};
  delayWeights_32 = _RAND_166[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{$random}};
  delayWeights_33 = _RAND_167[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{$random}};
  delayWeights_34 = _RAND_168[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{$random}};
  delayWeights_35 = _RAND_169[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{$random}};
  delayWeights_36 = _RAND_170[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{$random}};
  delayWeights_37 = _RAND_171[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{$random}};
  delayWeights_38 = _RAND_172[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{$random}};
  delayWeights_39 = _RAND_173[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{$random}};
  delayWeights_40 = _RAND_174[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{$random}};
  delayWeights_41 = _RAND_175[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{$random}};
  delayWeights_42 = _RAND_176[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{$random}};
  delayWeights_43 = _RAND_177[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{$random}};
  delayWeights_44 = _RAND_178[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{$random}};
  delayWeights_45 = _RAND_179[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{$random}};
  delayWeights_46 = _RAND_180[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{$random}};
  delayWeights_47 = _RAND_181[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{$random}};
  delayWeights_48 = _RAND_182[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{$random}};
  delayWeights_49 = _RAND_183[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{$random}};
  delayWeights_50 = _RAND_184[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{$random}};
  delayWeights_51 = _RAND_185[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{$random}};
  delayWeights_52 = _RAND_186[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{$random}};
  delayWeights_53 = _RAND_187[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{$random}};
  delayWeights_54 = _RAND_188[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{$random}};
  delayWeights_55 = _RAND_189[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{$random}};
  delayWeights_56 = _RAND_190[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{$random}};
  delayWeights_57 = _RAND_191[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{$random}};
  delayWeights_58 = _RAND_192[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{$random}};
  delayWeights_59 = _RAND_193[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{$random}};
  delayWeights_60 = _RAND_194[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{$random}};
  delayWeights_61 = _RAND_195[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{$random}};
  delayWeights_62 = _RAND_196[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{$random}};
  delayWeights_63 = _RAND_197[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{$random}};
  delayWeights_64 = _RAND_198[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{$random}};
  delayWeights_65 = _RAND_199[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{$random}};
  delayWeights_66 = _RAND_200[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{$random}};
  delayWeights_67 = _RAND_201[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{$random}};
  delayWeights_68 = _RAND_202[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{$random}};
  delayWeights_69 = _RAND_203[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{$random}};
  delayWeights_70 = _RAND_204[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{$random}};
  delayWeights_71 = _RAND_205[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{$random}};
  delayWeights_72 = _RAND_206[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{$random}};
  delayWeights_73 = _RAND_207[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{$random}};
  delayWeights_74 = _RAND_208[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{$random}};
  delayWeights_75 = _RAND_209[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{$random}};
  delayWeights_76 = _RAND_210[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{$random}};
  delayWeights_77 = _RAND_211[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{$random}};
  delayWeights_78 = _RAND_212[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{$random}};
  delayWeights_79 = _RAND_213[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{$random}};
  delayWeights_80 = _RAND_214[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{$random}};
  delayWeights_81 = _RAND_215[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{$random}};
  delayWeights_82 = _RAND_216[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{$random}};
  delayWeights_83 = _RAND_217[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{$random}};
  delayWeights_84 = _RAND_218[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{$random}};
  delayWeights_85 = _RAND_219[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{$random}};
  delayWeights_86 = _RAND_220[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{$random}};
  delayWeights_87 = _RAND_221[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{$random}};
  delayWeights_88 = _RAND_222[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{$random}};
  delayWeights_89 = _RAND_223[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{$random}};
  delayWeights_90 = _RAND_224[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{$random}};
  delayWeights_91 = _RAND_225[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{$random}};
  delayWeights_92 = _RAND_226[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{$random}};
  delayWeights_93 = _RAND_227[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{$random}};
  delayWeights_94 = _RAND_228[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{$random}};
  delayWeights_95 = _RAND_229[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{$random}};
  delayWeights_96 = _RAND_230[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{$random}};
  delayWeights_97 = _RAND_231[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{$random}};
  delayWeights_98 = _RAND_232[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{$random}};
  delayWeights_99 = _RAND_233[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{$random}};
  delayWeights_100 = _RAND_234[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{$random}};
  delayWeights_101 = _RAND_235[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{$random}};
  delayWeights_102 = _RAND_236[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{$random}};
  delayWeights_103 = _RAND_237[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{$random}};
  delayWeights_104 = _RAND_238[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{$random}};
  delayWeights_105 = _RAND_239[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{$random}};
  delayWeights_106 = _RAND_240[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{$random}};
  delayWeights_107 = _RAND_241[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{$random}};
  delayWeights_108 = _RAND_242[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{$random}};
  delayWeights_109 = _RAND_243[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{$random}};
  delayWeights_110 = _RAND_244[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{$random}};
  delayWeights_111 = _RAND_245[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{$random}};
  delayWeights_112 = _RAND_246[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{$random}};
  delayWeights_113 = _RAND_247[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{$random}};
  delayWeights_114 = _RAND_248[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{$random}};
  delayWeights_115 = _RAND_249[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{$random}};
  delayWeights_116 = _RAND_250[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{$random}};
  delayWeights_117 = _RAND_251[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{$random}};
  delayWeights_118 = _RAND_252[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{$random}};
  delayWeights_119 = _RAND_253[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{$random}};
  delayWeights_120 = _RAND_254[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{$random}};
  delayWeights_121 = _RAND_255[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{$random}};
  delayWeights_122 = _RAND_256[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{$random}};
  delayWeights_123 = _RAND_257[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{$random}};
  delayWeights_124 = _RAND_258[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{$random}};
  delayWeights_125 = _RAND_259[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{$random}};
  delayWeights_126 = _RAND_260[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{$random}};
  delayWeights_127 = _RAND_261[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{$random}};
  cummulativeSums_0 = _RAND_262[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{$random}};
  cummulativeSums_1 = _RAND_263[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{$random}};
  cummulativeSums_2 = _RAND_264[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{$random}};
  cummulativeSums_3 = _RAND_265[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{$random}};
  cummulativeSums_4 = _RAND_266[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{$random}};
  cummulativeSums_5 = _RAND_267[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{$random}};
  cummulativeSums_6 = _RAND_268[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{$random}};
  cummulativeSums_7 = _RAND_269[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{$random}};
  cummulativeSums_8 = _RAND_270[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{$random}};
  cummulativeSums_9 = _RAND_271[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{$random}};
  cummulativeSums_10 = _RAND_272[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{$random}};
  cummulativeSums_11 = _RAND_273[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{$random}};
  cummulativeSums_12 = _RAND_274[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{$random}};
  cummulativeSums_13 = _RAND_275[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{$random}};
  cummulativeSums_14 = _RAND_276[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{$random}};
  cummulativeSums_15 = _RAND_277[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{$random}};
  cummulativeSums_16 = _RAND_278[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{$random}};
  cummulativeSums_17 = _RAND_279[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{$random}};
  cummulativeSums_18 = _RAND_280[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{$random}};
  cummulativeSums_19 = _RAND_281[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{$random}};
  cummulativeSums_20 = _RAND_282[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{$random}};
  cummulativeSums_21 = _RAND_283[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{$random}};
  cummulativeSums_22 = _RAND_284[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{$random}};
  cummulativeSums_23 = _RAND_285[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{$random}};
  cummulativeSums_24 = _RAND_286[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{$random}};
  cummulativeSums_25 = _RAND_287[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{$random}};
  cummulativeSums_26 = _RAND_288[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{$random}};
  cummulativeSums_27 = _RAND_289[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{$random}};
  cummulativeSums_28 = _RAND_290[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{$random}};
  cummulativeSums_29 = _RAND_291[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{$random}};
  cummulativeSums_30 = _RAND_292[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{$random}};
  cummulativeSums_31 = _RAND_293[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{$random}};
  cummulativeSums_32 = _RAND_294[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{$random}};
  cummulativeSums_33 = _RAND_295[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{$random}};
  cummulativeSums_34 = _RAND_296[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{$random}};
  cummulativeSums_35 = _RAND_297[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{$random}};
  cummulativeSums_36 = _RAND_298[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{$random}};
  cummulativeSums_37 = _RAND_299[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{$random}};
  cummulativeSums_38 = _RAND_300[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{$random}};
  cummulativeSums_39 = _RAND_301[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{$random}};
  cummulativeSums_40 = _RAND_302[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{$random}};
  cummulativeSums_41 = _RAND_303[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{$random}};
  cummulativeSums_42 = _RAND_304[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{$random}};
  cummulativeSums_43 = _RAND_305[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{$random}};
  cummulativeSums_44 = _RAND_306[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{$random}};
  cummulativeSums_45 = _RAND_307[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{$random}};
  cummulativeSums_46 = _RAND_308[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{$random}};
  cummulativeSums_47 = _RAND_309[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{$random}};
  cummulativeSums_48 = _RAND_310[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{$random}};
  cummulativeSums_49 = _RAND_311[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{$random}};
  cummulativeSums_50 = _RAND_312[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{$random}};
  cummulativeSums_51 = _RAND_313[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{$random}};
  cummulativeSums_52 = _RAND_314[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{$random}};
  cummulativeSums_53 = _RAND_315[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{$random}};
  cummulativeSums_54 = _RAND_316[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{$random}};
  cummulativeSums_55 = _RAND_317[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{$random}};
  cummulativeSums_56 = _RAND_318[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{$random}};
  cummulativeSums_57 = _RAND_319[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{$random}};
  cummulativeSums_58 = _RAND_320[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{$random}};
  cummulativeSums_59 = _RAND_321[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{$random}};
  cummulativeSums_60 = _RAND_322[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{$random}};
  cummulativeSums_61 = _RAND_323[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{$random}};
  cummulativeSums_62 = _RAND_324[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{$random}};
  cummulativeSums_63 = _RAND_325[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{$random}};
  cummulativeSums_64 = _RAND_326[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{$random}};
  cummulativeSums_65 = _RAND_327[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{$random}};
  cummulativeSums_66 = _RAND_328[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{$random}};
  cummulativeSums_67 = _RAND_329[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{$random}};
  cummulativeSums_68 = _RAND_330[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{$random}};
  cummulativeSums_69 = _RAND_331[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{$random}};
  cummulativeSums_70 = _RAND_332[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{$random}};
  cummulativeSums_71 = _RAND_333[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{$random}};
  cummulativeSums_72 = _RAND_334[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{$random}};
  cummulativeSums_73 = _RAND_335[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{$random}};
  cummulativeSums_74 = _RAND_336[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{$random}};
  cummulativeSums_75 = _RAND_337[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{$random}};
  cummulativeSums_76 = _RAND_338[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{$random}};
  cummulativeSums_77 = _RAND_339[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{$random}};
  cummulativeSums_78 = _RAND_340[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{$random}};
  cummulativeSums_79 = _RAND_341[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{$random}};
  cummulativeSums_80 = _RAND_342[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{$random}};
  cummulativeSums_81 = _RAND_343[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{$random}};
  cummulativeSums_82 = _RAND_344[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{$random}};
  cummulativeSums_83 = _RAND_345[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{$random}};
  cummulativeSums_84 = _RAND_346[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{$random}};
  cummulativeSums_85 = _RAND_347[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{$random}};
  cummulativeSums_86 = _RAND_348[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{$random}};
  cummulativeSums_87 = _RAND_349[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{$random}};
  cummulativeSums_88 = _RAND_350[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{$random}};
  cummulativeSums_89 = _RAND_351[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{$random}};
  cummulativeSums_90 = _RAND_352[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{$random}};
  cummulativeSums_91 = _RAND_353[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{$random}};
  cummulativeSums_92 = _RAND_354[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{$random}};
  cummulativeSums_93 = _RAND_355[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{$random}};
  cummulativeSums_94 = _RAND_356[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{$random}};
  cummulativeSums_95 = _RAND_357[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{$random}};
  cummulativeSums_96 = _RAND_358[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{$random}};
  cummulativeSums_97 = _RAND_359[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{$random}};
  cummulativeSums_98 = _RAND_360[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{$random}};
  cummulativeSums_99 = _RAND_361[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{$random}};
  cummulativeSums_100 = _RAND_362[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{$random}};
  cummulativeSums_101 = _RAND_363[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{$random}};
  cummulativeSums_102 = _RAND_364[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{$random}};
  cummulativeSums_103 = _RAND_365[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{$random}};
  cummulativeSums_104 = _RAND_366[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{$random}};
  cummulativeSums_105 = _RAND_367[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{$random}};
  cummulativeSums_106 = _RAND_368[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{$random}};
  cummulativeSums_107 = _RAND_369[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{$random}};
  cummulativeSums_108 = _RAND_370[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{$random}};
  cummulativeSums_109 = _RAND_371[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{$random}};
  cummulativeSums_110 = _RAND_372[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{$random}};
  cummulativeSums_111 = _RAND_373[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{$random}};
  cummulativeSums_112 = _RAND_374[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{$random}};
  cummulativeSums_113 = _RAND_375[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{$random}};
  cummulativeSums_114 = _RAND_376[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{$random}};
  cummulativeSums_115 = _RAND_377[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{$random}};
  cummulativeSums_116 = _RAND_378[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{$random}};
  cummulativeSums_117 = _RAND_379[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{$random}};
  cummulativeSums_118 = _RAND_380[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{$random}};
  cummulativeSums_119 = _RAND_381[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{$random}};
  cummulativeSums_120 = _RAND_382[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{$random}};
  cummulativeSums_121 = _RAND_383[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{$random}};
  cummulativeSums_122 = _RAND_384[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{$random}};
  cummulativeSums_123 = _RAND_385[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{$random}};
  cummulativeSums_124 = _RAND_386[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{$random}};
  cummulativeSums_125 = _RAND_387[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{$random}};
  cummulativeSums_126 = _RAND_388[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{$random}};
  cummulativeSums_127 = _RAND_389[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{$random}};
  _T_2401 = _RAND_390[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{$random}};
  _T_2403 = _RAND_391[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{$random}};
  _T_2405 = _RAND_392[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{$random}};
  _T_2407 = _RAND_393[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{$random}};
  _T_2409 = _RAND_394[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{$random}};
  _T_2411 = _RAND_395[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{$random}};
  rst = _RAND_396[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{$random}};
  done = _RAND_397[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{$random}};
  _T_2422 = _RAND_398[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{$random}};
  _T_2424 = _RAND_399[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{$random}};
  _T_2426 = _RAND_400[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{$random}};
  _T_2428 = _RAND_401[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{$random}};
  _T_2430 = _RAND_402[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{$random}};
  _T_2432 = _RAND_403[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{$random}};
  vld = _RAND_404[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cntr <= 10'h0;
    end else begin
      if (io_dataIn_valid) begin
        cntr <= _T_159;
      end
    end
    _T_293 <= cntr;
    currActs_0 <= io_dataIn_bits_0;
    currActs_1 <= io_dataIn_bits_1;
    currActs_2 <= io_dataIn_bits_2;
    currActs_3 <= io_dataIn_bits_3;
    _T_711_0 <= currWeights_0;
    _T_711_1 <= currWeights_1;
    _T_711_2 <= currWeights_2;
    _T_711_3 <= currWeights_3;
    _T_711_4 <= currWeights_4;
    _T_711_5 <= currWeights_5;
    _T_711_6 <= currWeights_6;
    _T_711_7 <= currWeights_7;
    _T_711_8 <= currWeights_8;
    _T_711_9 <= currWeights_9;
    _T_711_10 <= currWeights_10;
    _T_711_11 <= currWeights_11;
    _T_711_12 <= currWeights_12;
    _T_711_13 <= currWeights_13;
    _T_711_14 <= currWeights_14;
    _T_711_15 <= currWeights_15;
    _T_711_16 <= currWeights_16;
    _T_711_17 <= currWeights_17;
    _T_711_18 <= currWeights_18;
    _T_711_19 <= currWeights_19;
    _T_711_20 <= currWeights_20;
    _T_711_21 <= currWeights_21;
    _T_711_22 <= currWeights_22;
    _T_711_23 <= currWeights_23;
    _T_711_24 <= currWeights_24;
    _T_711_25 <= currWeights_25;
    _T_711_26 <= currWeights_26;
    _T_711_27 <= currWeights_27;
    _T_711_28 <= currWeights_28;
    _T_711_29 <= currWeights_29;
    _T_711_30 <= currWeights_30;
    _T_711_31 <= currWeights_31;
    _T_711_32 <= currWeights_32;
    _T_711_33 <= currWeights_33;
    _T_711_34 <= currWeights_34;
    _T_711_35 <= currWeights_35;
    _T_711_36 <= currWeights_36;
    _T_711_37 <= currWeights_37;
    _T_711_38 <= currWeights_38;
    _T_711_39 <= currWeights_39;
    _T_711_40 <= currWeights_40;
    _T_711_41 <= currWeights_41;
    _T_711_42 <= currWeights_42;
    _T_711_43 <= currWeights_43;
    _T_711_44 <= currWeights_44;
    _T_711_45 <= currWeights_45;
    _T_711_46 <= currWeights_46;
    _T_711_47 <= currWeights_47;
    _T_711_48 <= currWeights_48;
    _T_711_49 <= currWeights_49;
    _T_711_50 <= currWeights_50;
    _T_711_51 <= currWeights_51;
    _T_711_52 <= currWeights_52;
    _T_711_53 <= currWeights_53;
    _T_711_54 <= currWeights_54;
    _T_711_55 <= currWeights_55;
    _T_711_56 <= currWeights_56;
    _T_711_57 <= currWeights_57;
    _T_711_58 <= currWeights_58;
    _T_711_59 <= currWeights_59;
    _T_711_60 <= currWeights_60;
    _T_711_61 <= currWeights_61;
    _T_711_62 <= currWeights_62;
    _T_711_63 <= currWeights_63;
    _T_711_64 <= currWeights_64;
    _T_711_65 <= currWeights_65;
    _T_711_66 <= currWeights_66;
    _T_711_67 <= currWeights_67;
    _T_711_68 <= currWeights_68;
    _T_711_69 <= currWeights_69;
    _T_711_70 <= currWeights_70;
    _T_711_71 <= currWeights_71;
    _T_711_72 <= currWeights_72;
    _T_711_73 <= currWeights_73;
    _T_711_74 <= currWeights_74;
    _T_711_75 <= currWeights_75;
    _T_711_76 <= currWeights_76;
    _T_711_77 <= currWeights_77;
    _T_711_78 <= currWeights_78;
    _T_711_79 <= currWeights_79;
    _T_711_80 <= currWeights_80;
    _T_711_81 <= currWeights_81;
    _T_711_82 <= currWeights_82;
    _T_711_83 <= currWeights_83;
    _T_711_84 <= currWeights_84;
    _T_711_85 <= currWeights_85;
    _T_711_86 <= currWeights_86;
    _T_711_87 <= currWeights_87;
    _T_711_88 <= currWeights_88;
    _T_711_89 <= currWeights_89;
    _T_711_90 <= currWeights_90;
    _T_711_91 <= currWeights_91;
    _T_711_92 <= currWeights_92;
    _T_711_93 <= currWeights_93;
    _T_711_94 <= currWeights_94;
    _T_711_95 <= currWeights_95;
    _T_711_96 <= currWeights_96;
    _T_711_97 <= currWeights_97;
    _T_711_98 <= currWeights_98;
    _T_711_99 <= currWeights_99;
    _T_711_100 <= currWeights_100;
    _T_711_101 <= currWeights_101;
    _T_711_102 <= currWeights_102;
    _T_711_103 <= currWeights_103;
    _T_711_104 <= currWeights_104;
    _T_711_105 <= currWeights_105;
    _T_711_106 <= currWeights_106;
    _T_711_107 <= currWeights_107;
    _T_711_108 <= currWeights_108;
    _T_711_109 <= currWeights_109;
    _T_711_110 <= currWeights_110;
    _T_711_111 <= currWeights_111;
    _T_711_112 <= currWeights_112;
    _T_711_113 <= currWeights_113;
    _T_711_114 <= currWeights_114;
    _T_711_115 <= currWeights_115;
    _T_711_116 <= currWeights_116;
    _T_711_117 <= currWeights_117;
    _T_711_118 <= currWeights_118;
    _T_711_119 <= currWeights_119;
    _T_711_120 <= currWeights_120;
    _T_711_121 <= currWeights_121;
    _T_711_122 <= currWeights_122;
    _T_711_123 <= currWeights_123;
    _T_711_124 <= currWeights_124;
    _T_711_125 <= currWeights_125;
    _T_711_126 <= currWeights_126;
    _T_711_127 <= currWeights_127;
    delayWeights_0 <= _T_711_0;
    delayWeights_1 <= _T_711_1;
    delayWeights_2 <= _T_711_2;
    delayWeights_3 <= _T_711_3;
    delayWeights_4 <= _T_711_4;
    delayWeights_5 <= _T_711_5;
    delayWeights_6 <= _T_711_6;
    delayWeights_7 <= _T_711_7;
    delayWeights_8 <= _T_711_8;
    delayWeights_9 <= _T_711_9;
    delayWeights_10 <= _T_711_10;
    delayWeights_11 <= _T_711_11;
    delayWeights_12 <= _T_711_12;
    delayWeights_13 <= _T_711_13;
    delayWeights_14 <= _T_711_14;
    delayWeights_15 <= _T_711_15;
    delayWeights_16 <= _T_711_16;
    delayWeights_17 <= _T_711_17;
    delayWeights_18 <= _T_711_18;
    delayWeights_19 <= _T_711_19;
    delayWeights_20 <= _T_711_20;
    delayWeights_21 <= _T_711_21;
    delayWeights_22 <= _T_711_22;
    delayWeights_23 <= _T_711_23;
    delayWeights_24 <= _T_711_24;
    delayWeights_25 <= _T_711_25;
    delayWeights_26 <= _T_711_26;
    delayWeights_27 <= _T_711_27;
    delayWeights_28 <= _T_711_28;
    delayWeights_29 <= _T_711_29;
    delayWeights_30 <= _T_711_30;
    delayWeights_31 <= _T_711_31;
    delayWeights_32 <= _T_711_32;
    delayWeights_33 <= _T_711_33;
    delayWeights_34 <= _T_711_34;
    delayWeights_35 <= _T_711_35;
    delayWeights_36 <= _T_711_36;
    delayWeights_37 <= _T_711_37;
    delayWeights_38 <= _T_711_38;
    delayWeights_39 <= _T_711_39;
    delayWeights_40 <= _T_711_40;
    delayWeights_41 <= _T_711_41;
    delayWeights_42 <= _T_711_42;
    delayWeights_43 <= _T_711_43;
    delayWeights_44 <= _T_711_44;
    delayWeights_45 <= _T_711_45;
    delayWeights_46 <= _T_711_46;
    delayWeights_47 <= _T_711_47;
    delayWeights_48 <= _T_711_48;
    delayWeights_49 <= _T_711_49;
    delayWeights_50 <= _T_711_50;
    delayWeights_51 <= _T_711_51;
    delayWeights_52 <= _T_711_52;
    delayWeights_53 <= _T_711_53;
    delayWeights_54 <= _T_711_54;
    delayWeights_55 <= _T_711_55;
    delayWeights_56 <= _T_711_56;
    delayWeights_57 <= _T_711_57;
    delayWeights_58 <= _T_711_58;
    delayWeights_59 <= _T_711_59;
    delayWeights_60 <= _T_711_60;
    delayWeights_61 <= _T_711_61;
    delayWeights_62 <= _T_711_62;
    delayWeights_63 <= _T_711_63;
    delayWeights_64 <= _T_711_64;
    delayWeights_65 <= _T_711_65;
    delayWeights_66 <= _T_711_66;
    delayWeights_67 <= _T_711_67;
    delayWeights_68 <= _T_711_68;
    delayWeights_69 <= _T_711_69;
    delayWeights_70 <= _T_711_70;
    delayWeights_71 <= _T_711_71;
    delayWeights_72 <= _T_711_72;
    delayWeights_73 <= _T_711_73;
    delayWeights_74 <= _T_711_74;
    delayWeights_75 <= _T_711_75;
    delayWeights_76 <= _T_711_76;
    delayWeights_77 <= _T_711_77;
    delayWeights_78 <= _T_711_78;
    delayWeights_79 <= _T_711_79;
    delayWeights_80 <= _T_711_80;
    delayWeights_81 <= _T_711_81;
    delayWeights_82 <= _T_711_82;
    delayWeights_83 <= _T_711_83;
    delayWeights_84 <= _T_711_84;
    delayWeights_85 <= _T_711_85;
    delayWeights_86 <= _T_711_86;
    delayWeights_87 <= _T_711_87;
    delayWeights_88 <= _T_711_88;
    delayWeights_89 <= _T_711_89;
    delayWeights_90 <= _T_711_90;
    delayWeights_91 <= _T_711_91;
    delayWeights_92 <= _T_711_92;
    delayWeights_93 <= _T_711_93;
    delayWeights_94 <= _T_711_94;
    delayWeights_95 <= _T_711_95;
    delayWeights_96 <= _T_711_96;
    delayWeights_97 <= _T_711_97;
    delayWeights_98 <= _T_711_98;
    delayWeights_99 <= _T_711_99;
    delayWeights_100 <= _T_711_100;
    delayWeights_101 <= _T_711_101;
    delayWeights_102 <= _T_711_102;
    delayWeights_103 <= _T_711_103;
    delayWeights_104 <= _T_711_104;
    delayWeights_105 <= _T_711_105;
    delayWeights_106 <= _T_711_106;
    delayWeights_107 <= _T_711_107;
    delayWeights_108 <= _T_711_108;
    delayWeights_109 <= _T_711_109;
    delayWeights_110 <= _T_711_110;
    delayWeights_111 <= _T_711_111;
    delayWeights_112 <= _T_711_112;
    delayWeights_113 <= _T_711_113;
    delayWeights_114 <= _T_711_114;
    delayWeights_115 <= _T_711_115;
    delayWeights_116 <= _T_711_116;
    delayWeights_117 <= _T_711_117;
    delayWeights_118 <= _T_711_118;
    delayWeights_119 <= _T_711_119;
    delayWeights_120 <= _T_711_120;
    delayWeights_121 <= _T_711_121;
    delayWeights_122 <= _T_711_122;
    delayWeights_123 <= _T_711_123;
    delayWeights_124 <= _T_711_124;
    delayWeights_125 <= _T_711_125;
    delayWeights_126 <= _T_711_126;
    delayWeights_127 <= _T_711_127;
    if (_T_2438) begin
      cummulativeSums_0 <= MultiplyAccumulate_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_0 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_0 <= _T_2436;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_1 <= MultiplyAccumulate_1_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_1 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_1 <= _T_2441;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_2 <= MultiplyAccumulate_2_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_2 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_2 <= _T_2446;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_3 <= MultiplyAccumulate_3_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_3 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_3 <= _T_2451;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_4 <= MultiplyAccumulate_4_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_4 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_4 <= _T_2456;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_5 <= MultiplyAccumulate_5_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_5 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_5 <= _T_2461;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_6 <= MultiplyAccumulate_6_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_6 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_6 <= _T_2466;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_7 <= MultiplyAccumulate_7_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_7 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_7 <= _T_2471;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_8 <= MultiplyAccumulate_8_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_8 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_8 <= _T_2476;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_9 <= MultiplyAccumulate_9_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_9 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_9 <= _T_2481;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_10 <= MultiplyAccumulate_10_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_10 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_10 <= _T_2486;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_11 <= MultiplyAccumulate_11_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_11 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_11 <= _T_2491;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_12 <= MultiplyAccumulate_12_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_12 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_12 <= _T_2496;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_13 <= MultiplyAccumulate_13_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_13 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_13 <= _T_2501;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_14 <= MultiplyAccumulate_14_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_14 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_14 <= _T_2506;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_15 <= MultiplyAccumulate_15_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_15 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_15 <= _T_2511;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_16 <= MultiplyAccumulate_16_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_16 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_16 <= _T_2516;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_17 <= MultiplyAccumulate_17_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_17 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_17 <= _T_2521;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_18 <= MultiplyAccumulate_18_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_18 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_18 <= _T_2526;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_19 <= MultiplyAccumulate_19_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_19 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_19 <= _T_2531;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_20 <= MultiplyAccumulate_20_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_20 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_20 <= _T_2536;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_21 <= MultiplyAccumulate_21_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_21 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_21 <= _T_2541;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_22 <= MultiplyAccumulate_22_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_22 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_22 <= _T_2546;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_23 <= MultiplyAccumulate_23_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_23 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_23 <= _T_2551;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_24 <= MultiplyAccumulate_24_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_24 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_24 <= _T_2556;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_25 <= MultiplyAccumulate_25_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_25 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_25 <= _T_2561;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_26 <= MultiplyAccumulate_26_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_26 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_26 <= _T_2566;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_27 <= MultiplyAccumulate_27_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_27 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_27 <= _T_2571;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_28 <= MultiplyAccumulate_28_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_28 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_28 <= _T_2576;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_29 <= MultiplyAccumulate_29_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_29 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_29 <= _T_2581;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_30 <= MultiplyAccumulate_30_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_30 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_30 <= _T_2586;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_31 <= MultiplyAccumulate_31_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_31 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_31 <= _T_2591;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_32 <= MultiplyAccumulate_32_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_32 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_32 <= _T_2596;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_33 <= MultiplyAccumulate_33_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_33 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_33 <= _T_2601;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_34 <= MultiplyAccumulate_34_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_34 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_34 <= _T_2606;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_35 <= MultiplyAccumulate_35_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_35 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_35 <= _T_2611;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_36 <= MultiplyAccumulate_36_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_36 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_36 <= _T_2616;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_37 <= MultiplyAccumulate_37_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_37 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_37 <= _T_2621;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_38 <= MultiplyAccumulate_38_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_38 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_38 <= _T_2626;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_39 <= MultiplyAccumulate_39_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_39 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_39 <= _T_2631;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_40 <= MultiplyAccumulate_40_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_40 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_40 <= _T_2636;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_41 <= MultiplyAccumulate_41_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_41 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_41 <= _T_2641;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_42 <= MultiplyAccumulate_42_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_42 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_42 <= _T_2646;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_43 <= MultiplyAccumulate_43_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_43 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_43 <= _T_2651;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_44 <= MultiplyAccumulate_44_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_44 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_44 <= _T_2656;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_45 <= MultiplyAccumulate_45_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_45 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_45 <= _T_2661;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_46 <= MultiplyAccumulate_46_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_46 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_46 <= _T_2666;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_47 <= MultiplyAccumulate_47_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_47 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_47 <= _T_2671;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_48 <= MultiplyAccumulate_48_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_48 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_48 <= _T_2676;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_49 <= MultiplyAccumulate_49_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_49 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_49 <= _T_2681;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_50 <= MultiplyAccumulate_50_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_50 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_50 <= _T_2686;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_51 <= MultiplyAccumulate_51_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_51 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_51 <= _T_2691;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_52 <= MultiplyAccumulate_52_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_52 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_52 <= _T_2696;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_53 <= MultiplyAccumulate_53_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_53 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_53 <= _T_2701;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_54 <= MultiplyAccumulate_54_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_54 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_54 <= _T_2706;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_55 <= MultiplyAccumulate_55_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_55 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_55 <= _T_2711;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_56 <= MultiplyAccumulate_56_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_56 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_56 <= _T_2716;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_57 <= MultiplyAccumulate_57_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_57 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_57 <= _T_2721;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_58 <= MultiplyAccumulate_58_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_58 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_58 <= _T_2726;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_59 <= MultiplyAccumulate_59_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_59 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_59 <= _T_2731;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_60 <= MultiplyAccumulate_60_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_60 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_60 <= _T_2736;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_61 <= MultiplyAccumulate_61_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_61 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_61 <= _T_2741;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_62 <= MultiplyAccumulate_62_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_62 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_62 <= _T_2746;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_63 <= MultiplyAccumulate_63_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_63 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_63 <= _T_2751;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_64 <= MultiplyAccumulate_64_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_64 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_64 <= _T_2756;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_65 <= MultiplyAccumulate_65_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_65 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_65 <= _T_2761;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_66 <= MultiplyAccumulate_66_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_66 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_66 <= _T_2766;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_67 <= MultiplyAccumulate_67_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_67 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_67 <= _T_2771;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_68 <= MultiplyAccumulate_68_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_68 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_68 <= _T_2776;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_69 <= MultiplyAccumulate_69_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_69 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_69 <= _T_2781;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_70 <= MultiplyAccumulate_70_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_70 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_70 <= _T_2786;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_71 <= MultiplyAccumulate_71_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_71 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_71 <= _T_2791;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_72 <= MultiplyAccumulate_72_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_72 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_72 <= _T_2796;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_73 <= MultiplyAccumulate_73_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_73 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_73 <= _T_2801;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_74 <= MultiplyAccumulate_74_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_74 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_74 <= _T_2806;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_75 <= MultiplyAccumulate_75_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_75 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_75 <= _T_2811;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_76 <= MultiplyAccumulate_76_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_76 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_76 <= _T_2816;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_77 <= MultiplyAccumulate_77_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_77 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_77 <= _T_2821;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_78 <= MultiplyAccumulate_78_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_78 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_78 <= _T_2826;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_79 <= MultiplyAccumulate_79_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_79 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_79 <= _T_2831;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_80 <= MultiplyAccumulate_80_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_80 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_80 <= _T_2836;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_81 <= MultiplyAccumulate_81_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_81 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_81 <= _T_2841;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_82 <= MultiplyAccumulate_82_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_82 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_82 <= _T_2846;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_83 <= MultiplyAccumulate_83_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_83 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_83 <= _T_2851;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_84 <= MultiplyAccumulate_84_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_84 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_84 <= _T_2856;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_85 <= MultiplyAccumulate_85_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_85 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_85 <= _T_2861;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_86 <= MultiplyAccumulate_86_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_86 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_86 <= _T_2866;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_87 <= MultiplyAccumulate_87_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_87 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_87 <= _T_2871;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_88 <= MultiplyAccumulate_88_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_88 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_88 <= _T_2876;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_89 <= MultiplyAccumulate_89_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_89 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_89 <= _T_2881;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_90 <= MultiplyAccumulate_90_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_90 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_90 <= _T_2886;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_91 <= MultiplyAccumulate_91_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_91 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_91 <= _T_2891;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_92 <= MultiplyAccumulate_92_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_92 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_92 <= _T_2896;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_93 <= MultiplyAccumulate_93_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_93 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_93 <= _T_2901;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_94 <= MultiplyAccumulate_94_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_94 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_94 <= _T_2906;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_95 <= MultiplyAccumulate_95_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_95 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_95 <= _T_2911;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_96 <= MultiplyAccumulate_96_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_96 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_96 <= _T_2916;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_97 <= MultiplyAccumulate_97_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_97 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_97 <= _T_2921;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_98 <= MultiplyAccumulate_98_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_98 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_98 <= _T_2926;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_99 <= MultiplyAccumulate_99_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_99 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_99 <= _T_2931;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_100 <= MultiplyAccumulate_100_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_100 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_100 <= _T_2936;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_101 <= MultiplyAccumulate_101_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_101 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_101 <= _T_2941;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_102 <= MultiplyAccumulate_102_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_102 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_102 <= _T_2946;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_103 <= MultiplyAccumulate_103_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_103 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_103 <= _T_2951;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_104 <= MultiplyAccumulate_104_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_104 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_104 <= _T_2956;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_105 <= MultiplyAccumulate_105_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_105 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_105 <= _T_2961;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_106 <= MultiplyAccumulate_106_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_106 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_106 <= _T_2966;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_107 <= MultiplyAccumulate_107_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_107 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_107 <= _T_2971;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_108 <= MultiplyAccumulate_108_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_108 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_108 <= _T_2976;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_109 <= MultiplyAccumulate_109_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_109 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_109 <= _T_2981;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_110 <= MultiplyAccumulate_110_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_110 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_110 <= _T_2986;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_111 <= MultiplyAccumulate_111_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_111 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_111 <= _T_2991;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_112 <= MultiplyAccumulate_112_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_112 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_112 <= _T_2996;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_113 <= MultiplyAccumulate_113_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_113 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_113 <= _T_3001;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_114 <= MultiplyAccumulate_114_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_114 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_114 <= _T_3006;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_115 <= MultiplyAccumulate_115_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_115 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_115 <= _T_3011;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_116 <= MultiplyAccumulate_116_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_116 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_116 <= _T_3016;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_117 <= MultiplyAccumulate_117_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_117 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_117 <= _T_3021;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_118 <= MultiplyAccumulate_118_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_118 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_118 <= _T_3026;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_119 <= MultiplyAccumulate_119_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_119 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_119 <= _T_3031;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_120 <= MultiplyAccumulate_120_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_120 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_120 <= _T_3036;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_121 <= MultiplyAccumulate_121_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_121 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_121 <= _T_3041;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_122 <= MultiplyAccumulate_122_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_122 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_122 <= _T_3046;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_123 <= MultiplyAccumulate_123_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_123 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_123 <= _T_3051;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_124 <= MultiplyAccumulate_124_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_124 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_124 <= _T_3056;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_125 <= MultiplyAccumulate_125_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_125 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_125 <= _T_3061;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_126 <= MultiplyAccumulate_126_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_126 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_126 <= _T_3066;
        end
      end
    end
    if (_T_2438) begin
      cummulativeSums_127 <= MultiplyAccumulate_127_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_127 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_127 <= _T_3071;
        end
      end
    end
    _T_2401 <= _T_2398;
    _T_2403 <= _T_2401;
    _T_2405 <= _T_2403;
    _T_2407 <= _T_2405;
    _T_2409 <= _T_2407;
    _T_2411 <= _T_2409;
    rst <= _T_2411;
    if (reset) begin
      done <= 1'h0;
    end else begin
      if (_T_2418) begin
        done <= 1'h0;
      end else begin
        if (_T_2416) begin
          done <= 1'h1;
        end
      end
    end
    _T_2422 <= io_dataIn_valid;
    _T_2424 <= _T_2422;
    _T_2426 <= _T_2424;
    _T_2428 <= _T_2426;
    _T_2430 <= _T_2428;
    _T_2432 <= _T_2430;
    vld <= _T_2432;
  end
endmodule
module SSILayerOut(
  input         clock,
  input         reset,
  input         io_dataIn_valid,
  input  [15:0] io_dataIn_bits_0,
  input  [15:0] io_dataIn_bits_1,
  input  [15:0] io_dataIn_bits_2,
  input  [15:0] io_dataIn_bits_3,
  input  [15:0] io_dataIn_bits_4,
  input  [15:0] io_dataIn_bits_5,
  input  [15:0] io_dataIn_bits_6,
  input  [15:0] io_dataIn_bits_7,
  input  [15:0] io_dataIn_bits_8,
  input  [15:0] io_dataIn_bits_9,
  input  [15:0] io_dataIn_bits_10,
  input  [15:0] io_dataIn_bits_11,
  input  [15:0] io_dataIn_bits_12,
  input  [15:0] io_dataIn_bits_13,
  input  [15:0] io_dataIn_bits_14,
  input  [15:0] io_dataIn_bits_15,
  input  [15:0] io_dataIn_bits_16,
  input  [15:0] io_dataIn_bits_17,
  input  [15:0] io_dataIn_bits_18,
  input  [15:0] io_dataIn_bits_19,
  input  [15:0] io_dataIn_bits_20,
  input  [15:0] io_dataIn_bits_21,
  input  [15:0] io_dataIn_bits_22,
  input  [15:0] io_dataIn_bits_23,
  input  [15:0] io_dataIn_bits_24,
  input  [15:0] io_dataIn_bits_25,
  input  [15:0] io_dataIn_bits_26,
  input  [15:0] io_dataIn_bits_27,
  input  [15:0] io_dataIn_bits_28,
  input  [15:0] io_dataIn_bits_29,
  input  [15:0] io_dataIn_bits_30,
  input  [15:0] io_dataIn_bits_31,
  input  [15:0] io_dataIn_bits_32,
  input  [15:0] io_dataIn_bits_33,
  input  [15:0] io_dataIn_bits_34,
  input  [15:0] io_dataIn_bits_35,
  input  [15:0] io_dataIn_bits_36,
  input  [15:0] io_dataIn_bits_37,
  input  [15:0] io_dataIn_bits_38,
  input  [15:0] io_dataIn_bits_39,
  input  [15:0] io_dataIn_bits_40,
  input  [15:0] io_dataIn_bits_41,
  input  [15:0] io_dataIn_bits_42,
  input  [15:0] io_dataIn_bits_43,
  input  [15:0] io_dataIn_bits_44,
  input  [15:0] io_dataIn_bits_45,
  input  [15:0] io_dataIn_bits_46,
  input  [15:0] io_dataIn_bits_47,
  input  [15:0] io_dataIn_bits_48,
  input  [15:0] io_dataIn_bits_49,
  input  [15:0] io_dataIn_bits_50,
  input  [15:0] io_dataIn_bits_51,
  input  [15:0] io_dataIn_bits_52,
  input  [15:0] io_dataIn_bits_53,
  input  [15:0] io_dataIn_bits_54,
  input  [15:0] io_dataIn_bits_55,
  input  [15:0] io_dataIn_bits_56,
  input  [15:0] io_dataIn_bits_57,
  input  [15:0] io_dataIn_bits_58,
  input  [15:0] io_dataIn_bits_59,
  input  [15:0] io_dataIn_bits_60,
  input  [15:0] io_dataIn_bits_61,
  input  [15:0] io_dataIn_bits_62,
  input  [15:0] io_dataIn_bits_63,
  input  [15:0] io_dataIn_bits_64,
  input  [15:0] io_dataIn_bits_65,
  input  [15:0] io_dataIn_bits_66,
  input  [15:0] io_dataIn_bits_67,
  input  [15:0] io_dataIn_bits_68,
  input  [15:0] io_dataIn_bits_69,
  input  [15:0] io_dataIn_bits_70,
  input  [15:0] io_dataIn_bits_71,
  input  [15:0] io_dataIn_bits_72,
  input  [15:0] io_dataIn_bits_73,
  input  [15:0] io_dataIn_bits_74,
  input  [15:0] io_dataIn_bits_75,
  input  [15:0] io_dataIn_bits_76,
  input  [15:0] io_dataIn_bits_77,
  input  [15:0] io_dataIn_bits_78,
  input  [15:0] io_dataIn_bits_79,
  input  [15:0] io_dataIn_bits_80,
  input  [15:0] io_dataIn_bits_81,
  input  [15:0] io_dataIn_bits_82,
  input  [15:0] io_dataIn_bits_83,
  input  [15:0] io_dataIn_bits_84,
  input  [15:0] io_dataIn_bits_85,
  input  [15:0] io_dataIn_bits_86,
  input  [15:0] io_dataIn_bits_87,
  input  [15:0] io_dataIn_bits_88,
  input  [15:0] io_dataIn_bits_89,
  input  [15:0] io_dataIn_bits_90,
  input  [15:0] io_dataIn_bits_91,
  input  [15:0] io_dataIn_bits_92,
  input  [15:0] io_dataIn_bits_93,
  input  [15:0] io_dataIn_bits_94,
  input  [15:0] io_dataIn_bits_95,
  input  [15:0] io_dataIn_bits_96,
  input  [15:0] io_dataIn_bits_97,
  input  [15:0] io_dataIn_bits_98,
  input  [15:0] io_dataIn_bits_99,
  input  [15:0] io_dataIn_bits_100,
  input  [15:0] io_dataIn_bits_101,
  input  [15:0] io_dataIn_bits_102,
  input  [15:0] io_dataIn_bits_103,
  input  [15:0] io_dataIn_bits_104,
  input  [15:0] io_dataIn_bits_105,
  input  [15:0] io_dataIn_bits_106,
  input  [15:0] io_dataIn_bits_107,
  input  [15:0] io_dataIn_bits_108,
  input  [15:0] io_dataIn_bits_109,
  input  [15:0] io_dataIn_bits_110,
  input  [15:0] io_dataIn_bits_111,
  input  [15:0] io_dataIn_bits_112,
  input  [15:0] io_dataIn_bits_113,
  input  [15:0] io_dataIn_bits_114,
  input  [15:0] io_dataIn_bits_115,
  input  [15:0] io_dataIn_bits_116,
  input  [15:0] io_dataIn_bits_117,
  input  [15:0] io_dataIn_bits_118,
  input  [15:0] io_dataIn_bits_119,
  input  [15:0] io_dataIn_bits_120,
  input  [15:0] io_dataIn_bits_121,
  input  [15:0] io_dataIn_bits_122,
  input  [15:0] io_dataIn_bits_123,
  input  [15:0] io_dataIn_bits_124,
  input  [15:0] io_dataIn_bits_125,
  input  [15:0] io_dataIn_bits_126,
  input  [15:0] io_dataIn_bits_127,
  output        io_dataOut_valid,
  output [15:0] io_dataOut_bits_0
);
  reg [15:0] buffer_0; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_0;
  reg [15:0] buffer_1; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_1;
  reg [15:0] buffer_2; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_2;
  reg [15:0] buffer_3; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_3;
  reg [15:0] buffer_4; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_4;
  reg [15:0] buffer_5; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_5;
  reg [15:0] buffer_6; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_6;
  reg [15:0] buffer_7; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_7;
  reg [15:0] buffer_8; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_8;
  reg [15:0] buffer_9; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_9;
  reg [15:0] buffer_10; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_10;
  reg [15:0] buffer_11; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_11;
  reg [15:0] buffer_12; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_12;
  reg [15:0] buffer_13; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_13;
  reg [15:0] buffer_14; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_14;
  reg [15:0] buffer_15; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_15;
  reg [15:0] buffer_16; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_16;
  reg [15:0] buffer_17; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_17;
  reg [15:0] buffer_18; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_18;
  reg [15:0] buffer_19; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_19;
  reg [15:0] buffer_20; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_20;
  reg [15:0] buffer_21; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_21;
  reg [15:0] buffer_22; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_22;
  reg [15:0] buffer_23; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_23;
  reg [15:0] buffer_24; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_24;
  reg [15:0] buffer_25; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_25;
  reg [15:0] buffer_26; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_26;
  reg [15:0] buffer_27; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_27;
  reg [15:0] buffer_28; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_28;
  reg [15:0] buffer_29; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_29;
  reg [15:0] buffer_30; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_30;
  reg [15:0] buffer_31; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_31;
  reg [15:0] buffer_32; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_32;
  reg [15:0] buffer_33; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_33;
  reg [15:0] buffer_34; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_34;
  reg [15:0] buffer_35; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_35;
  reg [15:0] buffer_36; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_36;
  reg [15:0] buffer_37; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_37;
  reg [15:0] buffer_38; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_38;
  reg [15:0] buffer_39; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_39;
  reg [15:0] buffer_40; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_40;
  reg [15:0] buffer_41; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_41;
  reg [15:0] buffer_42; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_42;
  reg [15:0] buffer_43; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_43;
  reg [15:0] buffer_44; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_44;
  reg [15:0] buffer_45; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_45;
  reg [15:0] buffer_46; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_46;
  reg [15:0] buffer_47; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_47;
  reg [15:0] buffer_48; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_48;
  reg [15:0] buffer_49; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_49;
  reg [15:0] buffer_50; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_50;
  reg [15:0] buffer_51; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_51;
  reg [15:0] buffer_52; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_52;
  reg [15:0] buffer_53; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_53;
  reg [15:0] buffer_54; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_54;
  reg [15:0] buffer_55; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_55;
  reg [15:0] buffer_56; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_56;
  reg [15:0] buffer_57; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_57;
  reg [15:0] buffer_58; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_58;
  reg [15:0] buffer_59; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_59;
  reg [15:0] buffer_60; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_60;
  reg [15:0] buffer_61; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_61;
  reg [15:0] buffer_62; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_62;
  reg [15:0] buffer_63; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_63;
  reg [15:0] buffer_64; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_64;
  reg [15:0] buffer_65; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_65;
  reg [15:0] buffer_66; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_66;
  reg [15:0] buffer_67; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_67;
  reg [15:0] buffer_68; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_68;
  reg [15:0] buffer_69; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_69;
  reg [15:0] buffer_70; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_70;
  reg [15:0] buffer_71; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_71;
  reg [15:0] buffer_72; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_72;
  reg [15:0] buffer_73; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_73;
  reg [15:0] buffer_74; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_74;
  reg [15:0] buffer_75; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_75;
  reg [15:0] buffer_76; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_76;
  reg [15:0] buffer_77; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_77;
  reg [15:0] buffer_78; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_78;
  reg [15:0] buffer_79; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_79;
  reg [15:0] buffer_80; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_80;
  reg [15:0] buffer_81; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_81;
  reg [15:0] buffer_82; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_82;
  reg [15:0] buffer_83; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_83;
  reg [15:0] buffer_84; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_84;
  reg [15:0] buffer_85; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_85;
  reg [15:0] buffer_86; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_86;
  reg [15:0] buffer_87; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_87;
  reg [15:0] buffer_88; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_88;
  reg [15:0] buffer_89; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_89;
  reg [15:0] buffer_90; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_90;
  reg [15:0] buffer_91; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_91;
  reg [15:0] buffer_92; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_92;
  reg [15:0] buffer_93; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_93;
  reg [15:0] buffer_94; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_94;
  reg [15:0] buffer_95; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_95;
  reg [15:0] buffer_96; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_96;
  reg [15:0] buffer_97; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_97;
  reg [15:0] buffer_98; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_98;
  reg [15:0] buffer_99; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_99;
  reg [15:0] buffer_100; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_100;
  reg [15:0] buffer_101; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_101;
  reg [15:0] buffer_102; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_102;
  reg [15:0] buffer_103; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_103;
  reg [15:0] buffer_104; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_104;
  reg [15:0] buffer_105; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_105;
  reg [15:0] buffer_106; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_106;
  reg [15:0] buffer_107; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_107;
  reg [15:0] buffer_108; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_108;
  reg [15:0] buffer_109; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_109;
  reg [15:0] buffer_110; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_110;
  reg [15:0] buffer_111; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_111;
  reg [15:0] buffer_112; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_112;
  reg [15:0] buffer_113; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_113;
  reg [15:0] buffer_114; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_114;
  reg [15:0] buffer_115; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_115;
  reg [15:0] buffer_116; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_116;
  reg [15:0] buffer_117; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_117;
  reg [15:0] buffer_118; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_118;
  reg [15:0] buffer_119; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_119;
  reg [15:0] buffer_120; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_120;
  reg [15:0] buffer_121; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_121;
  reg [15:0] buffer_122; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_122;
  reg [15:0] buffer_123; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_123;
  reg [15:0] buffer_124; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_124;
  reg [15:0] buffer_125; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_125;
  reg [15:0] buffer_126; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_126;
  reg [15:0] buffer_127; // @[SSILayerOut.scala 20:10]
  reg [31:0] _RAND_127;
  reg [127:0] _T_926; // @[SSILayerOut.scala 43:24]
  reg [127:0] _RAND_128;
  wire [15:0] _GEN_0; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_1; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_2; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_3; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_4; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_5; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_6; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_7; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_8; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_9; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_10; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_11; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_12; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_13; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_14; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_15; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_16; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_17; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_18; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_19; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_20; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_21; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_22; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_23; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_24; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_25; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_26; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_27; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_28; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_29; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_30; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_31; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_32; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_33; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_34; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_35; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_36; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_37; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_38; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_39; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_40; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_41; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_42; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_43; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_44; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_45; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_46; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_47; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_48; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_49; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_50; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_51; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_52; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_53; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_54; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_55; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_56; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_57; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_58; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_59; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_60; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_61; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_62; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_63; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_64; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_65; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_66; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_67; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_68; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_69; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_70; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_71; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_72; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_73; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_74; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_75; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_76; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_77; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_78; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_79; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_80; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_81; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_82; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_83; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_84; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_85; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_86; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_87; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_88; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_89; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_90; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_91; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_92; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_93; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_94; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_95; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_96; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_97; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_98; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_99; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_100; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_101; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_102; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_103; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_104; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_105; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_106; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_107; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_108; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_109; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_110; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_111; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_112; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_113; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_114; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_115; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_116; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_117; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_118; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_119; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_120; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_121; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_122; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_123; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_124; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_125; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_126; // @[SSILayerOut.scala 37:28]
  wire [15:0] _GEN_127; // @[SSILayerOut.scala 37:28]
  wire [128:0] _GEN_129; // @[SSILayerOut.scala 44:20]
  wire [128:0] _T_927; // @[SSILayerOut.scala 44:20]
  wire [128:0] _GEN_128; // @[SSILayerOut.scala 45:30]
  wire  _T_929; // @[SSILayerOut.scala 48:30]
  assign _GEN_0 = io_dataIn_valid ? $signed(io_dataIn_bits_0) : $signed(buffer_1); // @[SSILayerOut.scala 37:28]
  assign _GEN_1 = io_dataIn_valid ? $signed(io_dataIn_bits_1) : $signed(buffer_2); // @[SSILayerOut.scala 37:28]
  assign _GEN_2 = io_dataIn_valid ? $signed(io_dataIn_bits_2) : $signed(buffer_3); // @[SSILayerOut.scala 37:28]
  assign _GEN_3 = io_dataIn_valid ? $signed(io_dataIn_bits_3) : $signed(buffer_4); // @[SSILayerOut.scala 37:28]
  assign _GEN_4 = io_dataIn_valid ? $signed(io_dataIn_bits_4) : $signed(buffer_5); // @[SSILayerOut.scala 37:28]
  assign _GEN_5 = io_dataIn_valid ? $signed(io_dataIn_bits_5) : $signed(buffer_6); // @[SSILayerOut.scala 37:28]
  assign _GEN_6 = io_dataIn_valid ? $signed(io_dataIn_bits_6) : $signed(buffer_7); // @[SSILayerOut.scala 37:28]
  assign _GEN_7 = io_dataIn_valid ? $signed(io_dataIn_bits_7) : $signed(buffer_8); // @[SSILayerOut.scala 37:28]
  assign _GEN_8 = io_dataIn_valid ? $signed(io_dataIn_bits_8) : $signed(buffer_9); // @[SSILayerOut.scala 37:28]
  assign _GEN_9 = io_dataIn_valid ? $signed(io_dataIn_bits_9) : $signed(buffer_10); // @[SSILayerOut.scala 37:28]
  assign _GEN_10 = io_dataIn_valid ? $signed(io_dataIn_bits_10) : $signed(buffer_11); // @[SSILayerOut.scala 37:28]
  assign _GEN_11 = io_dataIn_valid ? $signed(io_dataIn_bits_11) : $signed(buffer_12); // @[SSILayerOut.scala 37:28]
  assign _GEN_12 = io_dataIn_valid ? $signed(io_dataIn_bits_12) : $signed(buffer_13); // @[SSILayerOut.scala 37:28]
  assign _GEN_13 = io_dataIn_valid ? $signed(io_dataIn_bits_13) : $signed(buffer_14); // @[SSILayerOut.scala 37:28]
  assign _GEN_14 = io_dataIn_valid ? $signed(io_dataIn_bits_14) : $signed(buffer_15); // @[SSILayerOut.scala 37:28]
  assign _GEN_15 = io_dataIn_valid ? $signed(io_dataIn_bits_15) : $signed(buffer_16); // @[SSILayerOut.scala 37:28]
  assign _GEN_16 = io_dataIn_valid ? $signed(io_dataIn_bits_16) : $signed(buffer_17); // @[SSILayerOut.scala 37:28]
  assign _GEN_17 = io_dataIn_valid ? $signed(io_dataIn_bits_17) : $signed(buffer_18); // @[SSILayerOut.scala 37:28]
  assign _GEN_18 = io_dataIn_valid ? $signed(io_dataIn_bits_18) : $signed(buffer_19); // @[SSILayerOut.scala 37:28]
  assign _GEN_19 = io_dataIn_valid ? $signed(io_dataIn_bits_19) : $signed(buffer_20); // @[SSILayerOut.scala 37:28]
  assign _GEN_20 = io_dataIn_valid ? $signed(io_dataIn_bits_20) : $signed(buffer_21); // @[SSILayerOut.scala 37:28]
  assign _GEN_21 = io_dataIn_valid ? $signed(io_dataIn_bits_21) : $signed(buffer_22); // @[SSILayerOut.scala 37:28]
  assign _GEN_22 = io_dataIn_valid ? $signed(io_dataIn_bits_22) : $signed(buffer_23); // @[SSILayerOut.scala 37:28]
  assign _GEN_23 = io_dataIn_valid ? $signed(io_dataIn_bits_23) : $signed(buffer_24); // @[SSILayerOut.scala 37:28]
  assign _GEN_24 = io_dataIn_valid ? $signed(io_dataIn_bits_24) : $signed(buffer_25); // @[SSILayerOut.scala 37:28]
  assign _GEN_25 = io_dataIn_valid ? $signed(io_dataIn_bits_25) : $signed(buffer_26); // @[SSILayerOut.scala 37:28]
  assign _GEN_26 = io_dataIn_valid ? $signed(io_dataIn_bits_26) : $signed(buffer_27); // @[SSILayerOut.scala 37:28]
  assign _GEN_27 = io_dataIn_valid ? $signed(io_dataIn_bits_27) : $signed(buffer_28); // @[SSILayerOut.scala 37:28]
  assign _GEN_28 = io_dataIn_valid ? $signed(io_dataIn_bits_28) : $signed(buffer_29); // @[SSILayerOut.scala 37:28]
  assign _GEN_29 = io_dataIn_valid ? $signed(io_dataIn_bits_29) : $signed(buffer_30); // @[SSILayerOut.scala 37:28]
  assign _GEN_30 = io_dataIn_valid ? $signed(io_dataIn_bits_30) : $signed(buffer_31); // @[SSILayerOut.scala 37:28]
  assign _GEN_31 = io_dataIn_valid ? $signed(io_dataIn_bits_31) : $signed(buffer_32); // @[SSILayerOut.scala 37:28]
  assign _GEN_32 = io_dataIn_valid ? $signed(io_dataIn_bits_32) : $signed(buffer_33); // @[SSILayerOut.scala 37:28]
  assign _GEN_33 = io_dataIn_valid ? $signed(io_dataIn_bits_33) : $signed(buffer_34); // @[SSILayerOut.scala 37:28]
  assign _GEN_34 = io_dataIn_valid ? $signed(io_dataIn_bits_34) : $signed(buffer_35); // @[SSILayerOut.scala 37:28]
  assign _GEN_35 = io_dataIn_valid ? $signed(io_dataIn_bits_35) : $signed(buffer_36); // @[SSILayerOut.scala 37:28]
  assign _GEN_36 = io_dataIn_valid ? $signed(io_dataIn_bits_36) : $signed(buffer_37); // @[SSILayerOut.scala 37:28]
  assign _GEN_37 = io_dataIn_valid ? $signed(io_dataIn_bits_37) : $signed(buffer_38); // @[SSILayerOut.scala 37:28]
  assign _GEN_38 = io_dataIn_valid ? $signed(io_dataIn_bits_38) : $signed(buffer_39); // @[SSILayerOut.scala 37:28]
  assign _GEN_39 = io_dataIn_valid ? $signed(io_dataIn_bits_39) : $signed(buffer_40); // @[SSILayerOut.scala 37:28]
  assign _GEN_40 = io_dataIn_valid ? $signed(io_dataIn_bits_40) : $signed(buffer_41); // @[SSILayerOut.scala 37:28]
  assign _GEN_41 = io_dataIn_valid ? $signed(io_dataIn_bits_41) : $signed(buffer_42); // @[SSILayerOut.scala 37:28]
  assign _GEN_42 = io_dataIn_valid ? $signed(io_dataIn_bits_42) : $signed(buffer_43); // @[SSILayerOut.scala 37:28]
  assign _GEN_43 = io_dataIn_valid ? $signed(io_dataIn_bits_43) : $signed(buffer_44); // @[SSILayerOut.scala 37:28]
  assign _GEN_44 = io_dataIn_valid ? $signed(io_dataIn_bits_44) : $signed(buffer_45); // @[SSILayerOut.scala 37:28]
  assign _GEN_45 = io_dataIn_valid ? $signed(io_dataIn_bits_45) : $signed(buffer_46); // @[SSILayerOut.scala 37:28]
  assign _GEN_46 = io_dataIn_valid ? $signed(io_dataIn_bits_46) : $signed(buffer_47); // @[SSILayerOut.scala 37:28]
  assign _GEN_47 = io_dataIn_valid ? $signed(io_dataIn_bits_47) : $signed(buffer_48); // @[SSILayerOut.scala 37:28]
  assign _GEN_48 = io_dataIn_valid ? $signed(io_dataIn_bits_48) : $signed(buffer_49); // @[SSILayerOut.scala 37:28]
  assign _GEN_49 = io_dataIn_valid ? $signed(io_dataIn_bits_49) : $signed(buffer_50); // @[SSILayerOut.scala 37:28]
  assign _GEN_50 = io_dataIn_valid ? $signed(io_dataIn_bits_50) : $signed(buffer_51); // @[SSILayerOut.scala 37:28]
  assign _GEN_51 = io_dataIn_valid ? $signed(io_dataIn_bits_51) : $signed(buffer_52); // @[SSILayerOut.scala 37:28]
  assign _GEN_52 = io_dataIn_valid ? $signed(io_dataIn_bits_52) : $signed(buffer_53); // @[SSILayerOut.scala 37:28]
  assign _GEN_53 = io_dataIn_valid ? $signed(io_dataIn_bits_53) : $signed(buffer_54); // @[SSILayerOut.scala 37:28]
  assign _GEN_54 = io_dataIn_valid ? $signed(io_dataIn_bits_54) : $signed(buffer_55); // @[SSILayerOut.scala 37:28]
  assign _GEN_55 = io_dataIn_valid ? $signed(io_dataIn_bits_55) : $signed(buffer_56); // @[SSILayerOut.scala 37:28]
  assign _GEN_56 = io_dataIn_valid ? $signed(io_dataIn_bits_56) : $signed(buffer_57); // @[SSILayerOut.scala 37:28]
  assign _GEN_57 = io_dataIn_valid ? $signed(io_dataIn_bits_57) : $signed(buffer_58); // @[SSILayerOut.scala 37:28]
  assign _GEN_58 = io_dataIn_valid ? $signed(io_dataIn_bits_58) : $signed(buffer_59); // @[SSILayerOut.scala 37:28]
  assign _GEN_59 = io_dataIn_valid ? $signed(io_dataIn_bits_59) : $signed(buffer_60); // @[SSILayerOut.scala 37:28]
  assign _GEN_60 = io_dataIn_valid ? $signed(io_dataIn_bits_60) : $signed(buffer_61); // @[SSILayerOut.scala 37:28]
  assign _GEN_61 = io_dataIn_valid ? $signed(io_dataIn_bits_61) : $signed(buffer_62); // @[SSILayerOut.scala 37:28]
  assign _GEN_62 = io_dataIn_valid ? $signed(io_dataIn_bits_62) : $signed(buffer_63); // @[SSILayerOut.scala 37:28]
  assign _GEN_63 = io_dataIn_valid ? $signed(io_dataIn_bits_63) : $signed(buffer_64); // @[SSILayerOut.scala 37:28]
  assign _GEN_64 = io_dataIn_valid ? $signed(io_dataIn_bits_64) : $signed(buffer_65); // @[SSILayerOut.scala 37:28]
  assign _GEN_65 = io_dataIn_valid ? $signed(io_dataIn_bits_65) : $signed(buffer_66); // @[SSILayerOut.scala 37:28]
  assign _GEN_66 = io_dataIn_valid ? $signed(io_dataIn_bits_66) : $signed(buffer_67); // @[SSILayerOut.scala 37:28]
  assign _GEN_67 = io_dataIn_valid ? $signed(io_dataIn_bits_67) : $signed(buffer_68); // @[SSILayerOut.scala 37:28]
  assign _GEN_68 = io_dataIn_valid ? $signed(io_dataIn_bits_68) : $signed(buffer_69); // @[SSILayerOut.scala 37:28]
  assign _GEN_69 = io_dataIn_valid ? $signed(io_dataIn_bits_69) : $signed(buffer_70); // @[SSILayerOut.scala 37:28]
  assign _GEN_70 = io_dataIn_valid ? $signed(io_dataIn_bits_70) : $signed(buffer_71); // @[SSILayerOut.scala 37:28]
  assign _GEN_71 = io_dataIn_valid ? $signed(io_dataIn_bits_71) : $signed(buffer_72); // @[SSILayerOut.scala 37:28]
  assign _GEN_72 = io_dataIn_valid ? $signed(io_dataIn_bits_72) : $signed(buffer_73); // @[SSILayerOut.scala 37:28]
  assign _GEN_73 = io_dataIn_valid ? $signed(io_dataIn_bits_73) : $signed(buffer_74); // @[SSILayerOut.scala 37:28]
  assign _GEN_74 = io_dataIn_valid ? $signed(io_dataIn_bits_74) : $signed(buffer_75); // @[SSILayerOut.scala 37:28]
  assign _GEN_75 = io_dataIn_valid ? $signed(io_dataIn_bits_75) : $signed(buffer_76); // @[SSILayerOut.scala 37:28]
  assign _GEN_76 = io_dataIn_valid ? $signed(io_dataIn_bits_76) : $signed(buffer_77); // @[SSILayerOut.scala 37:28]
  assign _GEN_77 = io_dataIn_valid ? $signed(io_dataIn_bits_77) : $signed(buffer_78); // @[SSILayerOut.scala 37:28]
  assign _GEN_78 = io_dataIn_valid ? $signed(io_dataIn_bits_78) : $signed(buffer_79); // @[SSILayerOut.scala 37:28]
  assign _GEN_79 = io_dataIn_valid ? $signed(io_dataIn_bits_79) : $signed(buffer_80); // @[SSILayerOut.scala 37:28]
  assign _GEN_80 = io_dataIn_valid ? $signed(io_dataIn_bits_80) : $signed(buffer_81); // @[SSILayerOut.scala 37:28]
  assign _GEN_81 = io_dataIn_valid ? $signed(io_dataIn_bits_81) : $signed(buffer_82); // @[SSILayerOut.scala 37:28]
  assign _GEN_82 = io_dataIn_valid ? $signed(io_dataIn_bits_82) : $signed(buffer_83); // @[SSILayerOut.scala 37:28]
  assign _GEN_83 = io_dataIn_valid ? $signed(io_dataIn_bits_83) : $signed(buffer_84); // @[SSILayerOut.scala 37:28]
  assign _GEN_84 = io_dataIn_valid ? $signed(io_dataIn_bits_84) : $signed(buffer_85); // @[SSILayerOut.scala 37:28]
  assign _GEN_85 = io_dataIn_valid ? $signed(io_dataIn_bits_85) : $signed(buffer_86); // @[SSILayerOut.scala 37:28]
  assign _GEN_86 = io_dataIn_valid ? $signed(io_dataIn_bits_86) : $signed(buffer_87); // @[SSILayerOut.scala 37:28]
  assign _GEN_87 = io_dataIn_valid ? $signed(io_dataIn_bits_87) : $signed(buffer_88); // @[SSILayerOut.scala 37:28]
  assign _GEN_88 = io_dataIn_valid ? $signed(io_dataIn_bits_88) : $signed(buffer_89); // @[SSILayerOut.scala 37:28]
  assign _GEN_89 = io_dataIn_valid ? $signed(io_dataIn_bits_89) : $signed(buffer_90); // @[SSILayerOut.scala 37:28]
  assign _GEN_90 = io_dataIn_valid ? $signed(io_dataIn_bits_90) : $signed(buffer_91); // @[SSILayerOut.scala 37:28]
  assign _GEN_91 = io_dataIn_valid ? $signed(io_dataIn_bits_91) : $signed(buffer_92); // @[SSILayerOut.scala 37:28]
  assign _GEN_92 = io_dataIn_valid ? $signed(io_dataIn_bits_92) : $signed(buffer_93); // @[SSILayerOut.scala 37:28]
  assign _GEN_93 = io_dataIn_valid ? $signed(io_dataIn_bits_93) : $signed(buffer_94); // @[SSILayerOut.scala 37:28]
  assign _GEN_94 = io_dataIn_valid ? $signed(io_dataIn_bits_94) : $signed(buffer_95); // @[SSILayerOut.scala 37:28]
  assign _GEN_95 = io_dataIn_valid ? $signed(io_dataIn_bits_95) : $signed(buffer_96); // @[SSILayerOut.scala 37:28]
  assign _GEN_96 = io_dataIn_valid ? $signed(io_dataIn_bits_96) : $signed(buffer_97); // @[SSILayerOut.scala 37:28]
  assign _GEN_97 = io_dataIn_valid ? $signed(io_dataIn_bits_97) : $signed(buffer_98); // @[SSILayerOut.scala 37:28]
  assign _GEN_98 = io_dataIn_valid ? $signed(io_dataIn_bits_98) : $signed(buffer_99); // @[SSILayerOut.scala 37:28]
  assign _GEN_99 = io_dataIn_valid ? $signed(io_dataIn_bits_99) : $signed(buffer_100); // @[SSILayerOut.scala 37:28]
  assign _GEN_100 = io_dataIn_valid ? $signed(io_dataIn_bits_100) : $signed(buffer_101); // @[SSILayerOut.scala 37:28]
  assign _GEN_101 = io_dataIn_valid ? $signed(io_dataIn_bits_101) : $signed(buffer_102); // @[SSILayerOut.scala 37:28]
  assign _GEN_102 = io_dataIn_valid ? $signed(io_dataIn_bits_102) : $signed(buffer_103); // @[SSILayerOut.scala 37:28]
  assign _GEN_103 = io_dataIn_valid ? $signed(io_dataIn_bits_103) : $signed(buffer_104); // @[SSILayerOut.scala 37:28]
  assign _GEN_104 = io_dataIn_valid ? $signed(io_dataIn_bits_104) : $signed(buffer_105); // @[SSILayerOut.scala 37:28]
  assign _GEN_105 = io_dataIn_valid ? $signed(io_dataIn_bits_105) : $signed(buffer_106); // @[SSILayerOut.scala 37:28]
  assign _GEN_106 = io_dataIn_valid ? $signed(io_dataIn_bits_106) : $signed(buffer_107); // @[SSILayerOut.scala 37:28]
  assign _GEN_107 = io_dataIn_valid ? $signed(io_dataIn_bits_107) : $signed(buffer_108); // @[SSILayerOut.scala 37:28]
  assign _GEN_108 = io_dataIn_valid ? $signed(io_dataIn_bits_108) : $signed(buffer_109); // @[SSILayerOut.scala 37:28]
  assign _GEN_109 = io_dataIn_valid ? $signed(io_dataIn_bits_109) : $signed(buffer_110); // @[SSILayerOut.scala 37:28]
  assign _GEN_110 = io_dataIn_valid ? $signed(io_dataIn_bits_110) : $signed(buffer_111); // @[SSILayerOut.scala 37:28]
  assign _GEN_111 = io_dataIn_valid ? $signed(io_dataIn_bits_111) : $signed(buffer_112); // @[SSILayerOut.scala 37:28]
  assign _GEN_112 = io_dataIn_valid ? $signed(io_dataIn_bits_112) : $signed(buffer_113); // @[SSILayerOut.scala 37:28]
  assign _GEN_113 = io_dataIn_valid ? $signed(io_dataIn_bits_113) : $signed(buffer_114); // @[SSILayerOut.scala 37:28]
  assign _GEN_114 = io_dataIn_valid ? $signed(io_dataIn_bits_114) : $signed(buffer_115); // @[SSILayerOut.scala 37:28]
  assign _GEN_115 = io_dataIn_valid ? $signed(io_dataIn_bits_115) : $signed(buffer_116); // @[SSILayerOut.scala 37:28]
  assign _GEN_116 = io_dataIn_valid ? $signed(io_dataIn_bits_116) : $signed(buffer_117); // @[SSILayerOut.scala 37:28]
  assign _GEN_117 = io_dataIn_valid ? $signed(io_dataIn_bits_117) : $signed(buffer_118); // @[SSILayerOut.scala 37:28]
  assign _GEN_118 = io_dataIn_valid ? $signed(io_dataIn_bits_118) : $signed(buffer_119); // @[SSILayerOut.scala 37:28]
  assign _GEN_119 = io_dataIn_valid ? $signed(io_dataIn_bits_119) : $signed(buffer_120); // @[SSILayerOut.scala 37:28]
  assign _GEN_120 = io_dataIn_valid ? $signed(io_dataIn_bits_120) : $signed(buffer_121); // @[SSILayerOut.scala 37:28]
  assign _GEN_121 = io_dataIn_valid ? $signed(io_dataIn_bits_121) : $signed(buffer_122); // @[SSILayerOut.scala 37:28]
  assign _GEN_122 = io_dataIn_valid ? $signed(io_dataIn_bits_122) : $signed(buffer_123); // @[SSILayerOut.scala 37:28]
  assign _GEN_123 = io_dataIn_valid ? $signed(io_dataIn_bits_123) : $signed(buffer_124); // @[SSILayerOut.scala 37:28]
  assign _GEN_124 = io_dataIn_valid ? $signed(io_dataIn_bits_124) : $signed(buffer_125); // @[SSILayerOut.scala 37:28]
  assign _GEN_125 = io_dataIn_valid ? $signed(io_dataIn_bits_125) : $signed(buffer_126); // @[SSILayerOut.scala 37:28]
  assign _GEN_126 = io_dataIn_valid ? $signed(io_dataIn_bits_126) : $signed(buffer_127); // @[SSILayerOut.scala 37:28]
  assign _GEN_127 = io_dataIn_valid ? $signed(io_dataIn_bits_127) : $signed(buffer_127); // @[SSILayerOut.scala 37:28]
  assign _GEN_129 = {{1'd0}, _T_926}; // @[SSILayerOut.scala 44:20]
  assign _T_927 = _GEN_129 << 1; // @[SSILayerOut.scala 44:20]
  assign _GEN_128 = io_dataIn_valid ? 129'hffffffffffffffffffffffffffffffff : _T_927; // @[SSILayerOut.scala 45:30]
  assign _T_929 = _T_926[127]; // @[SSILayerOut.scala 48:30]
  assign io_dataOut_valid = _T_929;
  assign io_dataOut_bits_0 = buffer_0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  buffer_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  buffer_1 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  buffer_2 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  buffer_3 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  buffer_4 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  buffer_5 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  buffer_6 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  buffer_7 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  buffer_8 = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  buffer_9 = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  buffer_10 = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  buffer_11 = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  buffer_12 = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  buffer_13 = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  buffer_14 = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  buffer_15 = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  buffer_16 = _RAND_16[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  buffer_17 = _RAND_17[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  buffer_18 = _RAND_18[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  buffer_19 = _RAND_19[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  buffer_20 = _RAND_20[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  buffer_21 = _RAND_21[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  buffer_22 = _RAND_22[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  buffer_23 = _RAND_23[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  buffer_24 = _RAND_24[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  buffer_25 = _RAND_25[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  buffer_26 = _RAND_26[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  buffer_27 = _RAND_27[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  buffer_28 = _RAND_28[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  buffer_29 = _RAND_29[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  buffer_30 = _RAND_30[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  buffer_31 = _RAND_31[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  buffer_32 = _RAND_32[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{$random}};
  buffer_33 = _RAND_33[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{$random}};
  buffer_34 = _RAND_34[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{$random}};
  buffer_35 = _RAND_35[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{$random}};
  buffer_36 = _RAND_36[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{$random}};
  buffer_37 = _RAND_37[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{$random}};
  buffer_38 = _RAND_38[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{$random}};
  buffer_39 = _RAND_39[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{$random}};
  buffer_40 = _RAND_40[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{$random}};
  buffer_41 = _RAND_41[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{$random}};
  buffer_42 = _RAND_42[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{$random}};
  buffer_43 = _RAND_43[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{$random}};
  buffer_44 = _RAND_44[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{$random}};
  buffer_45 = _RAND_45[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{$random}};
  buffer_46 = _RAND_46[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{$random}};
  buffer_47 = _RAND_47[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{$random}};
  buffer_48 = _RAND_48[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{$random}};
  buffer_49 = _RAND_49[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{$random}};
  buffer_50 = _RAND_50[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{$random}};
  buffer_51 = _RAND_51[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{$random}};
  buffer_52 = _RAND_52[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{$random}};
  buffer_53 = _RAND_53[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{$random}};
  buffer_54 = _RAND_54[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{$random}};
  buffer_55 = _RAND_55[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{$random}};
  buffer_56 = _RAND_56[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{$random}};
  buffer_57 = _RAND_57[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{$random}};
  buffer_58 = _RAND_58[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{$random}};
  buffer_59 = _RAND_59[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{$random}};
  buffer_60 = _RAND_60[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{$random}};
  buffer_61 = _RAND_61[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{$random}};
  buffer_62 = _RAND_62[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{$random}};
  buffer_63 = _RAND_63[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{$random}};
  buffer_64 = _RAND_64[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{$random}};
  buffer_65 = _RAND_65[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{$random}};
  buffer_66 = _RAND_66[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{$random}};
  buffer_67 = _RAND_67[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{$random}};
  buffer_68 = _RAND_68[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{$random}};
  buffer_69 = _RAND_69[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{$random}};
  buffer_70 = _RAND_70[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{$random}};
  buffer_71 = _RAND_71[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{$random}};
  buffer_72 = _RAND_72[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{$random}};
  buffer_73 = _RAND_73[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{$random}};
  buffer_74 = _RAND_74[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{$random}};
  buffer_75 = _RAND_75[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{$random}};
  buffer_76 = _RAND_76[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{$random}};
  buffer_77 = _RAND_77[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{$random}};
  buffer_78 = _RAND_78[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{$random}};
  buffer_79 = _RAND_79[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{$random}};
  buffer_80 = _RAND_80[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{$random}};
  buffer_81 = _RAND_81[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{$random}};
  buffer_82 = _RAND_82[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{$random}};
  buffer_83 = _RAND_83[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{$random}};
  buffer_84 = _RAND_84[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{$random}};
  buffer_85 = _RAND_85[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{$random}};
  buffer_86 = _RAND_86[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{$random}};
  buffer_87 = _RAND_87[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{$random}};
  buffer_88 = _RAND_88[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{$random}};
  buffer_89 = _RAND_89[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{$random}};
  buffer_90 = _RAND_90[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{$random}};
  buffer_91 = _RAND_91[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{$random}};
  buffer_92 = _RAND_92[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{$random}};
  buffer_93 = _RAND_93[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{$random}};
  buffer_94 = _RAND_94[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{$random}};
  buffer_95 = _RAND_95[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{$random}};
  buffer_96 = _RAND_96[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{$random}};
  buffer_97 = _RAND_97[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{$random}};
  buffer_98 = _RAND_98[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{$random}};
  buffer_99 = _RAND_99[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{$random}};
  buffer_100 = _RAND_100[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{$random}};
  buffer_101 = _RAND_101[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{$random}};
  buffer_102 = _RAND_102[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{$random}};
  buffer_103 = _RAND_103[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{$random}};
  buffer_104 = _RAND_104[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{$random}};
  buffer_105 = _RAND_105[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{$random}};
  buffer_106 = _RAND_106[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{$random}};
  buffer_107 = _RAND_107[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{$random}};
  buffer_108 = _RAND_108[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{$random}};
  buffer_109 = _RAND_109[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{$random}};
  buffer_110 = _RAND_110[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{$random}};
  buffer_111 = _RAND_111[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{$random}};
  buffer_112 = _RAND_112[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{$random}};
  buffer_113 = _RAND_113[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{$random}};
  buffer_114 = _RAND_114[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{$random}};
  buffer_115 = _RAND_115[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{$random}};
  buffer_116 = _RAND_116[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{$random}};
  buffer_117 = _RAND_117[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{$random}};
  buffer_118 = _RAND_118[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{$random}};
  buffer_119 = _RAND_119[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{$random}};
  buffer_120 = _RAND_120[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{$random}};
  buffer_121 = _RAND_121[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{$random}};
  buffer_122 = _RAND_122[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{$random}};
  buffer_123 = _RAND_123[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{$random}};
  buffer_124 = _RAND_124[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{$random}};
  buffer_125 = _RAND_125[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{$random}};
  buffer_126 = _RAND_126[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{$random}};
  buffer_127 = _RAND_127[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {4{$random}};
  _T_926 = _RAND_128[127:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (io_dataIn_valid) begin
      buffer_0 <= io_dataIn_bits_0;
    end else begin
      buffer_0 <= buffer_1;
    end
    if (io_dataIn_valid) begin
      buffer_1 <= io_dataIn_bits_1;
    end else begin
      buffer_1 <= buffer_2;
    end
    if (io_dataIn_valid) begin
      buffer_2 <= io_dataIn_bits_2;
    end else begin
      buffer_2 <= buffer_3;
    end
    if (io_dataIn_valid) begin
      buffer_3 <= io_dataIn_bits_3;
    end else begin
      buffer_3 <= buffer_4;
    end
    if (io_dataIn_valid) begin
      buffer_4 <= io_dataIn_bits_4;
    end else begin
      buffer_4 <= buffer_5;
    end
    if (io_dataIn_valid) begin
      buffer_5 <= io_dataIn_bits_5;
    end else begin
      buffer_5 <= buffer_6;
    end
    if (io_dataIn_valid) begin
      buffer_6 <= io_dataIn_bits_6;
    end else begin
      buffer_6 <= buffer_7;
    end
    if (io_dataIn_valid) begin
      buffer_7 <= io_dataIn_bits_7;
    end else begin
      buffer_7 <= buffer_8;
    end
    if (io_dataIn_valid) begin
      buffer_8 <= io_dataIn_bits_8;
    end else begin
      buffer_8 <= buffer_9;
    end
    if (io_dataIn_valid) begin
      buffer_9 <= io_dataIn_bits_9;
    end else begin
      buffer_9 <= buffer_10;
    end
    if (io_dataIn_valid) begin
      buffer_10 <= io_dataIn_bits_10;
    end else begin
      buffer_10 <= buffer_11;
    end
    if (io_dataIn_valid) begin
      buffer_11 <= io_dataIn_bits_11;
    end else begin
      buffer_11 <= buffer_12;
    end
    if (io_dataIn_valid) begin
      buffer_12 <= io_dataIn_bits_12;
    end else begin
      buffer_12 <= buffer_13;
    end
    if (io_dataIn_valid) begin
      buffer_13 <= io_dataIn_bits_13;
    end else begin
      buffer_13 <= buffer_14;
    end
    if (io_dataIn_valid) begin
      buffer_14 <= io_dataIn_bits_14;
    end else begin
      buffer_14 <= buffer_15;
    end
    if (io_dataIn_valid) begin
      buffer_15 <= io_dataIn_bits_15;
    end else begin
      buffer_15 <= buffer_16;
    end
    if (io_dataIn_valid) begin
      buffer_16 <= io_dataIn_bits_16;
    end else begin
      buffer_16 <= buffer_17;
    end
    if (io_dataIn_valid) begin
      buffer_17 <= io_dataIn_bits_17;
    end else begin
      buffer_17 <= buffer_18;
    end
    if (io_dataIn_valid) begin
      buffer_18 <= io_dataIn_bits_18;
    end else begin
      buffer_18 <= buffer_19;
    end
    if (io_dataIn_valid) begin
      buffer_19 <= io_dataIn_bits_19;
    end else begin
      buffer_19 <= buffer_20;
    end
    if (io_dataIn_valid) begin
      buffer_20 <= io_dataIn_bits_20;
    end else begin
      buffer_20 <= buffer_21;
    end
    if (io_dataIn_valid) begin
      buffer_21 <= io_dataIn_bits_21;
    end else begin
      buffer_21 <= buffer_22;
    end
    if (io_dataIn_valid) begin
      buffer_22 <= io_dataIn_bits_22;
    end else begin
      buffer_22 <= buffer_23;
    end
    if (io_dataIn_valid) begin
      buffer_23 <= io_dataIn_bits_23;
    end else begin
      buffer_23 <= buffer_24;
    end
    if (io_dataIn_valid) begin
      buffer_24 <= io_dataIn_bits_24;
    end else begin
      buffer_24 <= buffer_25;
    end
    if (io_dataIn_valid) begin
      buffer_25 <= io_dataIn_bits_25;
    end else begin
      buffer_25 <= buffer_26;
    end
    if (io_dataIn_valid) begin
      buffer_26 <= io_dataIn_bits_26;
    end else begin
      buffer_26 <= buffer_27;
    end
    if (io_dataIn_valid) begin
      buffer_27 <= io_dataIn_bits_27;
    end else begin
      buffer_27 <= buffer_28;
    end
    if (io_dataIn_valid) begin
      buffer_28 <= io_dataIn_bits_28;
    end else begin
      buffer_28 <= buffer_29;
    end
    if (io_dataIn_valid) begin
      buffer_29 <= io_dataIn_bits_29;
    end else begin
      buffer_29 <= buffer_30;
    end
    if (io_dataIn_valid) begin
      buffer_30 <= io_dataIn_bits_30;
    end else begin
      buffer_30 <= buffer_31;
    end
    if (io_dataIn_valid) begin
      buffer_31 <= io_dataIn_bits_31;
    end else begin
      buffer_31 <= buffer_32;
    end
    if (io_dataIn_valid) begin
      buffer_32 <= io_dataIn_bits_32;
    end else begin
      buffer_32 <= buffer_33;
    end
    if (io_dataIn_valid) begin
      buffer_33 <= io_dataIn_bits_33;
    end else begin
      buffer_33 <= buffer_34;
    end
    if (io_dataIn_valid) begin
      buffer_34 <= io_dataIn_bits_34;
    end else begin
      buffer_34 <= buffer_35;
    end
    if (io_dataIn_valid) begin
      buffer_35 <= io_dataIn_bits_35;
    end else begin
      buffer_35 <= buffer_36;
    end
    if (io_dataIn_valid) begin
      buffer_36 <= io_dataIn_bits_36;
    end else begin
      buffer_36 <= buffer_37;
    end
    if (io_dataIn_valid) begin
      buffer_37 <= io_dataIn_bits_37;
    end else begin
      buffer_37 <= buffer_38;
    end
    if (io_dataIn_valid) begin
      buffer_38 <= io_dataIn_bits_38;
    end else begin
      buffer_38 <= buffer_39;
    end
    if (io_dataIn_valid) begin
      buffer_39 <= io_dataIn_bits_39;
    end else begin
      buffer_39 <= buffer_40;
    end
    if (io_dataIn_valid) begin
      buffer_40 <= io_dataIn_bits_40;
    end else begin
      buffer_40 <= buffer_41;
    end
    if (io_dataIn_valid) begin
      buffer_41 <= io_dataIn_bits_41;
    end else begin
      buffer_41 <= buffer_42;
    end
    if (io_dataIn_valid) begin
      buffer_42 <= io_dataIn_bits_42;
    end else begin
      buffer_42 <= buffer_43;
    end
    if (io_dataIn_valid) begin
      buffer_43 <= io_dataIn_bits_43;
    end else begin
      buffer_43 <= buffer_44;
    end
    if (io_dataIn_valid) begin
      buffer_44 <= io_dataIn_bits_44;
    end else begin
      buffer_44 <= buffer_45;
    end
    if (io_dataIn_valid) begin
      buffer_45 <= io_dataIn_bits_45;
    end else begin
      buffer_45 <= buffer_46;
    end
    if (io_dataIn_valid) begin
      buffer_46 <= io_dataIn_bits_46;
    end else begin
      buffer_46 <= buffer_47;
    end
    if (io_dataIn_valid) begin
      buffer_47 <= io_dataIn_bits_47;
    end else begin
      buffer_47 <= buffer_48;
    end
    if (io_dataIn_valid) begin
      buffer_48 <= io_dataIn_bits_48;
    end else begin
      buffer_48 <= buffer_49;
    end
    if (io_dataIn_valid) begin
      buffer_49 <= io_dataIn_bits_49;
    end else begin
      buffer_49 <= buffer_50;
    end
    if (io_dataIn_valid) begin
      buffer_50 <= io_dataIn_bits_50;
    end else begin
      buffer_50 <= buffer_51;
    end
    if (io_dataIn_valid) begin
      buffer_51 <= io_dataIn_bits_51;
    end else begin
      buffer_51 <= buffer_52;
    end
    if (io_dataIn_valid) begin
      buffer_52 <= io_dataIn_bits_52;
    end else begin
      buffer_52 <= buffer_53;
    end
    if (io_dataIn_valid) begin
      buffer_53 <= io_dataIn_bits_53;
    end else begin
      buffer_53 <= buffer_54;
    end
    if (io_dataIn_valid) begin
      buffer_54 <= io_dataIn_bits_54;
    end else begin
      buffer_54 <= buffer_55;
    end
    if (io_dataIn_valid) begin
      buffer_55 <= io_dataIn_bits_55;
    end else begin
      buffer_55 <= buffer_56;
    end
    if (io_dataIn_valid) begin
      buffer_56 <= io_dataIn_bits_56;
    end else begin
      buffer_56 <= buffer_57;
    end
    if (io_dataIn_valid) begin
      buffer_57 <= io_dataIn_bits_57;
    end else begin
      buffer_57 <= buffer_58;
    end
    if (io_dataIn_valid) begin
      buffer_58 <= io_dataIn_bits_58;
    end else begin
      buffer_58 <= buffer_59;
    end
    if (io_dataIn_valid) begin
      buffer_59 <= io_dataIn_bits_59;
    end else begin
      buffer_59 <= buffer_60;
    end
    if (io_dataIn_valid) begin
      buffer_60 <= io_dataIn_bits_60;
    end else begin
      buffer_60 <= buffer_61;
    end
    if (io_dataIn_valid) begin
      buffer_61 <= io_dataIn_bits_61;
    end else begin
      buffer_61 <= buffer_62;
    end
    if (io_dataIn_valid) begin
      buffer_62 <= io_dataIn_bits_62;
    end else begin
      buffer_62 <= buffer_63;
    end
    if (io_dataIn_valid) begin
      buffer_63 <= io_dataIn_bits_63;
    end else begin
      buffer_63 <= buffer_64;
    end
    if (io_dataIn_valid) begin
      buffer_64 <= io_dataIn_bits_64;
    end else begin
      buffer_64 <= buffer_65;
    end
    if (io_dataIn_valid) begin
      buffer_65 <= io_dataIn_bits_65;
    end else begin
      buffer_65 <= buffer_66;
    end
    if (io_dataIn_valid) begin
      buffer_66 <= io_dataIn_bits_66;
    end else begin
      buffer_66 <= buffer_67;
    end
    if (io_dataIn_valid) begin
      buffer_67 <= io_dataIn_bits_67;
    end else begin
      buffer_67 <= buffer_68;
    end
    if (io_dataIn_valid) begin
      buffer_68 <= io_dataIn_bits_68;
    end else begin
      buffer_68 <= buffer_69;
    end
    if (io_dataIn_valid) begin
      buffer_69 <= io_dataIn_bits_69;
    end else begin
      buffer_69 <= buffer_70;
    end
    if (io_dataIn_valid) begin
      buffer_70 <= io_dataIn_bits_70;
    end else begin
      buffer_70 <= buffer_71;
    end
    if (io_dataIn_valid) begin
      buffer_71 <= io_dataIn_bits_71;
    end else begin
      buffer_71 <= buffer_72;
    end
    if (io_dataIn_valid) begin
      buffer_72 <= io_dataIn_bits_72;
    end else begin
      buffer_72 <= buffer_73;
    end
    if (io_dataIn_valid) begin
      buffer_73 <= io_dataIn_bits_73;
    end else begin
      buffer_73 <= buffer_74;
    end
    if (io_dataIn_valid) begin
      buffer_74 <= io_dataIn_bits_74;
    end else begin
      buffer_74 <= buffer_75;
    end
    if (io_dataIn_valid) begin
      buffer_75 <= io_dataIn_bits_75;
    end else begin
      buffer_75 <= buffer_76;
    end
    if (io_dataIn_valid) begin
      buffer_76 <= io_dataIn_bits_76;
    end else begin
      buffer_76 <= buffer_77;
    end
    if (io_dataIn_valid) begin
      buffer_77 <= io_dataIn_bits_77;
    end else begin
      buffer_77 <= buffer_78;
    end
    if (io_dataIn_valid) begin
      buffer_78 <= io_dataIn_bits_78;
    end else begin
      buffer_78 <= buffer_79;
    end
    if (io_dataIn_valid) begin
      buffer_79 <= io_dataIn_bits_79;
    end else begin
      buffer_79 <= buffer_80;
    end
    if (io_dataIn_valid) begin
      buffer_80 <= io_dataIn_bits_80;
    end else begin
      buffer_80 <= buffer_81;
    end
    if (io_dataIn_valid) begin
      buffer_81 <= io_dataIn_bits_81;
    end else begin
      buffer_81 <= buffer_82;
    end
    if (io_dataIn_valid) begin
      buffer_82 <= io_dataIn_bits_82;
    end else begin
      buffer_82 <= buffer_83;
    end
    if (io_dataIn_valid) begin
      buffer_83 <= io_dataIn_bits_83;
    end else begin
      buffer_83 <= buffer_84;
    end
    if (io_dataIn_valid) begin
      buffer_84 <= io_dataIn_bits_84;
    end else begin
      buffer_84 <= buffer_85;
    end
    if (io_dataIn_valid) begin
      buffer_85 <= io_dataIn_bits_85;
    end else begin
      buffer_85 <= buffer_86;
    end
    if (io_dataIn_valid) begin
      buffer_86 <= io_dataIn_bits_86;
    end else begin
      buffer_86 <= buffer_87;
    end
    if (io_dataIn_valid) begin
      buffer_87 <= io_dataIn_bits_87;
    end else begin
      buffer_87 <= buffer_88;
    end
    if (io_dataIn_valid) begin
      buffer_88 <= io_dataIn_bits_88;
    end else begin
      buffer_88 <= buffer_89;
    end
    if (io_dataIn_valid) begin
      buffer_89 <= io_dataIn_bits_89;
    end else begin
      buffer_89 <= buffer_90;
    end
    if (io_dataIn_valid) begin
      buffer_90 <= io_dataIn_bits_90;
    end else begin
      buffer_90 <= buffer_91;
    end
    if (io_dataIn_valid) begin
      buffer_91 <= io_dataIn_bits_91;
    end else begin
      buffer_91 <= buffer_92;
    end
    if (io_dataIn_valid) begin
      buffer_92 <= io_dataIn_bits_92;
    end else begin
      buffer_92 <= buffer_93;
    end
    if (io_dataIn_valid) begin
      buffer_93 <= io_dataIn_bits_93;
    end else begin
      buffer_93 <= buffer_94;
    end
    if (io_dataIn_valid) begin
      buffer_94 <= io_dataIn_bits_94;
    end else begin
      buffer_94 <= buffer_95;
    end
    if (io_dataIn_valid) begin
      buffer_95 <= io_dataIn_bits_95;
    end else begin
      buffer_95 <= buffer_96;
    end
    if (io_dataIn_valid) begin
      buffer_96 <= io_dataIn_bits_96;
    end else begin
      buffer_96 <= buffer_97;
    end
    if (io_dataIn_valid) begin
      buffer_97 <= io_dataIn_bits_97;
    end else begin
      buffer_97 <= buffer_98;
    end
    if (io_dataIn_valid) begin
      buffer_98 <= io_dataIn_bits_98;
    end else begin
      buffer_98 <= buffer_99;
    end
    if (io_dataIn_valid) begin
      buffer_99 <= io_dataIn_bits_99;
    end else begin
      buffer_99 <= buffer_100;
    end
    if (io_dataIn_valid) begin
      buffer_100 <= io_dataIn_bits_100;
    end else begin
      buffer_100 <= buffer_101;
    end
    if (io_dataIn_valid) begin
      buffer_101 <= io_dataIn_bits_101;
    end else begin
      buffer_101 <= buffer_102;
    end
    if (io_dataIn_valid) begin
      buffer_102 <= io_dataIn_bits_102;
    end else begin
      buffer_102 <= buffer_103;
    end
    if (io_dataIn_valid) begin
      buffer_103 <= io_dataIn_bits_103;
    end else begin
      buffer_103 <= buffer_104;
    end
    if (io_dataIn_valid) begin
      buffer_104 <= io_dataIn_bits_104;
    end else begin
      buffer_104 <= buffer_105;
    end
    if (io_dataIn_valid) begin
      buffer_105 <= io_dataIn_bits_105;
    end else begin
      buffer_105 <= buffer_106;
    end
    if (io_dataIn_valid) begin
      buffer_106 <= io_dataIn_bits_106;
    end else begin
      buffer_106 <= buffer_107;
    end
    if (io_dataIn_valid) begin
      buffer_107 <= io_dataIn_bits_107;
    end else begin
      buffer_107 <= buffer_108;
    end
    if (io_dataIn_valid) begin
      buffer_108 <= io_dataIn_bits_108;
    end else begin
      buffer_108 <= buffer_109;
    end
    if (io_dataIn_valid) begin
      buffer_109 <= io_dataIn_bits_109;
    end else begin
      buffer_109 <= buffer_110;
    end
    if (io_dataIn_valid) begin
      buffer_110 <= io_dataIn_bits_110;
    end else begin
      buffer_110 <= buffer_111;
    end
    if (io_dataIn_valid) begin
      buffer_111 <= io_dataIn_bits_111;
    end else begin
      buffer_111 <= buffer_112;
    end
    if (io_dataIn_valid) begin
      buffer_112 <= io_dataIn_bits_112;
    end else begin
      buffer_112 <= buffer_113;
    end
    if (io_dataIn_valid) begin
      buffer_113 <= io_dataIn_bits_113;
    end else begin
      buffer_113 <= buffer_114;
    end
    if (io_dataIn_valid) begin
      buffer_114 <= io_dataIn_bits_114;
    end else begin
      buffer_114 <= buffer_115;
    end
    if (io_dataIn_valid) begin
      buffer_115 <= io_dataIn_bits_115;
    end else begin
      buffer_115 <= buffer_116;
    end
    if (io_dataIn_valid) begin
      buffer_116 <= io_dataIn_bits_116;
    end else begin
      buffer_116 <= buffer_117;
    end
    if (io_dataIn_valid) begin
      buffer_117 <= io_dataIn_bits_117;
    end else begin
      buffer_117 <= buffer_118;
    end
    if (io_dataIn_valid) begin
      buffer_118 <= io_dataIn_bits_118;
    end else begin
      buffer_118 <= buffer_119;
    end
    if (io_dataIn_valid) begin
      buffer_119 <= io_dataIn_bits_119;
    end else begin
      buffer_119 <= buffer_120;
    end
    if (io_dataIn_valid) begin
      buffer_120 <= io_dataIn_bits_120;
    end else begin
      buffer_120 <= buffer_121;
    end
    if (io_dataIn_valid) begin
      buffer_121 <= io_dataIn_bits_121;
    end else begin
      buffer_121 <= buffer_122;
    end
    if (io_dataIn_valid) begin
      buffer_122 <= io_dataIn_bits_122;
    end else begin
      buffer_122 <= buffer_123;
    end
    if (io_dataIn_valid) begin
      buffer_123 <= io_dataIn_bits_123;
    end else begin
      buffer_123 <= buffer_124;
    end
    if (io_dataIn_valid) begin
      buffer_124 <= io_dataIn_bits_124;
    end else begin
      buffer_124 <= buffer_125;
    end
    if (io_dataIn_valid) begin
      buffer_125 <= io_dataIn_bits_125;
    end else begin
      buffer_125 <= buffer_126;
    end
    if (io_dataIn_valid) begin
      buffer_126 <= io_dataIn_bits_126;
    end else begin
      buffer_126 <= buffer_127;
    end
    if (io_dataIn_valid) begin
      buffer_127 <= io_dataIn_bits_127;
    end
    if (reset) begin
      _T_926 <= 128'h0;
    end else begin
      _T_926 <= _GEN_128[127:0];
    end
  end
endmodule
module DenseScale(
  input         clock,
  input         reset,
  input         io_dataIn_valid,
  input  [15:0] io_dataIn_bits_0,
  output        io_dataOut_valid,
  output [15:0] io_dataOut_bits_0
);
  reg [6:0] scaleCntr; // @[DenseScale.scala 23:26]
  reg [31:0] _RAND_0;
  wire [15:0] DenseBlackBoxe7682c2e6f_out; // @[DenseScale.scala 28:28]
  wire [6:0] DenseBlackBoxe7682c2e6f_readAddr; // @[DenseScale.scala 28:28]
  wire  DenseBlackBoxe7682c2e6f_clock; // @[DenseScale.scala 28:28]
  wire [15:0] DenseBlackBox4beeeb3293_out; // @[DenseScale.scala 29:28]
  wire [6:0] DenseBlackBox4beeeb3293_readAddr; // @[DenseScale.scala 29:28]
  wire  DenseBlackBox4beeeb3293_clock; // @[DenseScale.scala 29:28]
  reg [15:0] currAct; // @[DenseScale.scala 43:20]
  reg [31:0] _RAND_1;
  reg [15:0] bDelayed; // @[DenseScale.scala 50:25]
  reg [31:0] _RAND_2;
  reg [31:0] scale; // @[DenseScale.scala 52:22]
  reg [31:0] _RAND_3;
  reg [31:0] shift; // @[DenseScale.scala 53:22]
  reg [31:0] _RAND_4;
  reg [15:0] relu; // @[DenseScale.scala 55:17]
  reg [31:0] _RAND_5;
  reg  _T_44; // @[Reg.scala 19:20]
  reg [31:0] _RAND_6;
  reg  _T_46; // @[Reg.scala 19:20]
  reg [31:0] _RAND_7;
  reg  _T_48; // @[Reg.scala 19:20]
  reg [31:0] _RAND_8;
  reg  _T_50; // @[Reg.scala 19:20]
  reg [31:0] _RAND_9;
  wire [7:0] _T_26; // @[DenseScale.scala 25:28]
  wire [6:0] _T_27; // @[DenseScale.scala 25:28]
  wire [6:0] _GEN_0; // @[DenseScale.scala 24:28]
  wire [15:0] currA; // @[DenseScale.scala 47:24]
  wire [15:0] currB; // @[DenseScale.scala 48:24]
  wire [31:0] _T_31; // @[DenseScale.scala 52:32]
  wire [31:0] _GEN_6; // @[DenseScale.scala 53:30]
  wire [32:0] _T_33; // @[DenseScale.scala 53:30]
  wire [31:0] _T_34; // @[DenseScale.scala 53:30]
  wire [31:0] _T_35; // @[DenseScale.scala 53:30]
  wire [31:0] output$; // @[DenseScale.scala 54:22]
  wire  _T_40; // @[DenseScale.scala 57:16]
  wire [31:0] _GEN_1; // @[DenseScale.scala 57:24]
  wire [15:0] _GEN_7;
  DenseBlackBoxe7682c2e6f DenseBlackBoxe7682c2e6f ( // @[DenseScale.scala 28:28]
    .out(DenseBlackBoxe7682c2e6f_out),
    .readAddr(DenseBlackBoxe7682c2e6f_readAddr),
    .clock(DenseBlackBoxe7682c2e6f_clock)
  );
  DenseBlackBox4beeeb3293 DenseBlackBox4beeeb3293 ( // @[DenseScale.scala 29:28]
    .out(DenseBlackBox4beeeb3293_out),
    .readAddr(DenseBlackBox4beeeb3293_readAddr),
    .clock(DenseBlackBox4beeeb3293_clock)
  );
  assign _T_26 = scaleCntr + 7'h1; // @[DenseScale.scala 25:28]
  assign _T_27 = _T_26[6:0]; // @[DenseScale.scala 25:28]
  assign _GEN_0 = io_dataIn_valid ? _T_27 : scaleCntr; // @[DenseScale.scala 24:28]
  assign currA = $signed(DenseBlackBoxe7682c2e6f_out); // @[DenseScale.scala 47:24]
  assign currB = $signed(DenseBlackBox4beeeb3293_out); // @[DenseScale.scala 48:24]
  assign _T_31 = $signed(currAct) * $signed(currA); // @[DenseScale.scala 52:32]
  assign _GEN_6 = {{16{bDelayed[15]}},bDelayed}; // @[DenseScale.scala 53:30]
  assign _T_33 = $signed(scale) + $signed(_GEN_6); // @[DenseScale.scala 53:30]
  assign _T_34 = _T_33[31:0]; // @[DenseScale.scala 53:30]
  assign _T_35 = $signed(_T_34); // @[DenseScale.scala 53:30]
  assign output$ = $signed(shift) >>> 3'h6; // @[DenseScale.scala 54:22]
  assign _T_40 = $signed(shift) > $signed(32'sh0); // @[DenseScale.scala 57:16]
  assign _GEN_1 = _T_40 ? $signed(output$) : $signed(32'sh0); // @[DenseScale.scala 57:24]
  assign io_dataOut_valid = _T_50;
  assign io_dataOut_bits_0 = relu;
  assign DenseBlackBoxe7682c2e6f_readAddr = scaleCntr;
  assign DenseBlackBoxe7682c2e6f_clock = clock;
  assign DenseBlackBox4beeeb3293_readAddr = scaleCntr;
  assign DenseBlackBox4beeeb3293_clock = clock;
  assign _GEN_7 = _GEN_1[15:0];
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  scaleCntr = _RAND_0[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  currAct = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  bDelayed = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  scale = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  shift = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  relu = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  _T_44 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  _T_46 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  _T_48 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  _T_50 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      scaleCntr <= 7'h0;
    end else begin
      if (io_dataIn_valid) begin
        scaleCntr <= _T_27;
      end
    end
    currAct <= io_dataIn_bits_0;
    bDelayed <= currB;
    scale <= _T_31;
    shift <= _T_35;
    relu <= $signed(_GEN_7);
    if (reset) begin
      _T_44 <= 1'h0;
    end else begin
      _T_44 <= io_dataIn_valid;
    end
    if (reset) begin
      _T_46 <= 1'h0;
    end else begin
      _T_46 <= _T_44;
    end
    if (reset) begin
      _T_48 <= 1'h0;
    end else begin
      _T_48 <= _T_46;
    end
    if (reset) begin
      _T_50 <= 1'h0;
    end else begin
      _T_50 <= _T_48;
    end
  end
endmodule
module FanoutAWS_4(
  input         clock,
  input  [15:0] io_in,
  output [15:0] io_out_0,
  output [15:0] io_out_1,
  output [15:0] io_out_2,
  output [15:0] io_out_3,
  output [15:0] io_out_4,
  output [15:0] io_out_5,
  output [15:0] io_out_6,
  output [15:0] io_out_7,
  output [15:0] io_out_8,
  output [15:0] io_out_9
);
  reg [15:0] dataVecs_1_0; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_0;
  reg [15:0] dataVecs_1_1; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_1;
  reg [15:0] dataVecs_2_0; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_2;
  reg [15:0] dataVecs_2_1; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_3;
  reg [15:0] dataVecs_2_2; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_4;
  reg [15:0] dataVecs_2_3; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_5;
  reg [15:0] dataVecs_2_4; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_6;
  reg [15:0] dataVecs_3_0; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_7;
  reg [15:0] dataVecs_3_1; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_8;
  reg [15:0] dataVecs_3_2; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_9;
  reg [15:0] dataVecs_3_3; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_10;
  reg [15:0] dataVecs_3_4; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_11;
  reg [15:0] dataVecs_3_5; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_12;
  reg [15:0] dataVecs_3_6; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_13;
  reg [15:0] dataVecs_3_7; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_14;
  reg [15:0] dataVecs_3_8; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_15;
  reg [15:0] dataVecs_3_9; // @[FanoutAWS.scala 76:31]
  reg [31:0] _RAND_16;
  assign io_out_0 = dataVecs_3_0;
  assign io_out_1 = dataVecs_3_1;
  assign io_out_2 = dataVecs_3_2;
  assign io_out_3 = dataVecs_3_3;
  assign io_out_4 = dataVecs_3_4;
  assign io_out_5 = dataVecs_3_5;
  assign io_out_6 = dataVecs_3_6;
  assign io_out_7 = dataVecs_3_7;
  assign io_out_8 = dataVecs_3_8;
  assign io_out_9 = dataVecs_3_9;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  dataVecs_1_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  dataVecs_1_1 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  dataVecs_2_0 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  dataVecs_2_1 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  dataVecs_2_2 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  dataVecs_2_3 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  dataVecs_2_4 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  dataVecs_3_0 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  dataVecs_3_1 = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  dataVecs_3_2 = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  dataVecs_3_3 = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  dataVecs_3_4 = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  dataVecs_3_5 = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  dataVecs_3_6 = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  dataVecs_3_7 = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  dataVecs_3_8 = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  dataVecs_3_9 = _RAND_16[15:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    dataVecs_1_0 <= io_in;
    dataVecs_1_1 <= io_in;
    dataVecs_2_0 <= dataVecs_1_0;
    dataVecs_2_1 <= dataVecs_1_1;
    dataVecs_2_2 <= dataVecs_1_0;
    dataVecs_2_3 <= dataVecs_1_1;
    dataVecs_2_4 <= dataVecs_1_0;
    dataVecs_3_0 <= dataVecs_2_0;
    dataVecs_3_1 <= dataVecs_2_1;
    dataVecs_3_2 <= dataVecs_2_2;
    dataVecs_3_3 <= dataVecs_2_3;
    dataVecs_3_4 <= dataVecs_2_4;
    dataVecs_3_5 <= dataVecs_2_0;
    dataVecs_3_6 <= dataVecs_2_1;
    dataVecs_3_7 <= dataVecs_2_2;
    dataVecs_3_8 <= dataVecs_2_3;
    dataVecs_3_9 <= dataVecs_2_4;
  end
endmodule
module MultiplyAccumulate_128(
  input         clock,
  input  [15:0] io_activations_0,
  input  [1:0]  io_weights,
  output [15:0] io_sum
);
  reg [15:0] actMult_0; // @[DenseLayer.scala 40:20]
  reg [31:0] _RAND_0;
  wire  _T_11; // @[DenseLayer.scala 48:28]
  wire [15:0] _GEN_0; // @[DenseLayer.scala 48:44]
  wire  _T_14; // @[DenseLayer.scala 52:28]
  wire [16:0] _T_18; // @[DenseLayer.scala 53:31]
  wire [15:0] _T_19; // @[DenseLayer.scala 53:31]
  wire [15:0] _T_20; // @[DenseLayer.scala 53:31]
  wire [15:0] _GEN_1; // @[DenseLayer.scala 52:44]
  assign _T_11 = io_weights[0]; // @[DenseLayer.scala 48:28]
  assign _GEN_0 = _T_11 ? $signed(io_activations_0) : $signed(16'sh0); // @[DenseLayer.scala 48:44]
  assign _T_14 = io_weights[1]; // @[DenseLayer.scala 52:28]
  assign _T_18 = $signed(16'sh0) - $signed(io_activations_0); // @[DenseLayer.scala 53:31]
  assign _T_19 = _T_18[15:0]; // @[DenseLayer.scala 53:31]
  assign _T_20 = $signed(_T_19); // @[DenseLayer.scala 53:31]
  assign _GEN_1 = _T_14 ? $signed(_T_20) : $signed(_GEN_0); // @[DenseLayer.scala 52:44]
  assign io_sum = actMult_0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  actMult_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_14) begin
      actMult_0 <= _T_20;
    end else begin
      if (_T_11) begin
        actMult_0 <= io_activations_0;
      end else begin
        actMult_0 <= 16'sh0;
      end
    end
  end
endmodule
module DenseLayer_1(
  input         clock,
  input         reset,
  input         io_dataIn_valid,
  input  [15:0] io_dataIn_bits_0,
  output        io_dataOut_valid,
  output [15:0] io_dataOut_bits_0,
  output [15:0] io_dataOut_bits_1,
  output [15:0] io_dataOut_bits_2,
  output [15:0] io_dataOut_bits_3,
  output [15:0] io_dataOut_bits_4,
  output [15:0] io_dataOut_bits_5,
  output [15:0] io_dataOut_bits_6,
  output [15:0] io_dataOut_bits_7,
  output [15:0] io_dataOut_bits_8,
  output [15:0] io_dataOut_bits_9
);
  reg [6:0] cntr; // @[DenseLayer.scala 88:21]
  reg [31:0] _RAND_0;
  wire [19:0] weightsRAM_out; // @[DenseLayer.scala 96:34]
  wire [6:0] weightsRAM_readAddr; // @[DenseLayer.scala 96:34]
  wire  weightsRAM_clock; // @[DenseLayer.scala 96:34]
  reg [6:0] _T_51; // @[DenseLayer.scala 97:36]
  reg [31:0] _RAND_1;
  reg [15:0] currActs_0; // @[DenseLayer.scala 102:25]
  reg [31:0] _RAND_2;
  reg [1:0] _T_100_0; // @[Reg.scala 11:16]
  reg [31:0] _RAND_3;
  reg [1:0] _T_100_1; // @[Reg.scala 11:16]
  reg [31:0] _RAND_4;
  reg [1:0] _T_100_2; // @[Reg.scala 11:16]
  reg [31:0] _RAND_5;
  reg [1:0] _T_100_3; // @[Reg.scala 11:16]
  reg [31:0] _RAND_6;
  reg [1:0] _T_100_4; // @[Reg.scala 11:16]
  reg [31:0] _RAND_7;
  reg [1:0] _T_100_5; // @[Reg.scala 11:16]
  reg [31:0] _RAND_8;
  reg [1:0] _T_100_6; // @[Reg.scala 11:16]
  reg [31:0] _RAND_9;
  reg [1:0] _T_100_7; // @[Reg.scala 11:16]
  reg [31:0] _RAND_10;
  reg [1:0] _T_100_8; // @[Reg.scala 11:16]
  reg [31:0] _RAND_11;
  reg [1:0] _T_100_9; // @[Reg.scala 11:16]
  reg [31:0] _RAND_12;
  reg [1:0] delayWeights_0; // @[Reg.scala 11:16]
  reg [31:0] _RAND_13;
  reg [1:0] delayWeights_1; // @[Reg.scala 11:16]
  reg [31:0] _RAND_14;
  reg [1:0] delayWeights_2; // @[Reg.scala 11:16]
  reg [31:0] _RAND_15;
  reg [1:0] delayWeights_3; // @[Reg.scala 11:16]
  reg [31:0] _RAND_16;
  reg [1:0] delayWeights_4; // @[Reg.scala 11:16]
  reg [31:0] _RAND_17;
  reg [1:0] delayWeights_5; // @[Reg.scala 11:16]
  reg [31:0] _RAND_18;
  reg [1:0] delayWeights_6; // @[Reg.scala 11:16]
  reg [31:0] _RAND_19;
  reg [1:0] delayWeights_7; // @[Reg.scala 11:16]
  reg [31:0] _RAND_20;
  reg [1:0] delayWeights_8; // @[Reg.scala 11:16]
  reg [31:0] _RAND_21;
  reg [1:0] delayWeights_9; // @[Reg.scala 11:16]
  reg [31:0] _RAND_22;
  wire  FanoutAWS_clock; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_in; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_0; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_1; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_2; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_3; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_4; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_5; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_6; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_7; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_8; // @[FanoutAWS.scala 16:26]
  wire [15:0] FanoutAWS_io_out_9; // @[FanoutAWS.scala 16:26]
  wire  MultiplyAccumulate_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [1:0] MultiplyAccumulate_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_1_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_1_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [1:0] MultiplyAccumulate_1_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_1_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_2_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_2_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [1:0] MultiplyAccumulate_2_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_2_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_3_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_3_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [1:0] MultiplyAccumulate_3_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_3_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_4_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_4_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [1:0] MultiplyAccumulate_4_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_4_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_5_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_5_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [1:0] MultiplyAccumulate_5_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_5_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_6_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_6_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [1:0] MultiplyAccumulate_6_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_6_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_7_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_7_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [1:0] MultiplyAccumulate_7_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_7_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_8_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_8_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [1:0] MultiplyAccumulate_8_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_8_io_sum; // @[DenseLayer.scala 111:21]
  wire  MultiplyAccumulate_9_clock; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_9_io_activations_0; // @[DenseLayer.scala 111:21]
  wire [1:0] MultiplyAccumulate_9_io_weights; // @[DenseLayer.scala 111:21]
  wire [15:0] MultiplyAccumulate_9_io_sum; // @[DenseLayer.scala 111:21]
  reg [15:0] cummulativeSums_0; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_23;
  reg [15:0] cummulativeSums_1; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_24;
  reg [15:0] cummulativeSums_2; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_25;
  reg [15:0] cummulativeSums_3; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_26;
  reg [15:0] cummulativeSums_4; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_27;
  reg [15:0] cummulativeSums_5; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_28;
  reg [15:0] cummulativeSums_6; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_29;
  reg [15:0] cummulativeSums_7; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_30;
  reg [15:0] cummulativeSums_8; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_31;
  reg [15:0] cummulativeSums_9; // @[DenseLayer.scala 120:28]
  reg [31:0] _RAND_32;
  reg  _T_256; // @[Reg.scala 11:16]
  reg [31:0] _RAND_33;
  reg  _T_258; // @[Reg.scala 11:16]
  reg [31:0] _RAND_34;
  reg  _T_260; // @[Reg.scala 11:16]
  reg [31:0] _RAND_35;
  reg  _T_262; // @[Reg.scala 11:16]
  reg [31:0] _RAND_36;
  reg  rst; // @[Reg.scala 11:16]
  reg [31:0] _RAND_37;
  reg  done; // @[DenseLayer.scala 122:21]
  reg [31:0] _RAND_38;
  reg  _T_273; // @[Reg.scala 11:16]
  reg [31:0] _RAND_39;
  reg  _T_275; // @[Reg.scala 11:16]
  reg [31:0] _RAND_40;
  reg  _T_277; // @[Reg.scala 11:16]
  reg [31:0] _RAND_41;
  reg  _T_279; // @[Reg.scala 11:16]
  reg [31:0] _RAND_42;
  reg  vld; // @[Reg.scala 11:16]
  reg [31:0] _RAND_43;
  wire [7:0] _T_34; // @[DenseLayer.scala 90:18]
  wire [6:0] _T_35; // @[DenseLayer.scala 90:18]
  wire [6:0] _GEN_0; // @[DenseLayer.scala 89:28]
  wire [1:0] currWeights_0; // @[DenseLayer.scala 100:42]
  wire [1:0] currWeights_1; // @[DenseLayer.scala 100:42]
  wire [1:0] currWeights_2; // @[DenseLayer.scala 100:42]
  wire [1:0] currWeights_3; // @[DenseLayer.scala 100:42]
  wire [1:0] currWeights_4; // @[DenseLayer.scala 100:42]
  wire [1:0] currWeights_5; // @[DenseLayer.scala 100:42]
  wire [1:0] currWeights_6; // @[DenseLayer.scala 100:42]
  wire [1:0] currWeights_7; // @[DenseLayer.scala 100:42]
  wire [1:0] currWeights_8; // @[DenseLayer.scala 100:42]
  wire [1:0] currWeights_9; // @[DenseLayer.scala 100:42]
  wire  _T_253; // @[DenseLayer.scala 121:33]
  wire  _T_267; // @[DenseLayer.scala 123:16]
  wire  _GEN_26; // @[DenseLayer.scala 123:42]
  wire  _T_269; // @[DenseLayer.scala 126:14]
  wire  _GEN_27; // @[DenseLayer.scala 126:23]
  wire [16:0] _T_281; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_282; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_283; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_33; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_34; // @[DenseLayer.scala 135:18]
  wire  _T_285; // @[DenseLayer.scala 138:16]
  wire [15:0] _GEN_35; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_286; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_287; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_288; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_36; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_37; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_38; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_291; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_292; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_293; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_39; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_40; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_41; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_296; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_297; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_298; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_42; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_43; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_44; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_301; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_302; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_303; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_45; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_46; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_47; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_306; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_307; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_308; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_48; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_49; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_50; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_311; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_312; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_313; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_51; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_52; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_53; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_316; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_317; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_318; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_54; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_55; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_56; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_321; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_322; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_323; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_57; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_58; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_59; // @[DenseLayer.scala 138:24]
  wire [16:0] _T_326; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_327; // @[DenseLayer.scala 133:59]
  wire [15:0] _T_328; // @[DenseLayer.scala 133:59]
  wire [15:0] _GEN_60; // @[DenseLayer.scala 132:18]
  wire [15:0] _GEN_61; // @[DenseLayer.scala 135:18]
  wire [15:0] _GEN_62; // @[DenseLayer.scala 138:24]
  DenseBlackBox255c5dd06e weightsRAM ( // @[DenseLayer.scala 96:34]
    .out(weightsRAM_out),
    .readAddr(weightsRAM_readAddr),
    .clock(weightsRAM_clock)
  );
  FanoutAWS_4 FanoutAWS ( // @[FanoutAWS.scala 16:26]
    .clock(FanoutAWS_clock),
    .io_in(FanoutAWS_io_in),
    .io_out_0(FanoutAWS_io_out_0),
    .io_out_1(FanoutAWS_io_out_1),
    .io_out_2(FanoutAWS_io_out_2),
    .io_out_3(FanoutAWS_io_out_3),
    .io_out_4(FanoutAWS_io_out_4),
    .io_out_5(FanoutAWS_io_out_5),
    .io_out_6(FanoutAWS_io_out_6),
    .io_out_7(FanoutAWS_io_out_7),
    .io_out_8(FanoutAWS_io_out_8),
    .io_out_9(FanoutAWS_io_out_9)
  );
  MultiplyAccumulate_128 MultiplyAccumulate ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_clock),
    .io_activations_0(MultiplyAccumulate_io_activations_0),
    .io_weights(MultiplyAccumulate_io_weights),
    .io_sum(MultiplyAccumulate_io_sum)
  );
  MultiplyAccumulate_128 MultiplyAccumulate_1 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_1_clock),
    .io_activations_0(MultiplyAccumulate_1_io_activations_0),
    .io_weights(MultiplyAccumulate_1_io_weights),
    .io_sum(MultiplyAccumulate_1_io_sum)
  );
  MultiplyAccumulate_128 MultiplyAccumulate_2 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_2_clock),
    .io_activations_0(MultiplyAccumulate_2_io_activations_0),
    .io_weights(MultiplyAccumulate_2_io_weights),
    .io_sum(MultiplyAccumulate_2_io_sum)
  );
  MultiplyAccumulate_128 MultiplyAccumulate_3 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_3_clock),
    .io_activations_0(MultiplyAccumulate_3_io_activations_0),
    .io_weights(MultiplyAccumulate_3_io_weights),
    .io_sum(MultiplyAccumulate_3_io_sum)
  );
  MultiplyAccumulate_128 MultiplyAccumulate_4 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_4_clock),
    .io_activations_0(MultiplyAccumulate_4_io_activations_0),
    .io_weights(MultiplyAccumulate_4_io_weights),
    .io_sum(MultiplyAccumulate_4_io_sum)
  );
  MultiplyAccumulate_128 MultiplyAccumulate_5 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_5_clock),
    .io_activations_0(MultiplyAccumulate_5_io_activations_0),
    .io_weights(MultiplyAccumulate_5_io_weights),
    .io_sum(MultiplyAccumulate_5_io_sum)
  );
  MultiplyAccumulate_128 MultiplyAccumulate_6 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_6_clock),
    .io_activations_0(MultiplyAccumulate_6_io_activations_0),
    .io_weights(MultiplyAccumulate_6_io_weights),
    .io_sum(MultiplyAccumulate_6_io_sum)
  );
  MultiplyAccumulate_128 MultiplyAccumulate_7 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_7_clock),
    .io_activations_0(MultiplyAccumulate_7_io_activations_0),
    .io_weights(MultiplyAccumulate_7_io_weights),
    .io_sum(MultiplyAccumulate_7_io_sum)
  );
  MultiplyAccumulate_128 MultiplyAccumulate_8 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_8_clock),
    .io_activations_0(MultiplyAccumulate_8_io_activations_0),
    .io_weights(MultiplyAccumulate_8_io_weights),
    .io_sum(MultiplyAccumulate_8_io_sum)
  );
  MultiplyAccumulate_128 MultiplyAccumulate_9 ( // @[DenseLayer.scala 111:21]
    .clock(MultiplyAccumulate_9_clock),
    .io_activations_0(MultiplyAccumulate_9_io_activations_0),
    .io_weights(MultiplyAccumulate_9_io_weights),
    .io_sum(MultiplyAccumulate_9_io_sum)
  );
  assign _T_34 = cntr + 7'h1; // @[DenseLayer.scala 90:18]
  assign _T_35 = _T_34[6:0]; // @[DenseLayer.scala 90:18]
  assign _GEN_0 = io_dataIn_valid ? _T_35 : cntr; // @[DenseLayer.scala 89:28]
  assign currWeights_0 = weightsRAM_out[1:0]; // @[DenseLayer.scala 100:42]
  assign currWeights_1 = weightsRAM_out[3:2]; // @[DenseLayer.scala 100:42]
  assign currWeights_2 = weightsRAM_out[5:4]; // @[DenseLayer.scala 100:42]
  assign currWeights_3 = weightsRAM_out[7:6]; // @[DenseLayer.scala 100:42]
  assign currWeights_4 = weightsRAM_out[9:8]; // @[DenseLayer.scala 100:42]
  assign currWeights_5 = weightsRAM_out[11:10]; // @[DenseLayer.scala 100:42]
  assign currWeights_6 = weightsRAM_out[13:12]; // @[DenseLayer.scala 100:42]
  assign currWeights_7 = weightsRAM_out[15:14]; // @[DenseLayer.scala 100:42]
  assign currWeights_8 = weightsRAM_out[17:16]; // @[DenseLayer.scala 100:42]
  assign currWeights_9 = weightsRAM_out[19:18]; // @[DenseLayer.scala 100:42]
  assign _T_253 = cntr == 7'h0; // @[DenseLayer.scala 121:33]
  assign _T_267 = cntr == 7'h7f; // @[DenseLayer.scala 123:16]
  assign _GEN_26 = _T_267 ? 1'h1 : done; // @[DenseLayer.scala 123:42]
  assign _T_269 = rst & done; // @[DenseLayer.scala 126:14]
  assign _GEN_27 = _T_269 ? 1'h0 : _GEN_26; // @[DenseLayer.scala 126:23]
  assign _T_281 = $signed(cummulativeSums_0) + $signed(MultiplyAccumulate_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_282 = _T_281[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_283 = $signed(_T_282); // @[DenseLayer.scala 133:59]
  assign _GEN_33 = vld ? $signed(_T_283) : $signed(cummulativeSums_0); // @[DenseLayer.scala 132:18]
  assign _GEN_34 = rst ? $signed(16'sh0) : $signed(_GEN_33); // @[DenseLayer.scala 135:18]
  assign _T_285 = rst & vld; // @[DenseLayer.scala 138:16]
  assign _GEN_35 = _T_285 ? $signed(MultiplyAccumulate_io_sum) : $signed(_GEN_34); // @[DenseLayer.scala 138:24]
  assign _T_286 = $signed(cummulativeSums_1) + $signed(MultiplyAccumulate_1_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_287 = _T_286[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_288 = $signed(_T_287); // @[DenseLayer.scala 133:59]
  assign _GEN_36 = vld ? $signed(_T_288) : $signed(cummulativeSums_1); // @[DenseLayer.scala 132:18]
  assign _GEN_37 = rst ? $signed(16'sh0) : $signed(_GEN_36); // @[DenseLayer.scala 135:18]
  assign _GEN_38 = _T_285 ? $signed(MultiplyAccumulate_1_io_sum) : $signed(_GEN_37); // @[DenseLayer.scala 138:24]
  assign _T_291 = $signed(cummulativeSums_2) + $signed(MultiplyAccumulate_2_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_292 = _T_291[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_293 = $signed(_T_292); // @[DenseLayer.scala 133:59]
  assign _GEN_39 = vld ? $signed(_T_293) : $signed(cummulativeSums_2); // @[DenseLayer.scala 132:18]
  assign _GEN_40 = rst ? $signed(16'sh0) : $signed(_GEN_39); // @[DenseLayer.scala 135:18]
  assign _GEN_41 = _T_285 ? $signed(MultiplyAccumulate_2_io_sum) : $signed(_GEN_40); // @[DenseLayer.scala 138:24]
  assign _T_296 = $signed(cummulativeSums_3) + $signed(MultiplyAccumulate_3_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_297 = _T_296[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_298 = $signed(_T_297); // @[DenseLayer.scala 133:59]
  assign _GEN_42 = vld ? $signed(_T_298) : $signed(cummulativeSums_3); // @[DenseLayer.scala 132:18]
  assign _GEN_43 = rst ? $signed(16'sh0) : $signed(_GEN_42); // @[DenseLayer.scala 135:18]
  assign _GEN_44 = _T_285 ? $signed(MultiplyAccumulate_3_io_sum) : $signed(_GEN_43); // @[DenseLayer.scala 138:24]
  assign _T_301 = $signed(cummulativeSums_4) + $signed(MultiplyAccumulate_4_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_302 = _T_301[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_303 = $signed(_T_302); // @[DenseLayer.scala 133:59]
  assign _GEN_45 = vld ? $signed(_T_303) : $signed(cummulativeSums_4); // @[DenseLayer.scala 132:18]
  assign _GEN_46 = rst ? $signed(16'sh0) : $signed(_GEN_45); // @[DenseLayer.scala 135:18]
  assign _GEN_47 = _T_285 ? $signed(MultiplyAccumulate_4_io_sum) : $signed(_GEN_46); // @[DenseLayer.scala 138:24]
  assign _T_306 = $signed(cummulativeSums_5) + $signed(MultiplyAccumulate_5_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_307 = _T_306[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_308 = $signed(_T_307); // @[DenseLayer.scala 133:59]
  assign _GEN_48 = vld ? $signed(_T_308) : $signed(cummulativeSums_5); // @[DenseLayer.scala 132:18]
  assign _GEN_49 = rst ? $signed(16'sh0) : $signed(_GEN_48); // @[DenseLayer.scala 135:18]
  assign _GEN_50 = _T_285 ? $signed(MultiplyAccumulate_5_io_sum) : $signed(_GEN_49); // @[DenseLayer.scala 138:24]
  assign _T_311 = $signed(cummulativeSums_6) + $signed(MultiplyAccumulate_6_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_312 = _T_311[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_313 = $signed(_T_312); // @[DenseLayer.scala 133:59]
  assign _GEN_51 = vld ? $signed(_T_313) : $signed(cummulativeSums_6); // @[DenseLayer.scala 132:18]
  assign _GEN_52 = rst ? $signed(16'sh0) : $signed(_GEN_51); // @[DenseLayer.scala 135:18]
  assign _GEN_53 = _T_285 ? $signed(MultiplyAccumulate_6_io_sum) : $signed(_GEN_52); // @[DenseLayer.scala 138:24]
  assign _T_316 = $signed(cummulativeSums_7) + $signed(MultiplyAccumulate_7_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_317 = _T_316[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_318 = $signed(_T_317); // @[DenseLayer.scala 133:59]
  assign _GEN_54 = vld ? $signed(_T_318) : $signed(cummulativeSums_7); // @[DenseLayer.scala 132:18]
  assign _GEN_55 = rst ? $signed(16'sh0) : $signed(_GEN_54); // @[DenseLayer.scala 135:18]
  assign _GEN_56 = _T_285 ? $signed(MultiplyAccumulate_7_io_sum) : $signed(_GEN_55); // @[DenseLayer.scala 138:24]
  assign _T_321 = $signed(cummulativeSums_8) + $signed(MultiplyAccumulate_8_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_322 = _T_321[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_323 = $signed(_T_322); // @[DenseLayer.scala 133:59]
  assign _GEN_57 = vld ? $signed(_T_323) : $signed(cummulativeSums_8); // @[DenseLayer.scala 132:18]
  assign _GEN_58 = rst ? $signed(16'sh0) : $signed(_GEN_57); // @[DenseLayer.scala 135:18]
  assign _GEN_59 = _T_285 ? $signed(MultiplyAccumulate_8_io_sum) : $signed(_GEN_58); // @[DenseLayer.scala 138:24]
  assign _T_326 = $signed(cummulativeSums_9) + $signed(MultiplyAccumulate_9_io_sum); // @[DenseLayer.scala 133:59]
  assign _T_327 = _T_326[15:0]; // @[DenseLayer.scala 133:59]
  assign _T_328 = $signed(_T_327); // @[DenseLayer.scala 133:59]
  assign _GEN_60 = vld ? $signed(_T_328) : $signed(cummulativeSums_9); // @[DenseLayer.scala 132:18]
  assign _GEN_61 = rst ? $signed(16'sh0) : $signed(_GEN_60); // @[DenseLayer.scala 135:18]
  assign _GEN_62 = _T_285 ? $signed(MultiplyAccumulate_9_io_sum) : $signed(_GEN_61); // @[DenseLayer.scala 138:24]
  assign io_dataOut_valid = _T_269;
  assign io_dataOut_bits_0 = cummulativeSums_0;
  assign io_dataOut_bits_1 = cummulativeSums_1;
  assign io_dataOut_bits_2 = cummulativeSums_2;
  assign io_dataOut_bits_3 = cummulativeSums_3;
  assign io_dataOut_bits_4 = cummulativeSums_4;
  assign io_dataOut_bits_5 = cummulativeSums_5;
  assign io_dataOut_bits_6 = cummulativeSums_6;
  assign io_dataOut_bits_7 = cummulativeSums_7;
  assign io_dataOut_bits_8 = cummulativeSums_8;
  assign io_dataOut_bits_9 = cummulativeSums_9;
  assign weightsRAM_readAddr = _T_51;
  assign weightsRAM_clock = clock;
  assign FanoutAWS_clock = clock;
  assign FanoutAWS_io_in = currActs_0;
  assign MultiplyAccumulate_clock = clock;
  assign MultiplyAccumulate_io_activations_0 = FanoutAWS_io_out_0;
  assign MultiplyAccumulate_io_weights = delayWeights_0;
  assign MultiplyAccumulate_1_clock = clock;
  assign MultiplyAccumulate_1_io_activations_0 = FanoutAWS_io_out_1;
  assign MultiplyAccumulate_1_io_weights = delayWeights_1;
  assign MultiplyAccumulate_2_clock = clock;
  assign MultiplyAccumulate_2_io_activations_0 = FanoutAWS_io_out_2;
  assign MultiplyAccumulate_2_io_weights = delayWeights_2;
  assign MultiplyAccumulate_3_clock = clock;
  assign MultiplyAccumulate_3_io_activations_0 = FanoutAWS_io_out_3;
  assign MultiplyAccumulate_3_io_weights = delayWeights_3;
  assign MultiplyAccumulate_4_clock = clock;
  assign MultiplyAccumulate_4_io_activations_0 = FanoutAWS_io_out_4;
  assign MultiplyAccumulate_4_io_weights = delayWeights_4;
  assign MultiplyAccumulate_5_clock = clock;
  assign MultiplyAccumulate_5_io_activations_0 = FanoutAWS_io_out_5;
  assign MultiplyAccumulate_5_io_weights = delayWeights_5;
  assign MultiplyAccumulate_6_clock = clock;
  assign MultiplyAccumulate_6_io_activations_0 = FanoutAWS_io_out_6;
  assign MultiplyAccumulate_6_io_weights = delayWeights_6;
  assign MultiplyAccumulate_7_clock = clock;
  assign MultiplyAccumulate_7_io_activations_0 = FanoutAWS_io_out_7;
  assign MultiplyAccumulate_7_io_weights = delayWeights_7;
  assign MultiplyAccumulate_8_clock = clock;
  assign MultiplyAccumulate_8_io_activations_0 = FanoutAWS_io_out_8;
  assign MultiplyAccumulate_8_io_weights = delayWeights_8;
  assign MultiplyAccumulate_9_clock = clock;
  assign MultiplyAccumulate_9_io_activations_0 = FanoutAWS_io_out_9;
  assign MultiplyAccumulate_9_io_weights = delayWeights_9;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  cntr = _RAND_0[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  _T_51 = _RAND_1[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  currActs_0 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_100_0 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  _T_100_1 = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  _T_100_2 = _RAND_5[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  _T_100_3 = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  _T_100_4 = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  _T_100_5 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  _T_100_6 = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  _T_100_7 = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  _T_100_8 = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  _T_100_9 = _RAND_12[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  delayWeights_0 = _RAND_13[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  delayWeights_1 = _RAND_14[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  delayWeights_2 = _RAND_15[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  delayWeights_3 = _RAND_16[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  delayWeights_4 = _RAND_17[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  delayWeights_5 = _RAND_18[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  delayWeights_6 = _RAND_19[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  delayWeights_7 = _RAND_20[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  delayWeights_8 = _RAND_21[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  delayWeights_9 = _RAND_22[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  cummulativeSums_0 = _RAND_23[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  cummulativeSums_1 = _RAND_24[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  cummulativeSums_2 = _RAND_25[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  cummulativeSums_3 = _RAND_26[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  cummulativeSums_4 = _RAND_27[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  cummulativeSums_5 = _RAND_28[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  cummulativeSums_6 = _RAND_29[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  cummulativeSums_7 = _RAND_30[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  cummulativeSums_8 = _RAND_31[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  cummulativeSums_9 = _RAND_32[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{$random}};
  _T_256 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{$random}};
  _T_258 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{$random}};
  _T_260 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{$random}};
  _T_262 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{$random}};
  rst = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{$random}};
  done = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{$random}};
  _T_273 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{$random}};
  _T_275 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{$random}};
  _T_277 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{$random}};
  _T_279 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{$random}};
  vld = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cntr <= 7'h0;
    end else begin
      if (io_dataIn_valid) begin
        cntr <= _T_35;
      end
    end
    _T_51 <= cntr;
    currActs_0 <= io_dataIn_bits_0;
    _T_100_0 <= currWeights_0;
    _T_100_1 <= currWeights_1;
    _T_100_2 <= currWeights_2;
    _T_100_3 <= currWeights_3;
    _T_100_4 <= currWeights_4;
    _T_100_5 <= currWeights_5;
    _T_100_6 <= currWeights_6;
    _T_100_7 <= currWeights_7;
    _T_100_8 <= currWeights_8;
    _T_100_9 <= currWeights_9;
    delayWeights_0 <= _T_100_0;
    delayWeights_1 <= _T_100_1;
    delayWeights_2 <= _T_100_2;
    delayWeights_3 <= _T_100_3;
    delayWeights_4 <= _T_100_4;
    delayWeights_5 <= _T_100_5;
    delayWeights_6 <= _T_100_6;
    delayWeights_7 <= _T_100_7;
    delayWeights_8 <= _T_100_8;
    delayWeights_9 <= _T_100_9;
    if (_T_285) begin
      cummulativeSums_0 <= MultiplyAccumulate_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_0 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_0 <= _T_283;
        end
      end
    end
    if (_T_285) begin
      cummulativeSums_1 <= MultiplyAccumulate_1_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_1 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_1 <= _T_288;
        end
      end
    end
    if (_T_285) begin
      cummulativeSums_2 <= MultiplyAccumulate_2_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_2 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_2 <= _T_293;
        end
      end
    end
    if (_T_285) begin
      cummulativeSums_3 <= MultiplyAccumulate_3_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_3 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_3 <= _T_298;
        end
      end
    end
    if (_T_285) begin
      cummulativeSums_4 <= MultiplyAccumulate_4_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_4 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_4 <= _T_303;
        end
      end
    end
    if (_T_285) begin
      cummulativeSums_5 <= MultiplyAccumulate_5_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_5 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_5 <= _T_308;
        end
      end
    end
    if (_T_285) begin
      cummulativeSums_6 <= MultiplyAccumulate_6_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_6 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_6 <= _T_313;
        end
      end
    end
    if (_T_285) begin
      cummulativeSums_7 <= MultiplyAccumulate_7_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_7 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_7 <= _T_318;
        end
      end
    end
    if (_T_285) begin
      cummulativeSums_8 <= MultiplyAccumulate_8_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_8 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_8 <= _T_323;
        end
      end
    end
    if (_T_285) begin
      cummulativeSums_9 <= MultiplyAccumulate_9_io_sum;
    end else begin
      if (rst) begin
        cummulativeSums_9 <= 16'sh0;
      end else begin
        if (vld) begin
          cummulativeSums_9 <= _T_328;
        end
      end
    end
    _T_256 <= _T_253;
    _T_258 <= _T_256;
    _T_260 <= _T_258;
    _T_262 <= _T_260;
    rst <= _T_262;
    if (reset) begin
      done <= 1'h0;
    end else begin
      if (_T_269) begin
        done <= 1'h0;
      end else begin
        if (_T_267) begin
          done <= 1'h1;
        end
      end
    end
    _T_273 <= io_dataIn_valid;
    _T_275 <= _T_273;
    _T_277 <= _T_275;
    _T_279 <= _T_277;
    vld <= _T_279;
  end
endmodule
module AWSVggWrapper(
  input         clock,
  input         reset,
  output        io_dataIn_ready,
  input         io_dataIn_valid,
  input  [15:0] io_dataIn_bits_0,
  input  [15:0] io_dataIn_bits_1,
  input  [15:0] io_dataIn_bits_2,
  input         io_dataOut_ready,
  output        io_dataOut_valid,
  output [15:0] io_dataOut_bits_0,
  output [15:0] io_dataOut_bits_1,
  output [15:0] io_dataOut_bits_2,
  output [15:0] io_dataOut_bits_3,
  output [15:0] io_dataOut_bits_4,
  output [15:0] io_dataOut_bits_5,
  output [15:0] io_dataOut_bits_6,
  output [15:0] io_dataOut_bits_7,
  output [15:0] io_dataOut_bits_8,
  output [15:0] io_dataOut_bits_9
);
  wire  vgg_clock; // @[AWSVggWrapper.scala 47:27]
  wire  vgg_reset; // @[AWSVggWrapper.scala 47:27]
  wire  vgg_io_dataIn_ready; // @[AWSVggWrapper.scala 47:27]
  wire  vgg_io_dataIn_valid; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataIn_bits_0; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataIn_bits_1; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataIn_bits_2; // @[AWSVggWrapper.scala 47:27]
  wire  vgg_io_dataOut_ready; // @[AWSVggWrapper.scala 47:27]
  wire  vgg_io_dataOut_valid; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_0; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_1; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_2; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_3; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_4; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_5; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_6; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_7; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_8; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_9; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_10; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_11; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_12; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_13; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_14; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_15; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_16; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_17; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_18; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_19; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_20; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_21; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_22; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_23; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_24; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_25; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_26; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_27; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_28; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_29; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_30; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_31; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_32; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_33; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_34; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_35; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_36; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_37; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_38; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_39; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_40; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_41; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_42; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_43; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_44; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_45; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_46; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_47; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_48; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_49; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_50; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_51; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_52; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_53; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_54; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_55; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_56; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_57; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_58; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_59; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_60; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_61; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_62; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_63; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_64; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_65; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_66; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_67; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_68; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_69; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_70; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_71; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_72; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_73; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_74; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_75; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_76; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_77; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_78; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_79; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_80; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_81; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_82; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_83; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_84; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_85; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_86; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_87; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_88; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_89; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_90; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_91; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_92; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_93; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_94; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_95; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_96; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_97; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_98; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_99; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_100; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_101; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_102; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_103; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_104; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_105; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_106; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_107; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_108; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_109; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_110; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_111; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_112; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_113; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_114; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_115; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_116; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_117; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_118; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_119; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_120; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_121; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_122; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_123; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_124; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_125; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_126; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_127; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_128; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_129; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_130; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_131; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_132; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_133; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_134; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_135; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_136; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_137; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_138; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_139; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_140; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_141; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_142; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_143; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_144; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_145; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_146; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_147; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_148; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_149; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_150; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_151; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_152; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_153; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_154; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_155; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_156; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_157; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_158; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_159; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_160; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_161; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_162; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_163; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_164; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_165; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_166; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_167; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_168; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_169; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_170; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_171; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_172; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_173; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_174; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_175; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_176; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_177; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_178; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_179; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_180; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_181; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_182; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_183; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_184; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_185; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_186; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_187; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_188; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_189; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_190; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_191; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_192; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_193; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_194; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_195; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_196; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_197; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_198; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_199; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_200; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_201; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_202; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_203; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_204; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_205; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_206; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_207; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_208; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_209; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_210; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_211; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_212; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_213; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_214; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_215; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_216; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_217; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_218; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_219; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_220; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_221; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_222; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_223; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_224; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_225; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_226; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_227; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_228; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_229; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_230; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_231; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_232; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_233; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_234; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_235; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_236; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_237; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_238; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_239; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_240; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_241; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_242; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_243; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_244; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_245; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_246; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_247; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_248; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_249; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_250; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_251; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_252; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_253; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_254; // @[AWSVggWrapper.scala 47:27]
  wire [15:0] vgg_io_dataOut_bits_255; // @[AWSVggWrapper.scala 47:27]
  wire  queueIOOut_clock; // @[Decoupled.scala 289:19]
  wire  queueIOOut_reset; // @[Decoupled.scala 289:19]
  wire  queueIOOut_io_enq_ready; // @[Decoupled.scala 289:19]
  wire  queueIOOut_io_enq_valid; // @[Decoupled.scala 289:19]
  wire [4095:0] queueIOOut_io_enq_bits; // @[Decoupled.scala 289:19]
  wire  queueIOOut_io_deq_ready; // @[Decoupled.scala 289:19]
  wire  queueIOOut_io_deq_valid; // @[Decoupled.scala 289:19]
  wire [4095:0] queueIOOut_io_deq_bits; // @[Decoupled.scala 289:19]
  wire  muxLyr_clock; // @[AWSVggWrapper.scala 66:22]
  wire  muxLyr_reset; // @[AWSVggWrapper.scala 66:22]
  wire  muxLyr_io_dataIn_ready; // @[AWSVggWrapper.scala 66:22]
  wire  muxLyr_io_dataIn_valid; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_0; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_1; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_2; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_3; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_4; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_5; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_6; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_7; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_8; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_9; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_10; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_11; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_12; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_13; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_14; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_15; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_16; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_17; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_18; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_19; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_20; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_21; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_22; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_23; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_24; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_25; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_26; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_27; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_28; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_29; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_30; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_31; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_32; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_33; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_34; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_35; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_36; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_37; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_38; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_39; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_40; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_41; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_42; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_43; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_44; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_45; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_46; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_47; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_48; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_49; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_50; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_51; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_52; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_53; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_54; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_55; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_56; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_57; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_58; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_59; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_60; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_61; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_62; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_63; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_64; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_65; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_66; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_67; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_68; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_69; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_70; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_71; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_72; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_73; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_74; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_75; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_76; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_77; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_78; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_79; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_80; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_81; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_82; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_83; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_84; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_85; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_86; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_87; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_88; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_89; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_90; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_91; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_92; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_93; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_94; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_95; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_96; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_97; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_98; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_99; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_100; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_101; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_102; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_103; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_104; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_105; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_106; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_107; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_108; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_109; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_110; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_111; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_112; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_113; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_114; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_115; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_116; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_117; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_118; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_119; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_120; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_121; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_122; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_123; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_124; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_125; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_126; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_127; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_128; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_129; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_130; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_131; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_132; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_133; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_134; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_135; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_136; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_137; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_138; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_139; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_140; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_141; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_142; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_143; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_144; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_145; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_146; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_147; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_148; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_149; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_150; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_151; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_152; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_153; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_154; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_155; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_156; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_157; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_158; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_159; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_160; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_161; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_162; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_163; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_164; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_165; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_166; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_167; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_168; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_169; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_170; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_171; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_172; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_173; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_174; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_175; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_176; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_177; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_178; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_179; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_180; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_181; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_182; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_183; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_184; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_185; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_186; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_187; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_188; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_189; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_190; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_191; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_192; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_193; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_194; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_195; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_196; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_197; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_198; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_199; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_200; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_201; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_202; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_203; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_204; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_205; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_206; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_207; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_208; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_209; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_210; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_211; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_212; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_213; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_214; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_215; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_216; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_217; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_218; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_219; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_220; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_221; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_222; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_223; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_224; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_225; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_226; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_227; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_228; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_229; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_230; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_231; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_232; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_233; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_234; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_235; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_236; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_237; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_238; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_239; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_240; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_241; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_242; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_243; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_244; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_245; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_246; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_247; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_248; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_249; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_250; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_251; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_252; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_253; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_254; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataIn_bits_255; // @[AWSVggWrapper.scala 66:22]
  wire  muxLyr_io_dataOut_valid; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataOut_bits_0; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataOut_bits_1; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataOut_bits_2; // @[AWSVggWrapper.scala 66:22]
  wire [15:0] muxLyr_io_dataOut_bits_3; // @[AWSVggWrapper.scala 66:22]
  wire  dense_clock; // @[AWSVggWrapper.scala 75:21]
  wire  dense_reset; // @[AWSVggWrapper.scala 75:21]
  wire  dense_io_dataIn_valid; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataIn_bits_0; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataIn_bits_1; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataIn_bits_2; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataIn_bits_3; // @[AWSVggWrapper.scala 75:21]
  wire  dense_io_dataOut_valid; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_0; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_1; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_2; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_3; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_4; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_5; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_6; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_7; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_8; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_9; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_10; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_11; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_12; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_13; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_14; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_15; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_16; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_17; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_18; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_19; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_20; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_21; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_22; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_23; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_24; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_25; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_26; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_27; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_28; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_29; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_30; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_31; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_32; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_33; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_34; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_35; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_36; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_37; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_38; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_39; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_40; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_41; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_42; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_43; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_44; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_45; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_46; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_47; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_48; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_49; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_50; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_51; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_52; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_53; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_54; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_55; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_56; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_57; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_58; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_59; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_60; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_61; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_62; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_63; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_64; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_65; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_66; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_67; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_68; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_69; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_70; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_71; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_72; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_73; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_74; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_75; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_76; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_77; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_78; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_79; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_80; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_81; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_82; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_83; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_84; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_85; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_86; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_87; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_88; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_89; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_90; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_91; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_92; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_93; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_94; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_95; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_96; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_97; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_98; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_99; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_100; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_101; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_102; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_103; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_104; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_105; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_106; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_107; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_108; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_109; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_110; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_111; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_112; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_113; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_114; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_115; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_116; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_117; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_118; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_119; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_120; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_121; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_122; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_123; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_124; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_125; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_126; // @[AWSVggWrapper.scala 75:21]
  wire [15:0] dense_io_dataOut_bits_127; // @[AWSVggWrapper.scala 75:21]
  wire  muxLyr_2_clock; // @[AWSVggWrapper.scala 79:24]
  wire  muxLyr_2_reset; // @[AWSVggWrapper.scala 79:24]
  wire  muxLyr_2_io_dataIn_valid; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_0; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_1; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_2; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_3; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_4; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_5; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_6; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_7; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_8; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_9; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_10; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_11; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_12; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_13; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_14; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_15; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_16; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_17; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_18; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_19; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_20; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_21; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_22; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_23; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_24; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_25; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_26; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_27; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_28; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_29; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_30; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_31; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_32; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_33; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_34; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_35; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_36; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_37; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_38; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_39; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_40; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_41; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_42; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_43; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_44; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_45; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_46; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_47; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_48; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_49; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_50; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_51; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_52; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_53; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_54; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_55; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_56; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_57; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_58; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_59; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_60; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_61; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_62; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_63; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_64; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_65; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_66; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_67; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_68; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_69; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_70; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_71; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_72; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_73; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_74; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_75; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_76; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_77; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_78; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_79; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_80; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_81; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_82; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_83; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_84; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_85; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_86; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_87; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_88; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_89; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_90; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_91; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_92; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_93; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_94; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_95; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_96; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_97; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_98; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_99; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_100; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_101; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_102; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_103; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_104; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_105; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_106; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_107; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_108; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_109; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_110; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_111; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_112; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_113; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_114; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_115; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_116; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_117; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_118; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_119; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_120; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_121; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_122; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_123; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_124; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_125; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_126; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataIn_bits_127; // @[AWSVggWrapper.scala 79:24]
  wire  muxLyr_2_io_dataOut_valid; // @[AWSVggWrapper.scala 79:24]
  wire [15:0] muxLyr_2_io_dataOut_bits_0; // @[AWSVggWrapper.scala 79:24]
  wire  scale_clock; // @[AWSVggWrapper.scala 92:21]
  wire  scale_reset; // @[AWSVggWrapper.scala 92:21]
  wire  scale_io_dataIn_valid; // @[AWSVggWrapper.scala 92:21]
  wire [15:0] scale_io_dataIn_bits_0; // @[AWSVggWrapper.scala 92:21]
  wire  scale_io_dataOut_valid; // @[AWSVggWrapper.scala 92:21]
  wire [15:0] scale_io_dataOut_bits_0; // @[AWSVggWrapper.scala 92:21]
  wire  dense_2_clock; // @[AWSVggWrapper.scala 99:23]
  wire  dense_2_reset; // @[AWSVggWrapper.scala 99:23]
  wire  dense_2_io_dataIn_valid; // @[AWSVggWrapper.scala 99:23]
  wire [15:0] dense_2_io_dataIn_bits_0; // @[AWSVggWrapper.scala 99:23]
  wire  dense_2_io_dataOut_valid; // @[AWSVggWrapper.scala 99:23]
  wire [15:0] dense_2_io_dataOut_bits_0; // @[AWSVggWrapper.scala 99:23]
  wire [15:0] dense_2_io_dataOut_bits_1; // @[AWSVggWrapper.scala 99:23]
  wire [15:0] dense_2_io_dataOut_bits_2; // @[AWSVggWrapper.scala 99:23]
  wire [15:0] dense_2_io_dataOut_bits_3; // @[AWSVggWrapper.scala 99:23]
  wire [15:0] dense_2_io_dataOut_bits_4; // @[AWSVggWrapper.scala 99:23]
  wire [15:0] dense_2_io_dataOut_bits_5; // @[AWSVggWrapper.scala 99:23]
  wire [15:0] dense_2_io_dataOut_bits_6; // @[AWSVggWrapper.scala 99:23]
  wire [15:0] dense_2_io_dataOut_bits_7; // @[AWSVggWrapper.scala 99:23]
  wire [15:0] dense_2_io_dataOut_bits_8; // @[AWSVggWrapper.scala 99:23]
  wire [15:0] dense_2_io_dataOut_bits_9; // @[AWSVggWrapper.scala 99:23]
  reg [15:0] outputRegs_0; // @[AWSVggWrapper.scala 103:23]
  reg [31:0] _RAND_0;
  reg [15:0] outputRegs_1; // @[AWSVggWrapper.scala 103:23]
  reg [31:0] _RAND_1;
  reg [15:0] outputRegs_2; // @[AWSVggWrapper.scala 103:23]
  reg [31:0] _RAND_2;
  reg [15:0] outputRegs_3; // @[AWSVggWrapper.scala 103:23]
  reg [31:0] _RAND_3;
  reg [15:0] outputRegs_4; // @[AWSVggWrapper.scala 103:23]
  reg [31:0] _RAND_4;
  reg [15:0] outputRegs_5; // @[AWSVggWrapper.scala 103:23]
  reg [31:0] _RAND_5;
  reg [15:0] outputRegs_6; // @[AWSVggWrapper.scala 103:23]
  reg [31:0] _RAND_6;
  reg [15:0] outputRegs_7; // @[AWSVggWrapper.scala 103:23]
  reg [31:0] _RAND_7;
  reg [15:0] outputRegs_8; // @[AWSVggWrapper.scala 103:23]
  reg [31:0] _RAND_8;
  reg [15:0] outputRegs_9; // @[AWSVggWrapper.scala 103:23]
  reg [31:0] _RAND_9;
  reg  vldReg; // @[AWSVggWrapper.scala 106:23]
  reg [31:0] _RAND_10;
  wire [15:0] _T_35; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_36; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_37; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_38; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_39; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_40; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_41; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_42; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_43; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_44; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_45; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_46; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_47; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_48; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_49; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_50; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_51; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_52; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_53; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_54; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_55; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_56; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_57; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_58; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_59; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_60; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_61; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_62; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_63; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_64; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_65; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_66; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_67; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_68; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_69; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_70; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_71; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_72; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_73; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_74; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_75; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_76; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_77; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_78; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_79; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_80; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_81; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_82; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_83; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_84; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_85; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_86; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_87; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_88; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_89; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_90; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_91; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_92; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_93; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_94; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_95; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_96; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_97; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_98; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_99; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_100; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_101; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_102; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_103; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_104; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_105; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_106; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_107; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_108; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_109; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_110; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_111; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_112; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_113; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_114; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_115; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_116; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_117; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_118; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_119; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_120; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_121; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_122; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_123; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_124; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_125; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_126; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_127; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_128; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_129; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_130; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_131; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_132; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_133; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_134; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_135; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_136; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_137; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_138; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_139; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_140; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_141; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_142; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_143; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_144; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_145; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_146; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_147; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_148; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_149; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_150; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_151; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_152; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_153; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_154; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_155; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_156; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_157; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_158; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_159; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_160; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_161; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_162; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_163; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_164; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_165; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_166; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_167; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_168; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_169; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_170; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_171; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_172; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_173; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_174; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_175; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_176; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_177; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_178; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_179; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_180; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_181; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_182; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_183; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_184; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_185; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_186; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_187; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_188; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_189; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_190; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_191; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_192; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_193; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_194; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_195; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_196; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_197; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_198; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_199; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_200; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_201; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_202; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_203; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_204; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_205; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_206; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_207; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_208; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_209; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_210; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_211; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_212; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_213; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_214; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_215; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_216; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_217; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_218; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_219; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_220; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_221; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_222; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_223; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_224; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_225; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_226; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_227; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_228; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_229; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_230; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_231; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_232; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_233; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_234; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_235; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_236; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_237; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_238; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_239; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_240; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_241; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_242; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_243; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_244; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_245; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_246; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_247; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_248; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_249; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_250; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_251; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_252; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_253; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_254; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_255; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_256; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_257; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_258; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_259; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_260; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_261; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_262; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_263; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_264; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_265; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_266; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_267; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_268; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_269; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_270; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_271; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_272; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_273; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_274; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_275; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_276; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_277; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_278; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_279; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_280; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_281; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_282; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_283; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_284; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_285; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_286; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_287; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_288; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_289; // @[AWSVggWrapper.scala 53:79]
  wire [15:0] _T_290; // @[AWSVggWrapper.scala 53:79]
  wire [31:0] _T_291; // @[AWSVggWrapper.scala 53:94]
  wire [47:0] _T_292; // @[AWSVggWrapper.scala 53:94]
  wire [63:0] _T_293; // @[AWSVggWrapper.scala 53:94]
  wire [79:0] _T_294; // @[AWSVggWrapper.scala 53:94]
  wire [95:0] _T_295; // @[AWSVggWrapper.scala 53:94]
  wire [111:0] _T_296; // @[AWSVggWrapper.scala 53:94]
  wire [127:0] _T_297; // @[AWSVggWrapper.scala 53:94]
  wire [143:0] _T_298; // @[AWSVggWrapper.scala 53:94]
  wire [159:0] _T_299; // @[AWSVggWrapper.scala 53:94]
  wire [175:0] _T_300; // @[AWSVggWrapper.scala 53:94]
  wire [191:0] _T_301; // @[AWSVggWrapper.scala 53:94]
  wire [207:0] _T_302; // @[AWSVggWrapper.scala 53:94]
  wire [223:0] _T_303; // @[AWSVggWrapper.scala 53:94]
  wire [239:0] _T_304; // @[AWSVggWrapper.scala 53:94]
  wire [255:0] _T_305; // @[AWSVggWrapper.scala 53:94]
  wire [271:0] _T_306; // @[AWSVggWrapper.scala 53:94]
  wire [287:0] _T_307; // @[AWSVggWrapper.scala 53:94]
  wire [303:0] _T_308; // @[AWSVggWrapper.scala 53:94]
  wire [319:0] _T_309; // @[AWSVggWrapper.scala 53:94]
  wire [335:0] _T_310; // @[AWSVggWrapper.scala 53:94]
  wire [351:0] _T_311; // @[AWSVggWrapper.scala 53:94]
  wire [367:0] _T_312; // @[AWSVggWrapper.scala 53:94]
  wire [383:0] _T_313; // @[AWSVggWrapper.scala 53:94]
  wire [399:0] _T_314; // @[AWSVggWrapper.scala 53:94]
  wire [415:0] _T_315; // @[AWSVggWrapper.scala 53:94]
  wire [431:0] _T_316; // @[AWSVggWrapper.scala 53:94]
  wire [447:0] _T_317; // @[AWSVggWrapper.scala 53:94]
  wire [463:0] _T_318; // @[AWSVggWrapper.scala 53:94]
  wire [479:0] _T_319; // @[AWSVggWrapper.scala 53:94]
  wire [495:0] _T_320; // @[AWSVggWrapper.scala 53:94]
  wire [511:0] _T_321; // @[AWSVggWrapper.scala 53:94]
  wire [527:0] _T_322; // @[AWSVggWrapper.scala 53:94]
  wire [543:0] _T_323; // @[AWSVggWrapper.scala 53:94]
  wire [559:0] _T_324; // @[AWSVggWrapper.scala 53:94]
  wire [575:0] _T_325; // @[AWSVggWrapper.scala 53:94]
  wire [591:0] _T_326; // @[AWSVggWrapper.scala 53:94]
  wire [607:0] _T_327; // @[AWSVggWrapper.scala 53:94]
  wire [623:0] _T_328; // @[AWSVggWrapper.scala 53:94]
  wire [639:0] _T_329; // @[AWSVggWrapper.scala 53:94]
  wire [655:0] _T_330; // @[AWSVggWrapper.scala 53:94]
  wire [671:0] _T_331; // @[AWSVggWrapper.scala 53:94]
  wire [687:0] _T_332; // @[AWSVggWrapper.scala 53:94]
  wire [703:0] _T_333; // @[AWSVggWrapper.scala 53:94]
  wire [719:0] _T_334; // @[AWSVggWrapper.scala 53:94]
  wire [735:0] _T_335; // @[AWSVggWrapper.scala 53:94]
  wire [751:0] _T_336; // @[AWSVggWrapper.scala 53:94]
  wire [767:0] _T_337; // @[AWSVggWrapper.scala 53:94]
  wire [783:0] _T_338; // @[AWSVggWrapper.scala 53:94]
  wire [799:0] _T_339; // @[AWSVggWrapper.scala 53:94]
  wire [815:0] _T_340; // @[AWSVggWrapper.scala 53:94]
  wire [831:0] _T_341; // @[AWSVggWrapper.scala 53:94]
  wire [847:0] _T_342; // @[AWSVggWrapper.scala 53:94]
  wire [863:0] _T_343; // @[AWSVggWrapper.scala 53:94]
  wire [879:0] _T_344; // @[AWSVggWrapper.scala 53:94]
  wire [895:0] _T_345; // @[AWSVggWrapper.scala 53:94]
  wire [911:0] _T_346; // @[AWSVggWrapper.scala 53:94]
  wire [927:0] _T_347; // @[AWSVggWrapper.scala 53:94]
  wire [943:0] _T_348; // @[AWSVggWrapper.scala 53:94]
  wire [959:0] _T_349; // @[AWSVggWrapper.scala 53:94]
  wire [975:0] _T_350; // @[AWSVggWrapper.scala 53:94]
  wire [991:0] _T_351; // @[AWSVggWrapper.scala 53:94]
  wire [1007:0] _T_352; // @[AWSVggWrapper.scala 53:94]
  wire [1023:0] _T_353; // @[AWSVggWrapper.scala 53:94]
  wire [1039:0] _T_354; // @[AWSVggWrapper.scala 53:94]
  wire [1055:0] _T_355; // @[AWSVggWrapper.scala 53:94]
  wire [1071:0] _T_356; // @[AWSVggWrapper.scala 53:94]
  wire [1087:0] _T_357; // @[AWSVggWrapper.scala 53:94]
  wire [1103:0] _T_358; // @[AWSVggWrapper.scala 53:94]
  wire [1119:0] _T_359; // @[AWSVggWrapper.scala 53:94]
  wire [1135:0] _T_360; // @[AWSVggWrapper.scala 53:94]
  wire [1151:0] _T_361; // @[AWSVggWrapper.scala 53:94]
  wire [1167:0] _T_362; // @[AWSVggWrapper.scala 53:94]
  wire [1183:0] _T_363; // @[AWSVggWrapper.scala 53:94]
  wire [1199:0] _T_364; // @[AWSVggWrapper.scala 53:94]
  wire [1215:0] _T_365; // @[AWSVggWrapper.scala 53:94]
  wire [1231:0] _T_366; // @[AWSVggWrapper.scala 53:94]
  wire [1247:0] _T_367; // @[AWSVggWrapper.scala 53:94]
  wire [1263:0] _T_368; // @[AWSVggWrapper.scala 53:94]
  wire [1279:0] _T_369; // @[AWSVggWrapper.scala 53:94]
  wire [1295:0] _T_370; // @[AWSVggWrapper.scala 53:94]
  wire [1311:0] _T_371; // @[AWSVggWrapper.scala 53:94]
  wire [1327:0] _T_372; // @[AWSVggWrapper.scala 53:94]
  wire [1343:0] _T_373; // @[AWSVggWrapper.scala 53:94]
  wire [1359:0] _T_374; // @[AWSVggWrapper.scala 53:94]
  wire [1375:0] _T_375; // @[AWSVggWrapper.scala 53:94]
  wire [1391:0] _T_376; // @[AWSVggWrapper.scala 53:94]
  wire [1407:0] _T_377; // @[AWSVggWrapper.scala 53:94]
  wire [1423:0] _T_378; // @[AWSVggWrapper.scala 53:94]
  wire [1439:0] _T_379; // @[AWSVggWrapper.scala 53:94]
  wire [1455:0] _T_380; // @[AWSVggWrapper.scala 53:94]
  wire [1471:0] _T_381; // @[AWSVggWrapper.scala 53:94]
  wire [1487:0] _T_382; // @[AWSVggWrapper.scala 53:94]
  wire [1503:0] _T_383; // @[AWSVggWrapper.scala 53:94]
  wire [1519:0] _T_384; // @[AWSVggWrapper.scala 53:94]
  wire [1535:0] _T_385; // @[AWSVggWrapper.scala 53:94]
  wire [1551:0] _T_386; // @[AWSVggWrapper.scala 53:94]
  wire [1567:0] _T_387; // @[AWSVggWrapper.scala 53:94]
  wire [1583:0] _T_388; // @[AWSVggWrapper.scala 53:94]
  wire [1599:0] _T_389; // @[AWSVggWrapper.scala 53:94]
  wire [1615:0] _T_390; // @[AWSVggWrapper.scala 53:94]
  wire [1631:0] _T_391; // @[AWSVggWrapper.scala 53:94]
  wire [1647:0] _T_392; // @[AWSVggWrapper.scala 53:94]
  wire [1663:0] _T_393; // @[AWSVggWrapper.scala 53:94]
  wire [1679:0] _T_394; // @[AWSVggWrapper.scala 53:94]
  wire [1695:0] _T_395; // @[AWSVggWrapper.scala 53:94]
  wire [1711:0] _T_396; // @[AWSVggWrapper.scala 53:94]
  wire [1727:0] _T_397; // @[AWSVggWrapper.scala 53:94]
  wire [1743:0] _T_398; // @[AWSVggWrapper.scala 53:94]
  wire [1759:0] _T_399; // @[AWSVggWrapper.scala 53:94]
  wire [1775:0] _T_400; // @[AWSVggWrapper.scala 53:94]
  wire [1791:0] _T_401; // @[AWSVggWrapper.scala 53:94]
  wire [1807:0] _T_402; // @[AWSVggWrapper.scala 53:94]
  wire [1823:0] _T_403; // @[AWSVggWrapper.scala 53:94]
  wire [1839:0] _T_404; // @[AWSVggWrapper.scala 53:94]
  wire [1855:0] _T_405; // @[AWSVggWrapper.scala 53:94]
  wire [1871:0] _T_406; // @[AWSVggWrapper.scala 53:94]
  wire [1887:0] _T_407; // @[AWSVggWrapper.scala 53:94]
  wire [1903:0] _T_408; // @[AWSVggWrapper.scala 53:94]
  wire [1919:0] _T_409; // @[AWSVggWrapper.scala 53:94]
  wire [1935:0] _T_410; // @[AWSVggWrapper.scala 53:94]
  wire [1951:0] _T_411; // @[AWSVggWrapper.scala 53:94]
  wire [1967:0] _T_412; // @[AWSVggWrapper.scala 53:94]
  wire [1983:0] _T_413; // @[AWSVggWrapper.scala 53:94]
  wire [1999:0] _T_414; // @[AWSVggWrapper.scala 53:94]
  wire [2015:0] _T_415; // @[AWSVggWrapper.scala 53:94]
  wire [2031:0] _T_416; // @[AWSVggWrapper.scala 53:94]
  wire [2047:0] _T_417; // @[AWSVggWrapper.scala 53:94]
  wire [2063:0] _T_418; // @[AWSVggWrapper.scala 53:94]
  wire [2079:0] _T_419; // @[AWSVggWrapper.scala 53:94]
  wire [2095:0] _T_420; // @[AWSVggWrapper.scala 53:94]
  wire [2111:0] _T_421; // @[AWSVggWrapper.scala 53:94]
  wire [2127:0] _T_422; // @[AWSVggWrapper.scala 53:94]
  wire [2143:0] _T_423; // @[AWSVggWrapper.scala 53:94]
  wire [2159:0] _T_424; // @[AWSVggWrapper.scala 53:94]
  wire [2175:0] _T_425; // @[AWSVggWrapper.scala 53:94]
  wire [2191:0] _T_426; // @[AWSVggWrapper.scala 53:94]
  wire [2207:0] _T_427; // @[AWSVggWrapper.scala 53:94]
  wire [2223:0] _T_428; // @[AWSVggWrapper.scala 53:94]
  wire [2239:0] _T_429; // @[AWSVggWrapper.scala 53:94]
  wire [2255:0] _T_430; // @[AWSVggWrapper.scala 53:94]
  wire [2271:0] _T_431; // @[AWSVggWrapper.scala 53:94]
  wire [2287:0] _T_432; // @[AWSVggWrapper.scala 53:94]
  wire [2303:0] _T_433; // @[AWSVggWrapper.scala 53:94]
  wire [2319:0] _T_434; // @[AWSVggWrapper.scala 53:94]
  wire [2335:0] _T_435; // @[AWSVggWrapper.scala 53:94]
  wire [2351:0] _T_436; // @[AWSVggWrapper.scala 53:94]
  wire [2367:0] _T_437; // @[AWSVggWrapper.scala 53:94]
  wire [2383:0] _T_438; // @[AWSVggWrapper.scala 53:94]
  wire [2399:0] _T_439; // @[AWSVggWrapper.scala 53:94]
  wire [2415:0] _T_440; // @[AWSVggWrapper.scala 53:94]
  wire [2431:0] _T_441; // @[AWSVggWrapper.scala 53:94]
  wire [2447:0] _T_442; // @[AWSVggWrapper.scala 53:94]
  wire [2463:0] _T_443; // @[AWSVggWrapper.scala 53:94]
  wire [2479:0] _T_444; // @[AWSVggWrapper.scala 53:94]
  wire [2495:0] _T_445; // @[AWSVggWrapper.scala 53:94]
  wire [2511:0] _T_446; // @[AWSVggWrapper.scala 53:94]
  wire [2527:0] _T_447; // @[AWSVggWrapper.scala 53:94]
  wire [2543:0] _T_448; // @[AWSVggWrapper.scala 53:94]
  wire [2559:0] _T_449; // @[AWSVggWrapper.scala 53:94]
  wire [2575:0] _T_450; // @[AWSVggWrapper.scala 53:94]
  wire [2591:0] _T_451; // @[AWSVggWrapper.scala 53:94]
  wire [2607:0] _T_452; // @[AWSVggWrapper.scala 53:94]
  wire [2623:0] _T_453; // @[AWSVggWrapper.scala 53:94]
  wire [2639:0] _T_454; // @[AWSVggWrapper.scala 53:94]
  wire [2655:0] _T_455; // @[AWSVggWrapper.scala 53:94]
  wire [2671:0] _T_456; // @[AWSVggWrapper.scala 53:94]
  wire [2687:0] _T_457; // @[AWSVggWrapper.scala 53:94]
  wire [2703:0] _T_458; // @[AWSVggWrapper.scala 53:94]
  wire [2719:0] _T_459; // @[AWSVggWrapper.scala 53:94]
  wire [2735:0] _T_460; // @[AWSVggWrapper.scala 53:94]
  wire [2751:0] _T_461; // @[AWSVggWrapper.scala 53:94]
  wire [2767:0] _T_462; // @[AWSVggWrapper.scala 53:94]
  wire [2783:0] _T_463; // @[AWSVggWrapper.scala 53:94]
  wire [2799:0] _T_464; // @[AWSVggWrapper.scala 53:94]
  wire [2815:0] _T_465; // @[AWSVggWrapper.scala 53:94]
  wire [2831:0] _T_466; // @[AWSVggWrapper.scala 53:94]
  wire [2847:0] _T_467; // @[AWSVggWrapper.scala 53:94]
  wire [2863:0] _T_468; // @[AWSVggWrapper.scala 53:94]
  wire [2879:0] _T_469; // @[AWSVggWrapper.scala 53:94]
  wire [2895:0] _T_470; // @[AWSVggWrapper.scala 53:94]
  wire [2911:0] _T_471; // @[AWSVggWrapper.scala 53:94]
  wire [2927:0] _T_472; // @[AWSVggWrapper.scala 53:94]
  wire [2943:0] _T_473; // @[AWSVggWrapper.scala 53:94]
  wire [2959:0] _T_474; // @[AWSVggWrapper.scala 53:94]
  wire [2975:0] _T_475; // @[AWSVggWrapper.scala 53:94]
  wire [2991:0] _T_476; // @[AWSVggWrapper.scala 53:94]
  wire [3007:0] _T_477; // @[AWSVggWrapper.scala 53:94]
  wire [3023:0] _T_478; // @[AWSVggWrapper.scala 53:94]
  wire [3039:0] _T_479; // @[AWSVggWrapper.scala 53:94]
  wire [3055:0] _T_480; // @[AWSVggWrapper.scala 53:94]
  wire [3071:0] _T_481; // @[AWSVggWrapper.scala 53:94]
  wire [3087:0] _T_482; // @[AWSVggWrapper.scala 53:94]
  wire [3103:0] _T_483; // @[AWSVggWrapper.scala 53:94]
  wire [3119:0] _T_484; // @[AWSVggWrapper.scala 53:94]
  wire [3135:0] _T_485; // @[AWSVggWrapper.scala 53:94]
  wire [3151:0] _T_486; // @[AWSVggWrapper.scala 53:94]
  wire [3167:0] _T_487; // @[AWSVggWrapper.scala 53:94]
  wire [3183:0] _T_488; // @[AWSVggWrapper.scala 53:94]
  wire [3199:0] _T_489; // @[AWSVggWrapper.scala 53:94]
  wire [3215:0] _T_490; // @[AWSVggWrapper.scala 53:94]
  wire [3231:0] _T_491; // @[AWSVggWrapper.scala 53:94]
  wire [3247:0] _T_492; // @[AWSVggWrapper.scala 53:94]
  wire [3263:0] _T_493; // @[AWSVggWrapper.scala 53:94]
  wire [3279:0] _T_494; // @[AWSVggWrapper.scala 53:94]
  wire [3295:0] _T_495; // @[AWSVggWrapper.scala 53:94]
  wire [3311:0] _T_496; // @[AWSVggWrapper.scala 53:94]
  wire [3327:0] _T_497; // @[AWSVggWrapper.scala 53:94]
  wire [3343:0] _T_498; // @[AWSVggWrapper.scala 53:94]
  wire [3359:0] _T_499; // @[AWSVggWrapper.scala 53:94]
  wire [3375:0] _T_500; // @[AWSVggWrapper.scala 53:94]
  wire [3391:0] _T_501; // @[AWSVggWrapper.scala 53:94]
  wire [3407:0] _T_502; // @[AWSVggWrapper.scala 53:94]
  wire [3423:0] _T_503; // @[AWSVggWrapper.scala 53:94]
  wire [3439:0] _T_504; // @[AWSVggWrapper.scala 53:94]
  wire [3455:0] _T_505; // @[AWSVggWrapper.scala 53:94]
  wire [3471:0] _T_506; // @[AWSVggWrapper.scala 53:94]
  wire [3487:0] _T_507; // @[AWSVggWrapper.scala 53:94]
  wire [3503:0] _T_508; // @[AWSVggWrapper.scala 53:94]
  wire [3519:0] _T_509; // @[AWSVggWrapper.scala 53:94]
  wire [3535:0] _T_510; // @[AWSVggWrapper.scala 53:94]
  wire [3551:0] _T_511; // @[AWSVggWrapper.scala 53:94]
  wire [3567:0] _T_512; // @[AWSVggWrapper.scala 53:94]
  wire [3583:0] _T_513; // @[AWSVggWrapper.scala 53:94]
  wire [3599:0] _T_514; // @[AWSVggWrapper.scala 53:94]
  wire [3615:0] _T_515; // @[AWSVggWrapper.scala 53:94]
  wire [3631:0] _T_516; // @[AWSVggWrapper.scala 53:94]
  wire [3647:0] _T_517; // @[AWSVggWrapper.scala 53:94]
  wire [3663:0] _T_518; // @[AWSVggWrapper.scala 53:94]
  wire [3679:0] _T_519; // @[AWSVggWrapper.scala 53:94]
  wire [3695:0] _T_520; // @[AWSVggWrapper.scala 53:94]
  wire [3711:0] _T_521; // @[AWSVggWrapper.scala 53:94]
  wire [3727:0] _T_522; // @[AWSVggWrapper.scala 53:94]
  wire [3743:0] _T_523; // @[AWSVggWrapper.scala 53:94]
  wire [3759:0] _T_524; // @[AWSVggWrapper.scala 53:94]
  wire [3775:0] _T_525; // @[AWSVggWrapper.scala 53:94]
  wire [3791:0] _T_526; // @[AWSVggWrapper.scala 53:94]
  wire [3807:0] _T_527; // @[AWSVggWrapper.scala 53:94]
  wire [3823:0] _T_528; // @[AWSVggWrapper.scala 53:94]
  wire [3839:0] _T_529; // @[AWSVggWrapper.scala 53:94]
  wire [3855:0] _T_530; // @[AWSVggWrapper.scala 53:94]
  wire [3871:0] _T_531; // @[AWSVggWrapper.scala 53:94]
  wire [3887:0] _T_532; // @[AWSVggWrapper.scala 53:94]
  wire [3903:0] _T_533; // @[AWSVggWrapper.scala 53:94]
  wire [3919:0] _T_534; // @[AWSVggWrapper.scala 53:94]
  wire [3935:0] _T_535; // @[AWSVggWrapper.scala 53:94]
  wire [3951:0] _T_536; // @[AWSVggWrapper.scala 53:94]
  wire [3967:0] _T_537; // @[AWSVggWrapper.scala 53:94]
  wire [3983:0] _T_538; // @[AWSVggWrapper.scala 53:94]
  wire [3999:0] _T_539; // @[AWSVggWrapper.scala 53:94]
  wire [4015:0] _T_540; // @[AWSVggWrapper.scala 53:94]
  wire [4031:0] _T_541; // @[AWSVggWrapper.scala 53:94]
  wire [4047:0] _T_542; // @[AWSVggWrapper.scala 53:94]
  wire [4063:0] _T_543; // @[AWSVggWrapper.scala 53:94]
  wire [4079:0] _T_544; // @[AWSVggWrapper.scala 53:94]
  wire [4095:0] dataInAsUInt; // @[AWSVggWrapper.scala 53:94]
  wire [15:0] _T_1839; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_255; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1841; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_254; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1843; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_253; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1845; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_252; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1847; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_251; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1849; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_250; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1851; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_249; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1853; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_248; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1855; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_247; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1857; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_246; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1859; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_245; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1861; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_244; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1863; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_243; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1865; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_242; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1867; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_241; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1869; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_240; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1871; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_239; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1873; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_238; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1875; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_237; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1877; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_236; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1879; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_235; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1881; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_234; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1883; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_233; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1885; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_232; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1887; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_231; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1889; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_230; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1891; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_229; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1893; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_228; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1895; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_227; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1897; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_226; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1899; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_225; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1901; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_224; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1903; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_223; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1905; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_222; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1907; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_221; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1909; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_220; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1911; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_219; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1913; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_218; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1915; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_217; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1917; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_216; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1919; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_215; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1921; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_214; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1923; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_213; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1925; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_212; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1927; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_211; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1929; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_210; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1931; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_209; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1933; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_208; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1935; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_207; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1937; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_206; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1939; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_205; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1941; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_204; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1943; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_203; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1945; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_202; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1947; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_201; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1949; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_200; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1951; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_199; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1953; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_198; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1955; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_197; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1957; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_196; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1959; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_195; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1961; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_194; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1963; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_193; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1965; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_192; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1967; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_191; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1969; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_190; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1971; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_189; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1973; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_188; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1975; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_187; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1977; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_186; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1979; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_185; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1981; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_184; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1983; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_183; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1985; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_182; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1987; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_181; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1989; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_180; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1991; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_179; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1993; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_178; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1995; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_177; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1997; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_176; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_1999; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_175; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2001; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_174; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2003; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_173; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2005; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_172; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2007; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_171; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2009; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_170; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2011; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_169; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2013; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_168; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2015; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_167; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2017; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_166; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2019; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_165; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2021; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_164; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2023; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_163; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2025; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_162; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2027; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_161; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2029; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_160; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2031; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_159; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2033; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_158; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2035; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_157; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2037; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_156; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2039; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_155; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2041; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_154; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2043; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_153; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2045; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_152; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2047; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_151; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2049; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_150; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2051; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_149; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2053; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_148; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2055; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_147; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2057; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_146; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2059; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_145; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2061; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_144; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2063; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_143; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2065; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_142; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2067; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_141; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2069; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_140; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2071; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_139; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2073; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_138; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2075; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_137; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2077; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_136; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2079; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_135; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2081; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_134; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2083; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_133; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2085; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_132; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2087; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_131; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2089; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_130; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2091; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_129; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2093; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_128; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2095; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_127; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2097; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_126; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2099; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_125; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2101; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_124; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2103; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_123; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2105; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_122; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2107; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_121; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2109; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_120; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2111; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_119; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2113; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_118; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2115; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_117; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2117; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_116; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2119; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_115; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2121; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_114; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2123; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_113; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2125; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_112; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2127; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_111; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2129; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_110; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2131; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_109; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2133; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_108; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2135; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_107; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2137; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_106; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2139; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_105; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2141; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_104; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2143; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_103; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2145; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_102; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2147; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_101; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2149; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_100; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2151; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_99; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2153; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_98; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2155; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_97; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2157; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_96; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2159; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_95; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2161; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_94; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2163; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_93; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2165; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_92; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2167; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_91; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2169; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_90; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2171; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_89; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2173; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_88; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2175; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_87; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2177; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_86; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2179; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_85; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2181; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_84; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2183; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_83; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2185; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_82; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2187; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_81; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2189; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_80; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2191; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_79; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2193; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_78; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2195; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_77; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2197; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_76; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2199; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_75; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2201; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_74; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2203; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_73; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2205; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_72; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2207; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_71; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2209; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_70; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2211; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_69; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2213; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_68; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2215; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_67; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2217; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_66; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2219; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_65; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2221; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_64; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2223; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_63; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2225; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_62; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2227; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_61; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2229; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_60; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2231; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_59; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2233; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_58; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2235; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_57; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2237; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_56; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2239; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_55; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2241; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_54; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2243; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_53; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2245; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_52; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2247; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_51; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2249; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_50; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2251; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_49; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2253; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_48; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2255; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_47; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2257; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_46; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2259; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_45; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2261; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_44; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2263; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_43; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2265; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_42; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2267; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_41; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2269; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_40; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2271; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_39; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2273; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_38; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2275; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_37; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2277; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_36; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2279; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_35; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2281; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_34; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2283; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_33; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2285; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_32; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2287; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_31; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2289; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_30; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2291; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_29; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2293; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_28; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2295; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_27; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2297; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_26; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2299; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_25; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2301; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_24; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2303; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_23; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2305; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_22; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2307; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_21; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2309; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_20; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2311; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_19; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2313; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_18; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2315; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_17; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2317; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_16; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2319; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_15; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2321; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_14; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2323; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_13; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2325; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_12; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2327; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_11; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2329; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_10; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2331; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_9; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2333; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_8; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2335; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_7; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2337; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_6; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2339; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_5; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2341; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_4; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2343; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_3; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2345; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_2; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2347; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_1; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _T_2349; // @[AWSVggWrapper.scala 64:67]
  wire [15:0] sintOut_0; // @[AWSVggWrapper.scala 64:110]
  wire [15:0] _GEN_0; // @[AWSVggWrapper.scala 109:37]
  wire [15:0] _GEN_1; // @[AWSVggWrapper.scala 109:37]
  wire [15:0] _GEN_2; // @[AWSVggWrapper.scala 109:37]
  wire [15:0] _GEN_3; // @[AWSVggWrapper.scala 109:37]
  wire [15:0] _GEN_4; // @[AWSVggWrapper.scala 109:37]
  wire [15:0] _GEN_5; // @[AWSVggWrapper.scala 109:37]
  wire [15:0] _GEN_6; // @[AWSVggWrapper.scala 109:37]
  wire [15:0] _GEN_7; // @[AWSVggWrapper.scala 109:37]
  wire [15:0] _GEN_8; // @[AWSVggWrapper.scala 109:37]
  wire [15:0] _GEN_9; // @[AWSVggWrapper.scala 109:37]
  wire  _GEN_10; // @[AWSVggWrapper.scala 109:37]
  wire  queueIOIn_ready; // @[AWSVggWrapper.scala 54:23]
  wire  queueIOIn_valid; // @[AWSVggWrapper.scala 54:23]
  wire [15:0] _T_2353_0; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_1; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_2; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_3; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_4; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_5; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_6; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_7; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_8; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_9; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_10; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_11; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_12; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_13; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_14; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_15; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_16; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_17; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_18; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_19; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_20; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_21; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_22; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_23; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_24; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_25; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_26; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_27; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_28; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_29; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_30; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_31; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_32; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_33; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_34; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_35; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_36; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_37; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_38; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_39; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_40; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_41; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_42; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_43; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_44; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_45; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_46; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_47; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_48; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_49; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_50; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_51; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_52; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_53; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_54; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_55; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_56; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_57; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_58; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_59; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_60; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_61; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_62; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_63; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_64; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_65; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_66; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_67; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_68; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_69; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_70; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_71; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_72; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_73; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_74; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_75; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_76; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_77; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_78; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_79; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_80; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_81; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_82; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_83; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_84; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_85; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_86; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_87; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_88; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_89; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_90; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_91; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_92; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_93; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_94; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_95; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_96; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_97; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_98; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_99; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_100; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_101; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_102; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_103; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_104; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_105; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_106; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_107; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_108; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_109; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_110; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_111; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_112; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_113; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_114; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_115; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_116; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_117; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_118; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_119; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_120; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_121; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_122; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_123; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_124; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_125; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_126; // @[AWSVggWrapper.scala 83:33]
  wire [15:0] _T_2353_127; // @[AWSVggWrapper.scala 83:33]
  Vgg7 vgg ( // @[AWSVggWrapper.scala 47:27]
    .clock(vgg_clock),
    .reset(vgg_reset),
    .io_dataIn_ready(vgg_io_dataIn_ready),
    .io_dataIn_valid(vgg_io_dataIn_valid),
    .io_dataIn_bits_0(vgg_io_dataIn_bits_0),
    .io_dataIn_bits_1(vgg_io_dataIn_bits_1),
    .io_dataIn_bits_2(vgg_io_dataIn_bits_2),
    .io_dataOut_ready(vgg_io_dataOut_ready),
    .io_dataOut_valid(vgg_io_dataOut_valid),
    .io_dataOut_bits_0(vgg_io_dataOut_bits_0),
    .io_dataOut_bits_1(vgg_io_dataOut_bits_1),
    .io_dataOut_bits_2(vgg_io_dataOut_bits_2),
    .io_dataOut_bits_3(vgg_io_dataOut_bits_3),
    .io_dataOut_bits_4(vgg_io_dataOut_bits_4),
    .io_dataOut_bits_5(vgg_io_dataOut_bits_5),
    .io_dataOut_bits_6(vgg_io_dataOut_bits_6),
    .io_dataOut_bits_7(vgg_io_dataOut_bits_7),
    .io_dataOut_bits_8(vgg_io_dataOut_bits_8),
    .io_dataOut_bits_9(vgg_io_dataOut_bits_9),
    .io_dataOut_bits_10(vgg_io_dataOut_bits_10),
    .io_dataOut_bits_11(vgg_io_dataOut_bits_11),
    .io_dataOut_bits_12(vgg_io_dataOut_bits_12),
    .io_dataOut_bits_13(vgg_io_dataOut_bits_13),
    .io_dataOut_bits_14(vgg_io_dataOut_bits_14),
    .io_dataOut_bits_15(vgg_io_dataOut_bits_15),
    .io_dataOut_bits_16(vgg_io_dataOut_bits_16),
    .io_dataOut_bits_17(vgg_io_dataOut_bits_17),
    .io_dataOut_bits_18(vgg_io_dataOut_bits_18),
    .io_dataOut_bits_19(vgg_io_dataOut_bits_19),
    .io_dataOut_bits_20(vgg_io_dataOut_bits_20),
    .io_dataOut_bits_21(vgg_io_dataOut_bits_21),
    .io_dataOut_bits_22(vgg_io_dataOut_bits_22),
    .io_dataOut_bits_23(vgg_io_dataOut_bits_23),
    .io_dataOut_bits_24(vgg_io_dataOut_bits_24),
    .io_dataOut_bits_25(vgg_io_dataOut_bits_25),
    .io_dataOut_bits_26(vgg_io_dataOut_bits_26),
    .io_dataOut_bits_27(vgg_io_dataOut_bits_27),
    .io_dataOut_bits_28(vgg_io_dataOut_bits_28),
    .io_dataOut_bits_29(vgg_io_dataOut_bits_29),
    .io_dataOut_bits_30(vgg_io_dataOut_bits_30),
    .io_dataOut_bits_31(vgg_io_dataOut_bits_31),
    .io_dataOut_bits_32(vgg_io_dataOut_bits_32),
    .io_dataOut_bits_33(vgg_io_dataOut_bits_33),
    .io_dataOut_bits_34(vgg_io_dataOut_bits_34),
    .io_dataOut_bits_35(vgg_io_dataOut_bits_35),
    .io_dataOut_bits_36(vgg_io_dataOut_bits_36),
    .io_dataOut_bits_37(vgg_io_dataOut_bits_37),
    .io_dataOut_bits_38(vgg_io_dataOut_bits_38),
    .io_dataOut_bits_39(vgg_io_dataOut_bits_39),
    .io_dataOut_bits_40(vgg_io_dataOut_bits_40),
    .io_dataOut_bits_41(vgg_io_dataOut_bits_41),
    .io_dataOut_bits_42(vgg_io_dataOut_bits_42),
    .io_dataOut_bits_43(vgg_io_dataOut_bits_43),
    .io_dataOut_bits_44(vgg_io_dataOut_bits_44),
    .io_dataOut_bits_45(vgg_io_dataOut_bits_45),
    .io_dataOut_bits_46(vgg_io_dataOut_bits_46),
    .io_dataOut_bits_47(vgg_io_dataOut_bits_47),
    .io_dataOut_bits_48(vgg_io_dataOut_bits_48),
    .io_dataOut_bits_49(vgg_io_dataOut_bits_49),
    .io_dataOut_bits_50(vgg_io_dataOut_bits_50),
    .io_dataOut_bits_51(vgg_io_dataOut_bits_51),
    .io_dataOut_bits_52(vgg_io_dataOut_bits_52),
    .io_dataOut_bits_53(vgg_io_dataOut_bits_53),
    .io_dataOut_bits_54(vgg_io_dataOut_bits_54),
    .io_dataOut_bits_55(vgg_io_dataOut_bits_55),
    .io_dataOut_bits_56(vgg_io_dataOut_bits_56),
    .io_dataOut_bits_57(vgg_io_dataOut_bits_57),
    .io_dataOut_bits_58(vgg_io_dataOut_bits_58),
    .io_dataOut_bits_59(vgg_io_dataOut_bits_59),
    .io_dataOut_bits_60(vgg_io_dataOut_bits_60),
    .io_dataOut_bits_61(vgg_io_dataOut_bits_61),
    .io_dataOut_bits_62(vgg_io_dataOut_bits_62),
    .io_dataOut_bits_63(vgg_io_dataOut_bits_63),
    .io_dataOut_bits_64(vgg_io_dataOut_bits_64),
    .io_dataOut_bits_65(vgg_io_dataOut_bits_65),
    .io_dataOut_bits_66(vgg_io_dataOut_bits_66),
    .io_dataOut_bits_67(vgg_io_dataOut_bits_67),
    .io_dataOut_bits_68(vgg_io_dataOut_bits_68),
    .io_dataOut_bits_69(vgg_io_dataOut_bits_69),
    .io_dataOut_bits_70(vgg_io_dataOut_bits_70),
    .io_dataOut_bits_71(vgg_io_dataOut_bits_71),
    .io_dataOut_bits_72(vgg_io_dataOut_bits_72),
    .io_dataOut_bits_73(vgg_io_dataOut_bits_73),
    .io_dataOut_bits_74(vgg_io_dataOut_bits_74),
    .io_dataOut_bits_75(vgg_io_dataOut_bits_75),
    .io_dataOut_bits_76(vgg_io_dataOut_bits_76),
    .io_dataOut_bits_77(vgg_io_dataOut_bits_77),
    .io_dataOut_bits_78(vgg_io_dataOut_bits_78),
    .io_dataOut_bits_79(vgg_io_dataOut_bits_79),
    .io_dataOut_bits_80(vgg_io_dataOut_bits_80),
    .io_dataOut_bits_81(vgg_io_dataOut_bits_81),
    .io_dataOut_bits_82(vgg_io_dataOut_bits_82),
    .io_dataOut_bits_83(vgg_io_dataOut_bits_83),
    .io_dataOut_bits_84(vgg_io_dataOut_bits_84),
    .io_dataOut_bits_85(vgg_io_dataOut_bits_85),
    .io_dataOut_bits_86(vgg_io_dataOut_bits_86),
    .io_dataOut_bits_87(vgg_io_dataOut_bits_87),
    .io_dataOut_bits_88(vgg_io_dataOut_bits_88),
    .io_dataOut_bits_89(vgg_io_dataOut_bits_89),
    .io_dataOut_bits_90(vgg_io_dataOut_bits_90),
    .io_dataOut_bits_91(vgg_io_dataOut_bits_91),
    .io_dataOut_bits_92(vgg_io_dataOut_bits_92),
    .io_dataOut_bits_93(vgg_io_dataOut_bits_93),
    .io_dataOut_bits_94(vgg_io_dataOut_bits_94),
    .io_dataOut_bits_95(vgg_io_dataOut_bits_95),
    .io_dataOut_bits_96(vgg_io_dataOut_bits_96),
    .io_dataOut_bits_97(vgg_io_dataOut_bits_97),
    .io_dataOut_bits_98(vgg_io_dataOut_bits_98),
    .io_dataOut_bits_99(vgg_io_dataOut_bits_99),
    .io_dataOut_bits_100(vgg_io_dataOut_bits_100),
    .io_dataOut_bits_101(vgg_io_dataOut_bits_101),
    .io_dataOut_bits_102(vgg_io_dataOut_bits_102),
    .io_dataOut_bits_103(vgg_io_dataOut_bits_103),
    .io_dataOut_bits_104(vgg_io_dataOut_bits_104),
    .io_dataOut_bits_105(vgg_io_dataOut_bits_105),
    .io_dataOut_bits_106(vgg_io_dataOut_bits_106),
    .io_dataOut_bits_107(vgg_io_dataOut_bits_107),
    .io_dataOut_bits_108(vgg_io_dataOut_bits_108),
    .io_dataOut_bits_109(vgg_io_dataOut_bits_109),
    .io_dataOut_bits_110(vgg_io_dataOut_bits_110),
    .io_dataOut_bits_111(vgg_io_dataOut_bits_111),
    .io_dataOut_bits_112(vgg_io_dataOut_bits_112),
    .io_dataOut_bits_113(vgg_io_dataOut_bits_113),
    .io_dataOut_bits_114(vgg_io_dataOut_bits_114),
    .io_dataOut_bits_115(vgg_io_dataOut_bits_115),
    .io_dataOut_bits_116(vgg_io_dataOut_bits_116),
    .io_dataOut_bits_117(vgg_io_dataOut_bits_117),
    .io_dataOut_bits_118(vgg_io_dataOut_bits_118),
    .io_dataOut_bits_119(vgg_io_dataOut_bits_119),
    .io_dataOut_bits_120(vgg_io_dataOut_bits_120),
    .io_dataOut_bits_121(vgg_io_dataOut_bits_121),
    .io_dataOut_bits_122(vgg_io_dataOut_bits_122),
    .io_dataOut_bits_123(vgg_io_dataOut_bits_123),
    .io_dataOut_bits_124(vgg_io_dataOut_bits_124),
    .io_dataOut_bits_125(vgg_io_dataOut_bits_125),
    .io_dataOut_bits_126(vgg_io_dataOut_bits_126),
    .io_dataOut_bits_127(vgg_io_dataOut_bits_127),
    .io_dataOut_bits_128(vgg_io_dataOut_bits_128),
    .io_dataOut_bits_129(vgg_io_dataOut_bits_129),
    .io_dataOut_bits_130(vgg_io_dataOut_bits_130),
    .io_dataOut_bits_131(vgg_io_dataOut_bits_131),
    .io_dataOut_bits_132(vgg_io_dataOut_bits_132),
    .io_dataOut_bits_133(vgg_io_dataOut_bits_133),
    .io_dataOut_bits_134(vgg_io_dataOut_bits_134),
    .io_dataOut_bits_135(vgg_io_dataOut_bits_135),
    .io_dataOut_bits_136(vgg_io_dataOut_bits_136),
    .io_dataOut_bits_137(vgg_io_dataOut_bits_137),
    .io_dataOut_bits_138(vgg_io_dataOut_bits_138),
    .io_dataOut_bits_139(vgg_io_dataOut_bits_139),
    .io_dataOut_bits_140(vgg_io_dataOut_bits_140),
    .io_dataOut_bits_141(vgg_io_dataOut_bits_141),
    .io_dataOut_bits_142(vgg_io_dataOut_bits_142),
    .io_dataOut_bits_143(vgg_io_dataOut_bits_143),
    .io_dataOut_bits_144(vgg_io_dataOut_bits_144),
    .io_dataOut_bits_145(vgg_io_dataOut_bits_145),
    .io_dataOut_bits_146(vgg_io_dataOut_bits_146),
    .io_dataOut_bits_147(vgg_io_dataOut_bits_147),
    .io_dataOut_bits_148(vgg_io_dataOut_bits_148),
    .io_dataOut_bits_149(vgg_io_dataOut_bits_149),
    .io_dataOut_bits_150(vgg_io_dataOut_bits_150),
    .io_dataOut_bits_151(vgg_io_dataOut_bits_151),
    .io_dataOut_bits_152(vgg_io_dataOut_bits_152),
    .io_dataOut_bits_153(vgg_io_dataOut_bits_153),
    .io_dataOut_bits_154(vgg_io_dataOut_bits_154),
    .io_dataOut_bits_155(vgg_io_dataOut_bits_155),
    .io_dataOut_bits_156(vgg_io_dataOut_bits_156),
    .io_dataOut_bits_157(vgg_io_dataOut_bits_157),
    .io_dataOut_bits_158(vgg_io_dataOut_bits_158),
    .io_dataOut_bits_159(vgg_io_dataOut_bits_159),
    .io_dataOut_bits_160(vgg_io_dataOut_bits_160),
    .io_dataOut_bits_161(vgg_io_dataOut_bits_161),
    .io_dataOut_bits_162(vgg_io_dataOut_bits_162),
    .io_dataOut_bits_163(vgg_io_dataOut_bits_163),
    .io_dataOut_bits_164(vgg_io_dataOut_bits_164),
    .io_dataOut_bits_165(vgg_io_dataOut_bits_165),
    .io_dataOut_bits_166(vgg_io_dataOut_bits_166),
    .io_dataOut_bits_167(vgg_io_dataOut_bits_167),
    .io_dataOut_bits_168(vgg_io_dataOut_bits_168),
    .io_dataOut_bits_169(vgg_io_dataOut_bits_169),
    .io_dataOut_bits_170(vgg_io_dataOut_bits_170),
    .io_dataOut_bits_171(vgg_io_dataOut_bits_171),
    .io_dataOut_bits_172(vgg_io_dataOut_bits_172),
    .io_dataOut_bits_173(vgg_io_dataOut_bits_173),
    .io_dataOut_bits_174(vgg_io_dataOut_bits_174),
    .io_dataOut_bits_175(vgg_io_dataOut_bits_175),
    .io_dataOut_bits_176(vgg_io_dataOut_bits_176),
    .io_dataOut_bits_177(vgg_io_dataOut_bits_177),
    .io_dataOut_bits_178(vgg_io_dataOut_bits_178),
    .io_dataOut_bits_179(vgg_io_dataOut_bits_179),
    .io_dataOut_bits_180(vgg_io_dataOut_bits_180),
    .io_dataOut_bits_181(vgg_io_dataOut_bits_181),
    .io_dataOut_bits_182(vgg_io_dataOut_bits_182),
    .io_dataOut_bits_183(vgg_io_dataOut_bits_183),
    .io_dataOut_bits_184(vgg_io_dataOut_bits_184),
    .io_dataOut_bits_185(vgg_io_dataOut_bits_185),
    .io_dataOut_bits_186(vgg_io_dataOut_bits_186),
    .io_dataOut_bits_187(vgg_io_dataOut_bits_187),
    .io_dataOut_bits_188(vgg_io_dataOut_bits_188),
    .io_dataOut_bits_189(vgg_io_dataOut_bits_189),
    .io_dataOut_bits_190(vgg_io_dataOut_bits_190),
    .io_dataOut_bits_191(vgg_io_dataOut_bits_191),
    .io_dataOut_bits_192(vgg_io_dataOut_bits_192),
    .io_dataOut_bits_193(vgg_io_dataOut_bits_193),
    .io_dataOut_bits_194(vgg_io_dataOut_bits_194),
    .io_dataOut_bits_195(vgg_io_dataOut_bits_195),
    .io_dataOut_bits_196(vgg_io_dataOut_bits_196),
    .io_dataOut_bits_197(vgg_io_dataOut_bits_197),
    .io_dataOut_bits_198(vgg_io_dataOut_bits_198),
    .io_dataOut_bits_199(vgg_io_dataOut_bits_199),
    .io_dataOut_bits_200(vgg_io_dataOut_bits_200),
    .io_dataOut_bits_201(vgg_io_dataOut_bits_201),
    .io_dataOut_bits_202(vgg_io_dataOut_bits_202),
    .io_dataOut_bits_203(vgg_io_dataOut_bits_203),
    .io_dataOut_bits_204(vgg_io_dataOut_bits_204),
    .io_dataOut_bits_205(vgg_io_dataOut_bits_205),
    .io_dataOut_bits_206(vgg_io_dataOut_bits_206),
    .io_dataOut_bits_207(vgg_io_dataOut_bits_207),
    .io_dataOut_bits_208(vgg_io_dataOut_bits_208),
    .io_dataOut_bits_209(vgg_io_dataOut_bits_209),
    .io_dataOut_bits_210(vgg_io_dataOut_bits_210),
    .io_dataOut_bits_211(vgg_io_dataOut_bits_211),
    .io_dataOut_bits_212(vgg_io_dataOut_bits_212),
    .io_dataOut_bits_213(vgg_io_dataOut_bits_213),
    .io_dataOut_bits_214(vgg_io_dataOut_bits_214),
    .io_dataOut_bits_215(vgg_io_dataOut_bits_215),
    .io_dataOut_bits_216(vgg_io_dataOut_bits_216),
    .io_dataOut_bits_217(vgg_io_dataOut_bits_217),
    .io_dataOut_bits_218(vgg_io_dataOut_bits_218),
    .io_dataOut_bits_219(vgg_io_dataOut_bits_219),
    .io_dataOut_bits_220(vgg_io_dataOut_bits_220),
    .io_dataOut_bits_221(vgg_io_dataOut_bits_221),
    .io_dataOut_bits_222(vgg_io_dataOut_bits_222),
    .io_dataOut_bits_223(vgg_io_dataOut_bits_223),
    .io_dataOut_bits_224(vgg_io_dataOut_bits_224),
    .io_dataOut_bits_225(vgg_io_dataOut_bits_225),
    .io_dataOut_bits_226(vgg_io_dataOut_bits_226),
    .io_dataOut_bits_227(vgg_io_dataOut_bits_227),
    .io_dataOut_bits_228(vgg_io_dataOut_bits_228),
    .io_dataOut_bits_229(vgg_io_dataOut_bits_229),
    .io_dataOut_bits_230(vgg_io_dataOut_bits_230),
    .io_dataOut_bits_231(vgg_io_dataOut_bits_231),
    .io_dataOut_bits_232(vgg_io_dataOut_bits_232),
    .io_dataOut_bits_233(vgg_io_dataOut_bits_233),
    .io_dataOut_bits_234(vgg_io_dataOut_bits_234),
    .io_dataOut_bits_235(vgg_io_dataOut_bits_235),
    .io_dataOut_bits_236(vgg_io_dataOut_bits_236),
    .io_dataOut_bits_237(vgg_io_dataOut_bits_237),
    .io_dataOut_bits_238(vgg_io_dataOut_bits_238),
    .io_dataOut_bits_239(vgg_io_dataOut_bits_239),
    .io_dataOut_bits_240(vgg_io_dataOut_bits_240),
    .io_dataOut_bits_241(vgg_io_dataOut_bits_241),
    .io_dataOut_bits_242(vgg_io_dataOut_bits_242),
    .io_dataOut_bits_243(vgg_io_dataOut_bits_243),
    .io_dataOut_bits_244(vgg_io_dataOut_bits_244),
    .io_dataOut_bits_245(vgg_io_dataOut_bits_245),
    .io_dataOut_bits_246(vgg_io_dataOut_bits_246),
    .io_dataOut_bits_247(vgg_io_dataOut_bits_247),
    .io_dataOut_bits_248(vgg_io_dataOut_bits_248),
    .io_dataOut_bits_249(vgg_io_dataOut_bits_249),
    .io_dataOut_bits_250(vgg_io_dataOut_bits_250),
    .io_dataOut_bits_251(vgg_io_dataOut_bits_251),
    .io_dataOut_bits_252(vgg_io_dataOut_bits_252),
    .io_dataOut_bits_253(vgg_io_dataOut_bits_253),
    .io_dataOut_bits_254(vgg_io_dataOut_bits_254),
    .io_dataOut_bits_255(vgg_io_dataOut_bits_255)
  );
  Queue_4096 queueIOOut ( // @[Decoupled.scala 289:19]
    .clock(queueIOOut_clock),
    .reset(queueIOOut_reset),
    .io_enq_ready(queueIOOut_io_enq_ready),
    .io_enq_valid(queueIOOut_io_enq_valid),
    .io_enq_bits(queueIOOut_io_enq_bits),
    .io_deq_ready(queueIOOut_io_deq_ready),
    .io_deq_valid(queueIOOut_io_deq_valid),
    .io_deq_bits(queueIOOut_io_deq_bits)
  );
  MuxLayer muxLyr ( // @[AWSVggWrapper.scala 66:22]
    .clock(muxLyr_clock),
    .reset(muxLyr_reset),
    .io_dataIn_ready(muxLyr_io_dataIn_ready),
    .io_dataIn_valid(muxLyr_io_dataIn_valid),
    .io_dataIn_bits_0(muxLyr_io_dataIn_bits_0),
    .io_dataIn_bits_1(muxLyr_io_dataIn_bits_1),
    .io_dataIn_bits_2(muxLyr_io_dataIn_bits_2),
    .io_dataIn_bits_3(muxLyr_io_dataIn_bits_3),
    .io_dataIn_bits_4(muxLyr_io_dataIn_bits_4),
    .io_dataIn_bits_5(muxLyr_io_dataIn_bits_5),
    .io_dataIn_bits_6(muxLyr_io_dataIn_bits_6),
    .io_dataIn_bits_7(muxLyr_io_dataIn_bits_7),
    .io_dataIn_bits_8(muxLyr_io_dataIn_bits_8),
    .io_dataIn_bits_9(muxLyr_io_dataIn_bits_9),
    .io_dataIn_bits_10(muxLyr_io_dataIn_bits_10),
    .io_dataIn_bits_11(muxLyr_io_dataIn_bits_11),
    .io_dataIn_bits_12(muxLyr_io_dataIn_bits_12),
    .io_dataIn_bits_13(muxLyr_io_dataIn_bits_13),
    .io_dataIn_bits_14(muxLyr_io_dataIn_bits_14),
    .io_dataIn_bits_15(muxLyr_io_dataIn_bits_15),
    .io_dataIn_bits_16(muxLyr_io_dataIn_bits_16),
    .io_dataIn_bits_17(muxLyr_io_dataIn_bits_17),
    .io_dataIn_bits_18(muxLyr_io_dataIn_bits_18),
    .io_dataIn_bits_19(muxLyr_io_dataIn_bits_19),
    .io_dataIn_bits_20(muxLyr_io_dataIn_bits_20),
    .io_dataIn_bits_21(muxLyr_io_dataIn_bits_21),
    .io_dataIn_bits_22(muxLyr_io_dataIn_bits_22),
    .io_dataIn_bits_23(muxLyr_io_dataIn_bits_23),
    .io_dataIn_bits_24(muxLyr_io_dataIn_bits_24),
    .io_dataIn_bits_25(muxLyr_io_dataIn_bits_25),
    .io_dataIn_bits_26(muxLyr_io_dataIn_bits_26),
    .io_dataIn_bits_27(muxLyr_io_dataIn_bits_27),
    .io_dataIn_bits_28(muxLyr_io_dataIn_bits_28),
    .io_dataIn_bits_29(muxLyr_io_dataIn_bits_29),
    .io_dataIn_bits_30(muxLyr_io_dataIn_bits_30),
    .io_dataIn_bits_31(muxLyr_io_dataIn_bits_31),
    .io_dataIn_bits_32(muxLyr_io_dataIn_bits_32),
    .io_dataIn_bits_33(muxLyr_io_dataIn_bits_33),
    .io_dataIn_bits_34(muxLyr_io_dataIn_bits_34),
    .io_dataIn_bits_35(muxLyr_io_dataIn_bits_35),
    .io_dataIn_bits_36(muxLyr_io_dataIn_bits_36),
    .io_dataIn_bits_37(muxLyr_io_dataIn_bits_37),
    .io_dataIn_bits_38(muxLyr_io_dataIn_bits_38),
    .io_dataIn_bits_39(muxLyr_io_dataIn_bits_39),
    .io_dataIn_bits_40(muxLyr_io_dataIn_bits_40),
    .io_dataIn_bits_41(muxLyr_io_dataIn_bits_41),
    .io_dataIn_bits_42(muxLyr_io_dataIn_bits_42),
    .io_dataIn_bits_43(muxLyr_io_dataIn_bits_43),
    .io_dataIn_bits_44(muxLyr_io_dataIn_bits_44),
    .io_dataIn_bits_45(muxLyr_io_dataIn_bits_45),
    .io_dataIn_bits_46(muxLyr_io_dataIn_bits_46),
    .io_dataIn_bits_47(muxLyr_io_dataIn_bits_47),
    .io_dataIn_bits_48(muxLyr_io_dataIn_bits_48),
    .io_dataIn_bits_49(muxLyr_io_dataIn_bits_49),
    .io_dataIn_bits_50(muxLyr_io_dataIn_bits_50),
    .io_dataIn_bits_51(muxLyr_io_dataIn_bits_51),
    .io_dataIn_bits_52(muxLyr_io_dataIn_bits_52),
    .io_dataIn_bits_53(muxLyr_io_dataIn_bits_53),
    .io_dataIn_bits_54(muxLyr_io_dataIn_bits_54),
    .io_dataIn_bits_55(muxLyr_io_dataIn_bits_55),
    .io_dataIn_bits_56(muxLyr_io_dataIn_bits_56),
    .io_dataIn_bits_57(muxLyr_io_dataIn_bits_57),
    .io_dataIn_bits_58(muxLyr_io_dataIn_bits_58),
    .io_dataIn_bits_59(muxLyr_io_dataIn_bits_59),
    .io_dataIn_bits_60(muxLyr_io_dataIn_bits_60),
    .io_dataIn_bits_61(muxLyr_io_dataIn_bits_61),
    .io_dataIn_bits_62(muxLyr_io_dataIn_bits_62),
    .io_dataIn_bits_63(muxLyr_io_dataIn_bits_63),
    .io_dataIn_bits_64(muxLyr_io_dataIn_bits_64),
    .io_dataIn_bits_65(muxLyr_io_dataIn_bits_65),
    .io_dataIn_bits_66(muxLyr_io_dataIn_bits_66),
    .io_dataIn_bits_67(muxLyr_io_dataIn_bits_67),
    .io_dataIn_bits_68(muxLyr_io_dataIn_bits_68),
    .io_dataIn_bits_69(muxLyr_io_dataIn_bits_69),
    .io_dataIn_bits_70(muxLyr_io_dataIn_bits_70),
    .io_dataIn_bits_71(muxLyr_io_dataIn_bits_71),
    .io_dataIn_bits_72(muxLyr_io_dataIn_bits_72),
    .io_dataIn_bits_73(muxLyr_io_dataIn_bits_73),
    .io_dataIn_bits_74(muxLyr_io_dataIn_bits_74),
    .io_dataIn_bits_75(muxLyr_io_dataIn_bits_75),
    .io_dataIn_bits_76(muxLyr_io_dataIn_bits_76),
    .io_dataIn_bits_77(muxLyr_io_dataIn_bits_77),
    .io_dataIn_bits_78(muxLyr_io_dataIn_bits_78),
    .io_dataIn_bits_79(muxLyr_io_dataIn_bits_79),
    .io_dataIn_bits_80(muxLyr_io_dataIn_bits_80),
    .io_dataIn_bits_81(muxLyr_io_dataIn_bits_81),
    .io_dataIn_bits_82(muxLyr_io_dataIn_bits_82),
    .io_dataIn_bits_83(muxLyr_io_dataIn_bits_83),
    .io_dataIn_bits_84(muxLyr_io_dataIn_bits_84),
    .io_dataIn_bits_85(muxLyr_io_dataIn_bits_85),
    .io_dataIn_bits_86(muxLyr_io_dataIn_bits_86),
    .io_dataIn_bits_87(muxLyr_io_dataIn_bits_87),
    .io_dataIn_bits_88(muxLyr_io_dataIn_bits_88),
    .io_dataIn_bits_89(muxLyr_io_dataIn_bits_89),
    .io_dataIn_bits_90(muxLyr_io_dataIn_bits_90),
    .io_dataIn_bits_91(muxLyr_io_dataIn_bits_91),
    .io_dataIn_bits_92(muxLyr_io_dataIn_bits_92),
    .io_dataIn_bits_93(muxLyr_io_dataIn_bits_93),
    .io_dataIn_bits_94(muxLyr_io_dataIn_bits_94),
    .io_dataIn_bits_95(muxLyr_io_dataIn_bits_95),
    .io_dataIn_bits_96(muxLyr_io_dataIn_bits_96),
    .io_dataIn_bits_97(muxLyr_io_dataIn_bits_97),
    .io_dataIn_bits_98(muxLyr_io_dataIn_bits_98),
    .io_dataIn_bits_99(muxLyr_io_dataIn_bits_99),
    .io_dataIn_bits_100(muxLyr_io_dataIn_bits_100),
    .io_dataIn_bits_101(muxLyr_io_dataIn_bits_101),
    .io_dataIn_bits_102(muxLyr_io_dataIn_bits_102),
    .io_dataIn_bits_103(muxLyr_io_dataIn_bits_103),
    .io_dataIn_bits_104(muxLyr_io_dataIn_bits_104),
    .io_dataIn_bits_105(muxLyr_io_dataIn_bits_105),
    .io_dataIn_bits_106(muxLyr_io_dataIn_bits_106),
    .io_dataIn_bits_107(muxLyr_io_dataIn_bits_107),
    .io_dataIn_bits_108(muxLyr_io_dataIn_bits_108),
    .io_dataIn_bits_109(muxLyr_io_dataIn_bits_109),
    .io_dataIn_bits_110(muxLyr_io_dataIn_bits_110),
    .io_dataIn_bits_111(muxLyr_io_dataIn_bits_111),
    .io_dataIn_bits_112(muxLyr_io_dataIn_bits_112),
    .io_dataIn_bits_113(muxLyr_io_dataIn_bits_113),
    .io_dataIn_bits_114(muxLyr_io_dataIn_bits_114),
    .io_dataIn_bits_115(muxLyr_io_dataIn_bits_115),
    .io_dataIn_bits_116(muxLyr_io_dataIn_bits_116),
    .io_dataIn_bits_117(muxLyr_io_dataIn_bits_117),
    .io_dataIn_bits_118(muxLyr_io_dataIn_bits_118),
    .io_dataIn_bits_119(muxLyr_io_dataIn_bits_119),
    .io_dataIn_bits_120(muxLyr_io_dataIn_bits_120),
    .io_dataIn_bits_121(muxLyr_io_dataIn_bits_121),
    .io_dataIn_bits_122(muxLyr_io_dataIn_bits_122),
    .io_dataIn_bits_123(muxLyr_io_dataIn_bits_123),
    .io_dataIn_bits_124(muxLyr_io_dataIn_bits_124),
    .io_dataIn_bits_125(muxLyr_io_dataIn_bits_125),
    .io_dataIn_bits_126(muxLyr_io_dataIn_bits_126),
    .io_dataIn_bits_127(muxLyr_io_dataIn_bits_127),
    .io_dataIn_bits_128(muxLyr_io_dataIn_bits_128),
    .io_dataIn_bits_129(muxLyr_io_dataIn_bits_129),
    .io_dataIn_bits_130(muxLyr_io_dataIn_bits_130),
    .io_dataIn_bits_131(muxLyr_io_dataIn_bits_131),
    .io_dataIn_bits_132(muxLyr_io_dataIn_bits_132),
    .io_dataIn_bits_133(muxLyr_io_dataIn_bits_133),
    .io_dataIn_bits_134(muxLyr_io_dataIn_bits_134),
    .io_dataIn_bits_135(muxLyr_io_dataIn_bits_135),
    .io_dataIn_bits_136(muxLyr_io_dataIn_bits_136),
    .io_dataIn_bits_137(muxLyr_io_dataIn_bits_137),
    .io_dataIn_bits_138(muxLyr_io_dataIn_bits_138),
    .io_dataIn_bits_139(muxLyr_io_dataIn_bits_139),
    .io_dataIn_bits_140(muxLyr_io_dataIn_bits_140),
    .io_dataIn_bits_141(muxLyr_io_dataIn_bits_141),
    .io_dataIn_bits_142(muxLyr_io_dataIn_bits_142),
    .io_dataIn_bits_143(muxLyr_io_dataIn_bits_143),
    .io_dataIn_bits_144(muxLyr_io_dataIn_bits_144),
    .io_dataIn_bits_145(muxLyr_io_dataIn_bits_145),
    .io_dataIn_bits_146(muxLyr_io_dataIn_bits_146),
    .io_dataIn_bits_147(muxLyr_io_dataIn_bits_147),
    .io_dataIn_bits_148(muxLyr_io_dataIn_bits_148),
    .io_dataIn_bits_149(muxLyr_io_dataIn_bits_149),
    .io_dataIn_bits_150(muxLyr_io_dataIn_bits_150),
    .io_dataIn_bits_151(muxLyr_io_dataIn_bits_151),
    .io_dataIn_bits_152(muxLyr_io_dataIn_bits_152),
    .io_dataIn_bits_153(muxLyr_io_dataIn_bits_153),
    .io_dataIn_bits_154(muxLyr_io_dataIn_bits_154),
    .io_dataIn_bits_155(muxLyr_io_dataIn_bits_155),
    .io_dataIn_bits_156(muxLyr_io_dataIn_bits_156),
    .io_dataIn_bits_157(muxLyr_io_dataIn_bits_157),
    .io_dataIn_bits_158(muxLyr_io_dataIn_bits_158),
    .io_dataIn_bits_159(muxLyr_io_dataIn_bits_159),
    .io_dataIn_bits_160(muxLyr_io_dataIn_bits_160),
    .io_dataIn_bits_161(muxLyr_io_dataIn_bits_161),
    .io_dataIn_bits_162(muxLyr_io_dataIn_bits_162),
    .io_dataIn_bits_163(muxLyr_io_dataIn_bits_163),
    .io_dataIn_bits_164(muxLyr_io_dataIn_bits_164),
    .io_dataIn_bits_165(muxLyr_io_dataIn_bits_165),
    .io_dataIn_bits_166(muxLyr_io_dataIn_bits_166),
    .io_dataIn_bits_167(muxLyr_io_dataIn_bits_167),
    .io_dataIn_bits_168(muxLyr_io_dataIn_bits_168),
    .io_dataIn_bits_169(muxLyr_io_dataIn_bits_169),
    .io_dataIn_bits_170(muxLyr_io_dataIn_bits_170),
    .io_dataIn_bits_171(muxLyr_io_dataIn_bits_171),
    .io_dataIn_bits_172(muxLyr_io_dataIn_bits_172),
    .io_dataIn_bits_173(muxLyr_io_dataIn_bits_173),
    .io_dataIn_bits_174(muxLyr_io_dataIn_bits_174),
    .io_dataIn_bits_175(muxLyr_io_dataIn_bits_175),
    .io_dataIn_bits_176(muxLyr_io_dataIn_bits_176),
    .io_dataIn_bits_177(muxLyr_io_dataIn_bits_177),
    .io_dataIn_bits_178(muxLyr_io_dataIn_bits_178),
    .io_dataIn_bits_179(muxLyr_io_dataIn_bits_179),
    .io_dataIn_bits_180(muxLyr_io_dataIn_bits_180),
    .io_dataIn_bits_181(muxLyr_io_dataIn_bits_181),
    .io_dataIn_bits_182(muxLyr_io_dataIn_bits_182),
    .io_dataIn_bits_183(muxLyr_io_dataIn_bits_183),
    .io_dataIn_bits_184(muxLyr_io_dataIn_bits_184),
    .io_dataIn_bits_185(muxLyr_io_dataIn_bits_185),
    .io_dataIn_bits_186(muxLyr_io_dataIn_bits_186),
    .io_dataIn_bits_187(muxLyr_io_dataIn_bits_187),
    .io_dataIn_bits_188(muxLyr_io_dataIn_bits_188),
    .io_dataIn_bits_189(muxLyr_io_dataIn_bits_189),
    .io_dataIn_bits_190(muxLyr_io_dataIn_bits_190),
    .io_dataIn_bits_191(muxLyr_io_dataIn_bits_191),
    .io_dataIn_bits_192(muxLyr_io_dataIn_bits_192),
    .io_dataIn_bits_193(muxLyr_io_dataIn_bits_193),
    .io_dataIn_bits_194(muxLyr_io_dataIn_bits_194),
    .io_dataIn_bits_195(muxLyr_io_dataIn_bits_195),
    .io_dataIn_bits_196(muxLyr_io_dataIn_bits_196),
    .io_dataIn_bits_197(muxLyr_io_dataIn_bits_197),
    .io_dataIn_bits_198(muxLyr_io_dataIn_bits_198),
    .io_dataIn_bits_199(muxLyr_io_dataIn_bits_199),
    .io_dataIn_bits_200(muxLyr_io_dataIn_bits_200),
    .io_dataIn_bits_201(muxLyr_io_dataIn_bits_201),
    .io_dataIn_bits_202(muxLyr_io_dataIn_bits_202),
    .io_dataIn_bits_203(muxLyr_io_dataIn_bits_203),
    .io_dataIn_bits_204(muxLyr_io_dataIn_bits_204),
    .io_dataIn_bits_205(muxLyr_io_dataIn_bits_205),
    .io_dataIn_bits_206(muxLyr_io_dataIn_bits_206),
    .io_dataIn_bits_207(muxLyr_io_dataIn_bits_207),
    .io_dataIn_bits_208(muxLyr_io_dataIn_bits_208),
    .io_dataIn_bits_209(muxLyr_io_dataIn_bits_209),
    .io_dataIn_bits_210(muxLyr_io_dataIn_bits_210),
    .io_dataIn_bits_211(muxLyr_io_dataIn_bits_211),
    .io_dataIn_bits_212(muxLyr_io_dataIn_bits_212),
    .io_dataIn_bits_213(muxLyr_io_dataIn_bits_213),
    .io_dataIn_bits_214(muxLyr_io_dataIn_bits_214),
    .io_dataIn_bits_215(muxLyr_io_dataIn_bits_215),
    .io_dataIn_bits_216(muxLyr_io_dataIn_bits_216),
    .io_dataIn_bits_217(muxLyr_io_dataIn_bits_217),
    .io_dataIn_bits_218(muxLyr_io_dataIn_bits_218),
    .io_dataIn_bits_219(muxLyr_io_dataIn_bits_219),
    .io_dataIn_bits_220(muxLyr_io_dataIn_bits_220),
    .io_dataIn_bits_221(muxLyr_io_dataIn_bits_221),
    .io_dataIn_bits_222(muxLyr_io_dataIn_bits_222),
    .io_dataIn_bits_223(muxLyr_io_dataIn_bits_223),
    .io_dataIn_bits_224(muxLyr_io_dataIn_bits_224),
    .io_dataIn_bits_225(muxLyr_io_dataIn_bits_225),
    .io_dataIn_bits_226(muxLyr_io_dataIn_bits_226),
    .io_dataIn_bits_227(muxLyr_io_dataIn_bits_227),
    .io_dataIn_bits_228(muxLyr_io_dataIn_bits_228),
    .io_dataIn_bits_229(muxLyr_io_dataIn_bits_229),
    .io_dataIn_bits_230(muxLyr_io_dataIn_bits_230),
    .io_dataIn_bits_231(muxLyr_io_dataIn_bits_231),
    .io_dataIn_bits_232(muxLyr_io_dataIn_bits_232),
    .io_dataIn_bits_233(muxLyr_io_dataIn_bits_233),
    .io_dataIn_bits_234(muxLyr_io_dataIn_bits_234),
    .io_dataIn_bits_235(muxLyr_io_dataIn_bits_235),
    .io_dataIn_bits_236(muxLyr_io_dataIn_bits_236),
    .io_dataIn_bits_237(muxLyr_io_dataIn_bits_237),
    .io_dataIn_bits_238(muxLyr_io_dataIn_bits_238),
    .io_dataIn_bits_239(muxLyr_io_dataIn_bits_239),
    .io_dataIn_bits_240(muxLyr_io_dataIn_bits_240),
    .io_dataIn_bits_241(muxLyr_io_dataIn_bits_241),
    .io_dataIn_bits_242(muxLyr_io_dataIn_bits_242),
    .io_dataIn_bits_243(muxLyr_io_dataIn_bits_243),
    .io_dataIn_bits_244(muxLyr_io_dataIn_bits_244),
    .io_dataIn_bits_245(muxLyr_io_dataIn_bits_245),
    .io_dataIn_bits_246(muxLyr_io_dataIn_bits_246),
    .io_dataIn_bits_247(muxLyr_io_dataIn_bits_247),
    .io_dataIn_bits_248(muxLyr_io_dataIn_bits_248),
    .io_dataIn_bits_249(muxLyr_io_dataIn_bits_249),
    .io_dataIn_bits_250(muxLyr_io_dataIn_bits_250),
    .io_dataIn_bits_251(muxLyr_io_dataIn_bits_251),
    .io_dataIn_bits_252(muxLyr_io_dataIn_bits_252),
    .io_dataIn_bits_253(muxLyr_io_dataIn_bits_253),
    .io_dataIn_bits_254(muxLyr_io_dataIn_bits_254),
    .io_dataIn_bits_255(muxLyr_io_dataIn_bits_255),
    .io_dataOut_valid(muxLyr_io_dataOut_valid),
    .io_dataOut_bits_0(muxLyr_io_dataOut_bits_0),
    .io_dataOut_bits_1(muxLyr_io_dataOut_bits_1),
    .io_dataOut_bits_2(muxLyr_io_dataOut_bits_2),
    .io_dataOut_bits_3(muxLyr_io_dataOut_bits_3)
  );
  DenseLayer dense ( // @[AWSVggWrapper.scala 75:21]
    .clock(dense_clock),
    .reset(dense_reset),
    .io_dataIn_valid(dense_io_dataIn_valid),
    .io_dataIn_bits_0(dense_io_dataIn_bits_0),
    .io_dataIn_bits_1(dense_io_dataIn_bits_1),
    .io_dataIn_bits_2(dense_io_dataIn_bits_2),
    .io_dataIn_bits_3(dense_io_dataIn_bits_3),
    .io_dataOut_valid(dense_io_dataOut_valid),
    .io_dataOut_bits_0(dense_io_dataOut_bits_0),
    .io_dataOut_bits_1(dense_io_dataOut_bits_1),
    .io_dataOut_bits_2(dense_io_dataOut_bits_2),
    .io_dataOut_bits_3(dense_io_dataOut_bits_3),
    .io_dataOut_bits_4(dense_io_dataOut_bits_4),
    .io_dataOut_bits_5(dense_io_dataOut_bits_5),
    .io_dataOut_bits_6(dense_io_dataOut_bits_6),
    .io_dataOut_bits_7(dense_io_dataOut_bits_7),
    .io_dataOut_bits_8(dense_io_dataOut_bits_8),
    .io_dataOut_bits_9(dense_io_dataOut_bits_9),
    .io_dataOut_bits_10(dense_io_dataOut_bits_10),
    .io_dataOut_bits_11(dense_io_dataOut_bits_11),
    .io_dataOut_bits_12(dense_io_dataOut_bits_12),
    .io_dataOut_bits_13(dense_io_dataOut_bits_13),
    .io_dataOut_bits_14(dense_io_dataOut_bits_14),
    .io_dataOut_bits_15(dense_io_dataOut_bits_15),
    .io_dataOut_bits_16(dense_io_dataOut_bits_16),
    .io_dataOut_bits_17(dense_io_dataOut_bits_17),
    .io_dataOut_bits_18(dense_io_dataOut_bits_18),
    .io_dataOut_bits_19(dense_io_dataOut_bits_19),
    .io_dataOut_bits_20(dense_io_dataOut_bits_20),
    .io_dataOut_bits_21(dense_io_dataOut_bits_21),
    .io_dataOut_bits_22(dense_io_dataOut_bits_22),
    .io_dataOut_bits_23(dense_io_dataOut_bits_23),
    .io_dataOut_bits_24(dense_io_dataOut_bits_24),
    .io_dataOut_bits_25(dense_io_dataOut_bits_25),
    .io_dataOut_bits_26(dense_io_dataOut_bits_26),
    .io_dataOut_bits_27(dense_io_dataOut_bits_27),
    .io_dataOut_bits_28(dense_io_dataOut_bits_28),
    .io_dataOut_bits_29(dense_io_dataOut_bits_29),
    .io_dataOut_bits_30(dense_io_dataOut_bits_30),
    .io_dataOut_bits_31(dense_io_dataOut_bits_31),
    .io_dataOut_bits_32(dense_io_dataOut_bits_32),
    .io_dataOut_bits_33(dense_io_dataOut_bits_33),
    .io_dataOut_bits_34(dense_io_dataOut_bits_34),
    .io_dataOut_bits_35(dense_io_dataOut_bits_35),
    .io_dataOut_bits_36(dense_io_dataOut_bits_36),
    .io_dataOut_bits_37(dense_io_dataOut_bits_37),
    .io_dataOut_bits_38(dense_io_dataOut_bits_38),
    .io_dataOut_bits_39(dense_io_dataOut_bits_39),
    .io_dataOut_bits_40(dense_io_dataOut_bits_40),
    .io_dataOut_bits_41(dense_io_dataOut_bits_41),
    .io_dataOut_bits_42(dense_io_dataOut_bits_42),
    .io_dataOut_bits_43(dense_io_dataOut_bits_43),
    .io_dataOut_bits_44(dense_io_dataOut_bits_44),
    .io_dataOut_bits_45(dense_io_dataOut_bits_45),
    .io_dataOut_bits_46(dense_io_dataOut_bits_46),
    .io_dataOut_bits_47(dense_io_dataOut_bits_47),
    .io_dataOut_bits_48(dense_io_dataOut_bits_48),
    .io_dataOut_bits_49(dense_io_dataOut_bits_49),
    .io_dataOut_bits_50(dense_io_dataOut_bits_50),
    .io_dataOut_bits_51(dense_io_dataOut_bits_51),
    .io_dataOut_bits_52(dense_io_dataOut_bits_52),
    .io_dataOut_bits_53(dense_io_dataOut_bits_53),
    .io_dataOut_bits_54(dense_io_dataOut_bits_54),
    .io_dataOut_bits_55(dense_io_dataOut_bits_55),
    .io_dataOut_bits_56(dense_io_dataOut_bits_56),
    .io_dataOut_bits_57(dense_io_dataOut_bits_57),
    .io_dataOut_bits_58(dense_io_dataOut_bits_58),
    .io_dataOut_bits_59(dense_io_dataOut_bits_59),
    .io_dataOut_bits_60(dense_io_dataOut_bits_60),
    .io_dataOut_bits_61(dense_io_dataOut_bits_61),
    .io_dataOut_bits_62(dense_io_dataOut_bits_62),
    .io_dataOut_bits_63(dense_io_dataOut_bits_63),
    .io_dataOut_bits_64(dense_io_dataOut_bits_64),
    .io_dataOut_bits_65(dense_io_dataOut_bits_65),
    .io_dataOut_bits_66(dense_io_dataOut_bits_66),
    .io_dataOut_bits_67(dense_io_dataOut_bits_67),
    .io_dataOut_bits_68(dense_io_dataOut_bits_68),
    .io_dataOut_bits_69(dense_io_dataOut_bits_69),
    .io_dataOut_bits_70(dense_io_dataOut_bits_70),
    .io_dataOut_bits_71(dense_io_dataOut_bits_71),
    .io_dataOut_bits_72(dense_io_dataOut_bits_72),
    .io_dataOut_bits_73(dense_io_dataOut_bits_73),
    .io_dataOut_bits_74(dense_io_dataOut_bits_74),
    .io_dataOut_bits_75(dense_io_dataOut_bits_75),
    .io_dataOut_bits_76(dense_io_dataOut_bits_76),
    .io_dataOut_bits_77(dense_io_dataOut_bits_77),
    .io_dataOut_bits_78(dense_io_dataOut_bits_78),
    .io_dataOut_bits_79(dense_io_dataOut_bits_79),
    .io_dataOut_bits_80(dense_io_dataOut_bits_80),
    .io_dataOut_bits_81(dense_io_dataOut_bits_81),
    .io_dataOut_bits_82(dense_io_dataOut_bits_82),
    .io_dataOut_bits_83(dense_io_dataOut_bits_83),
    .io_dataOut_bits_84(dense_io_dataOut_bits_84),
    .io_dataOut_bits_85(dense_io_dataOut_bits_85),
    .io_dataOut_bits_86(dense_io_dataOut_bits_86),
    .io_dataOut_bits_87(dense_io_dataOut_bits_87),
    .io_dataOut_bits_88(dense_io_dataOut_bits_88),
    .io_dataOut_bits_89(dense_io_dataOut_bits_89),
    .io_dataOut_bits_90(dense_io_dataOut_bits_90),
    .io_dataOut_bits_91(dense_io_dataOut_bits_91),
    .io_dataOut_bits_92(dense_io_dataOut_bits_92),
    .io_dataOut_bits_93(dense_io_dataOut_bits_93),
    .io_dataOut_bits_94(dense_io_dataOut_bits_94),
    .io_dataOut_bits_95(dense_io_dataOut_bits_95),
    .io_dataOut_bits_96(dense_io_dataOut_bits_96),
    .io_dataOut_bits_97(dense_io_dataOut_bits_97),
    .io_dataOut_bits_98(dense_io_dataOut_bits_98),
    .io_dataOut_bits_99(dense_io_dataOut_bits_99),
    .io_dataOut_bits_100(dense_io_dataOut_bits_100),
    .io_dataOut_bits_101(dense_io_dataOut_bits_101),
    .io_dataOut_bits_102(dense_io_dataOut_bits_102),
    .io_dataOut_bits_103(dense_io_dataOut_bits_103),
    .io_dataOut_bits_104(dense_io_dataOut_bits_104),
    .io_dataOut_bits_105(dense_io_dataOut_bits_105),
    .io_dataOut_bits_106(dense_io_dataOut_bits_106),
    .io_dataOut_bits_107(dense_io_dataOut_bits_107),
    .io_dataOut_bits_108(dense_io_dataOut_bits_108),
    .io_dataOut_bits_109(dense_io_dataOut_bits_109),
    .io_dataOut_bits_110(dense_io_dataOut_bits_110),
    .io_dataOut_bits_111(dense_io_dataOut_bits_111),
    .io_dataOut_bits_112(dense_io_dataOut_bits_112),
    .io_dataOut_bits_113(dense_io_dataOut_bits_113),
    .io_dataOut_bits_114(dense_io_dataOut_bits_114),
    .io_dataOut_bits_115(dense_io_dataOut_bits_115),
    .io_dataOut_bits_116(dense_io_dataOut_bits_116),
    .io_dataOut_bits_117(dense_io_dataOut_bits_117),
    .io_dataOut_bits_118(dense_io_dataOut_bits_118),
    .io_dataOut_bits_119(dense_io_dataOut_bits_119),
    .io_dataOut_bits_120(dense_io_dataOut_bits_120),
    .io_dataOut_bits_121(dense_io_dataOut_bits_121),
    .io_dataOut_bits_122(dense_io_dataOut_bits_122),
    .io_dataOut_bits_123(dense_io_dataOut_bits_123),
    .io_dataOut_bits_124(dense_io_dataOut_bits_124),
    .io_dataOut_bits_125(dense_io_dataOut_bits_125),
    .io_dataOut_bits_126(dense_io_dataOut_bits_126),
    .io_dataOut_bits_127(dense_io_dataOut_bits_127)
  );
  SSILayerOut muxLyr_2 ( // @[AWSVggWrapper.scala 79:24]
    .clock(muxLyr_2_clock),
    .reset(muxLyr_2_reset),
    .io_dataIn_valid(muxLyr_2_io_dataIn_valid),
    .io_dataIn_bits_0(muxLyr_2_io_dataIn_bits_0),
    .io_dataIn_bits_1(muxLyr_2_io_dataIn_bits_1),
    .io_dataIn_bits_2(muxLyr_2_io_dataIn_bits_2),
    .io_dataIn_bits_3(muxLyr_2_io_dataIn_bits_3),
    .io_dataIn_bits_4(muxLyr_2_io_dataIn_bits_4),
    .io_dataIn_bits_5(muxLyr_2_io_dataIn_bits_5),
    .io_dataIn_bits_6(muxLyr_2_io_dataIn_bits_6),
    .io_dataIn_bits_7(muxLyr_2_io_dataIn_bits_7),
    .io_dataIn_bits_8(muxLyr_2_io_dataIn_bits_8),
    .io_dataIn_bits_9(muxLyr_2_io_dataIn_bits_9),
    .io_dataIn_bits_10(muxLyr_2_io_dataIn_bits_10),
    .io_dataIn_bits_11(muxLyr_2_io_dataIn_bits_11),
    .io_dataIn_bits_12(muxLyr_2_io_dataIn_bits_12),
    .io_dataIn_bits_13(muxLyr_2_io_dataIn_bits_13),
    .io_dataIn_bits_14(muxLyr_2_io_dataIn_bits_14),
    .io_dataIn_bits_15(muxLyr_2_io_dataIn_bits_15),
    .io_dataIn_bits_16(muxLyr_2_io_dataIn_bits_16),
    .io_dataIn_bits_17(muxLyr_2_io_dataIn_bits_17),
    .io_dataIn_bits_18(muxLyr_2_io_dataIn_bits_18),
    .io_dataIn_bits_19(muxLyr_2_io_dataIn_bits_19),
    .io_dataIn_bits_20(muxLyr_2_io_dataIn_bits_20),
    .io_dataIn_bits_21(muxLyr_2_io_dataIn_bits_21),
    .io_dataIn_bits_22(muxLyr_2_io_dataIn_bits_22),
    .io_dataIn_bits_23(muxLyr_2_io_dataIn_bits_23),
    .io_dataIn_bits_24(muxLyr_2_io_dataIn_bits_24),
    .io_dataIn_bits_25(muxLyr_2_io_dataIn_bits_25),
    .io_dataIn_bits_26(muxLyr_2_io_dataIn_bits_26),
    .io_dataIn_bits_27(muxLyr_2_io_dataIn_bits_27),
    .io_dataIn_bits_28(muxLyr_2_io_dataIn_bits_28),
    .io_dataIn_bits_29(muxLyr_2_io_dataIn_bits_29),
    .io_dataIn_bits_30(muxLyr_2_io_dataIn_bits_30),
    .io_dataIn_bits_31(muxLyr_2_io_dataIn_bits_31),
    .io_dataIn_bits_32(muxLyr_2_io_dataIn_bits_32),
    .io_dataIn_bits_33(muxLyr_2_io_dataIn_bits_33),
    .io_dataIn_bits_34(muxLyr_2_io_dataIn_bits_34),
    .io_dataIn_bits_35(muxLyr_2_io_dataIn_bits_35),
    .io_dataIn_bits_36(muxLyr_2_io_dataIn_bits_36),
    .io_dataIn_bits_37(muxLyr_2_io_dataIn_bits_37),
    .io_dataIn_bits_38(muxLyr_2_io_dataIn_bits_38),
    .io_dataIn_bits_39(muxLyr_2_io_dataIn_bits_39),
    .io_dataIn_bits_40(muxLyr_2_io_dataIn_bits_40),
    .io_dataIn_bits_41(muxLyr_2_io_dataIn_bits_41),
    .io_dataIn_bits_42(muxLyr_2_io_dataIn_bits_42),
    .io_dataIn_bits_43(muxLyr_2_io_dataIn_bits_43),
    .io_dataIn_bits_44(muxLyr_2_io_dataIn_bits_44),
    .io_dataIn_bits_45(muxLyr_2_io_dataIn_bits_45),
    .io_dataIn_bits_46(muxLyr_2_io_dataIn_bits_46),
    .io_dataIn_bits_47(muxLyr_2_io_dataIn_bits_47),
    .io_dataIn_bits_48(muxLyr_2_io_dataIn_bits_48),
    .io_dataIn_bits_49(muxLyr_2_io_dataIn_bits_49),
    .io_dataIn_bits_50(muxLyr_2_io_dataIn_bits_50),
    .io_dataIn_bits_51(muxLyr_2_io_dataIn_bits_51),
    .io_dataIn_bits_52(muxLyr_2_io_dataIn_bits_52),
    .io_dataIn_bits_53(muxLyr_2_io_dataIn_bits_53),
    .io_dataIn_bits_54(muxLyr_2_io_dataIn_bits_54),
    .io_dataIn_bits_55(muxLyr_2_io_dataIn_bits_55),
    .io_dataIn_bits_56(muxLyr_2_io_dataIn_bits_56),
    .io_dataIn_bits_57(muxLyr_2_io_dataIn_bits_57),
    .io_dataIn_bits_58(muxLyr_2_io_dataIn_bits_58),
    .io_dataIn_bits_59(muxLyr_2_io_dataIn_bits_59),
    .io_dataIn_bits_60(muxLyr_2_io_dataIn_bits_60),
    .io_dataIn_bits_61(muxLyr_2_io_dataIn_bits_61),
    .io_dataIn_bits_62(muxLyr_2_io_dataIn_bits_62),
    .io_dataIn_bits_63(muxLyr_2_io_dataIn_bits_63),
    .io_dataIn_bits_64(muxLyr_2_io_dataIn_bits_64),
    .io_dataIn_bits_65(muxLyr_2_io_dataIn_bits_65),
    .io_dataIn_bits_66(muxLyr_2_io_dataIn_bits_66),
    .io_dataIn_bits_67(muxLyr_2_io_dataIn_bits_67),
    .io_dataIn_bits_68(muxLyr_2_io_dataIn_bits_68),
    .io_dataIn_bits_69(muxLyr_2_io_dataIn_bits_69),
    .io_dataIn_bits_70(muxLyr_2_io_dataIn_bits_70),
    .io_dataIn_bits_71(muxLyr_2_io_dataIn_bits_71),
    .io_dataIn_bits_72(muxLyr_2_io_dataIn_bits_72),
    .io_dataIn_bits_73(muxLyr_2_io_dataIn_bits_73),
    .io_dataIn_bits_74(muxLyr_2_io_dataIn_bits_74),
    .io_dataIn_bits_75(muxLyr_2_io_dataIn_bits_75),
    .io_dataIn_bits_76(muxLyr_2_io_dataIn_bits_76),
    .io_dataIn_bits_77(muxLyr_2_io_dataIn_bits_77),
    .io_dataIn_bits_78(muxLyr_2_io_dataIn_bits_78),
    .io_dataIn_bits_79(muxLyr_2_io_dataIn_bits_79),
    .io_dataIn_bits_80(muxLyr_2_io_dataIn_bits_80),
    .io_dataIn_bits_81(muxLyr_2_io_dataIn_bits_81),
    .io_dataIn_bits_82(muxLyr_2_io_dataIn_bits_82),
    .io_dataIn_bits_83(muxLyr_2_io_dataIn_bits_83),
    .io_dataIn_bits_84(muxLyr_2_io_dataIn_bits_84),
    .io_dataIn_bits_85(muxLyr_2_io_dataIn_bits_85),
    .io_dataIn_bits_86(muxLyr_2_io_dataIn_bits_86),
    .io_dataIn_bits_87(muxLyr_2_io_dataIn_bits_87),
    .io_dataIn_bits_88(muxLyr_2_io_dataIn_bits_88),
    .io_dataIn_bits_89(muxLyr_2_io_dataIn_bits_89),
    .io_dataIn_bits_90(muxLyr_2_io_dataIn_bits_90),
    .io_dataIn_bits_91(muxLyr_2_io_dataIn_bits_91),
    .io_dataIn_bits_92(muxLyr_2_io_dataIn_bits_92),
    .io_dataIn_bits_93(muxLyr_2_io_dataIn_bits_93),
    .io_dataIn_bits_94(muxLyr_2_io_dataIn_bits_94),
    .io_dataIn_bits_95(muxLyr_2_io_dataIn_bits_95),
    .io_dataIn_bits_96(muxLyr_2_io_dataIn_bits_96),
    .io_dataIn_bits_97(muxLyr_2_io_dataIn_bits_97),
    .io_dataIn_bits_98(muxLyr_2_io_dataIn_bits_98),
    .io_dataIn_bits_99(muxLyr_2_io_dataIn_bits_99),
    .io_dataIn_bits_100(muxLyr_2_io_dataIn_bits_100),
    .io_dataIn_bits_101(muxLyr_2_io_dataIn_bits_101),
    .io_dataIn_bits_102(muxLyr_2_io_dataIn_bits_102),
    .io_dataIn_bits_103(muxLyr_2_io_dataIn_bits_103),
    .io_dataIn_bits_104(muxLyr_2_io_dataIn_bits_104),
    .io_dataIn_bits_105(muxLyr_2_io_dataIn_bits_105),
    .io_dataIn_bits_106(muxLyr_2_io_dataIn_bits_106),
    .io_dataIn_bits_107(muxLyr_2_io_dataIn_bits_107),
    .io_dataIn_bits_108(muxLyr_2_io_dataIn_bits_108),
    .io_dataIn_bits_109(muxLyr_2_io_dataIn_bits_109),
    .io_dataIn_bits_110(muxLyr_2_io_dataIn_bits_110),
    .io_dataIn_bits_111(muxLyr_2_io_dataIn_bits_111),
    .io_dataIn_bits_112(muxLyr_2_io_dataIn_bits_112),
    .io_dataIn_bits_113(muxLyr_2_io_dataIn_bits_113),
    .io_dataIn_bits_114(muxLyr_2_io_dataIn_bits_114),
    .io_dataIn_bits_115(muxLyr_2_io_dataIn_bits_115),
    .io_dataIn_bits_116(muxLyr_2_io_dataIn_bits_116),
    .io_dataIn_bits_117(muxLyr_2_io_dataIn_bits_117),
    .io_dataIn_bits_118(muxLyr_2_io_dataIn_bits_118),
    .io_dataIn_bits_119(muxLyr_2_io_dataIn_bits_119),
    .io_dataIn_bits_120(muxLyr_2_io_dataIn_bits_120),
    .io_dataIn_bits_121(muxLyr_2_io_dataIn_bits_121),
    .io_dataIn_bits_122(muxLyr_2_io_dataIn_bits_122),
    .io_dataIn_bits_123(muxLyr_2_io_dataIn_bits_123),
    .io_dataIn_bits_124(muxLyr_2_io_dataIn_bits_124),
    .io_dataIn_bits_125(muxLyr_2_io_dataIn_bits_125),
    .io_dataIn_bits_126(muxLyr_2_io_dataIn_bits_126),
    .io_dataIn_bits_127(muxLyr_2_io_dataIn_bits_127),
    .io_dataOut_valid(muxLyr_2_io_dataOut_valid),
    .io_dataOut_bits_0(muxLyr_2_io_dataOut_bits_0)
  );
  DenseScale scale ( // @[AWSVggWrapper.scala 92:21]
    .clock(scale_clock),
    .reset(scale_reset),
    .io_dataIn_valid(scale_io_dataIn_valid),
    .io_dataIn_bits_0(scale_io_dataIn_bits_0),
    .io_dataOut_valid(scale_io_dataOut_valid),
    .io_dataOut_bits_0(scale_io_dataOut_bits_0)
  );
  DenseLayer_1 dense_2 ( // @[AWSVggWrapper.scala 99:23]
    .clock(dense_2_clock),
    .reset(dense_2_reset),
    .io_dataIn_valid(dense_2_io_dataIn_valid),
    .io_dataIn_bits_0(dense_2_io_dataIn_bits_0),
    .io_dataOut_valid(dense_2_io_dataOut_valid),
    .io_dataOut_bits_0(dense_2_io_dataOut_bits_0),
    .io_dataOut_bits_1(dense_2_io_dataOut_bits_1),
    .io_dataOut_bits_2(dense_2_io_dataOut_bits_2),
    .io_dataOut_bits_3(dense_2_io_dataOut_bits_3),
    .io_dataOut_bits_4(dense_2_io_dataOut_bits_4),
    .io_dataOut_bits_5(dense_2_io_dataOut_bits_5),
    .io_dataOut_bits_6(dense_2_io_dataOut_bits_6),
    .io_dataOut_bits_7(dense_2_io_dataOut_bits_7),
    .io_dataOut_bits_8(dense_2_io_dataOut_bits_8),
    .io_dataOut_bits_9(dense_2_io_dataOut_bits_9)
  );
  assign _T_35 = $unsigned(vgg_io_dataOut_bits_0); // @[AWSVggWrapper.scala 53:79]
  assign _T_36 = $unsigned(vgg_io_dataOut_bits_1); // @[AWSVggWrapper.scala 53:79]
  assign _T_37 = $unsigned(vgg_io_dataOut_bits_2); // @[AWSVggWrapper.scala 53:79]
  assign _T_38 = $unsigned(vgg_io_dataOut_bits_3); // @[AWSVggWrapper.scala 53:79]
  assign _T_39 = $unsigned(vgg_io_dataOut_bits_4); // @[AWSVggWrapper.scala 53:79]
  assign _T_40 = $unsigned(vgg_io_dataOut_bits_5); // @[AWSVggWrapper.scala 53:79]
  assign _T_41 = $unsigned(vgg_io_dataOut_bits_6); // @[AWSVggWrapper.scala 53:79]
  assign _T_42 = $unsigned(vgg_io_dataOut_bits_7); // @[AWSVggWrapper.scala 53:79]
  assign _T_43 = $unsigned(vgg_io_dataOut_bits_8); // @[AWSVggWrapper.scala 53:79]
  assign _T_44 = $unsigned(vgg_io_dataOut_bits_9); // @[AWSVggWrapper.scala 53:79]
  assign _T_45 = $unsigned(vgg_io_dataOut_bits_10); // @[AWSVggWrapper.scala 53:79]
  assign _T_46 = $unsigned(vgg_io_dataOut_bits_11); // @[AWSVggWrapper.scala 53:79]
  assign _T_47 = $unsigned(vgg_io_dataOut_bits_12); // @[AWSVggWrapper.scala 53:79]
  assign _T_48 = $unsigned(vgg_io_dataOut_bits_13); // @[AWSVggWrapper.scala 53:79]
  assign _T_49 = $unsigned(vgg_io_dataOut_bits_14); // @[AWSVggWrapper.scala 53:79]
  assign _T_50 = $unsigned(vgg_io_dataOut_bits_15); // @[AWSVggWrapper.scala 53:79]
  assign _T_51 = $unsigned(vgg_io_dataOut_bits_16); // @[AWSVggWrapper.scala 53:79]
  assign _T_52 = $unsigned(vgg_io_dataOut_bits_17); // @[AWSVggWrapper.scala 53:79]
  assign _T_53 = $unsigned(vgg_io_dataOut_bits_18); // @[AWSVggWrapper.scala 53:79]
  assign _T_54 = $unsigned(vgg_io_dataOut_bits_19); // @[AWSVggWrapper.scala 53:79]
  assign _T_55 = $unsigned(vgg_io_dataOut_bits_20); // @[AWSVggWrapper.scala 53:79]
  assign _T_56 = $unsigned(vgg_io_dataOut_bits_21); // @[AWSVggWrapper.scala 53:79]
  assign _T_57 = $unsigned(vgg_io_dataOut_bits_22); // @[AWSVggWrapper.scala 53:79]
  assign _T_58 = $unsigned(vgg_io_dataOut_bits_23); // @[AWSVggWrapper.scala 53:79]
  assign _T_59 = $unsigned(vgg_io_dataOut_bits_24); // @[AWSVggWrapper.scala 53:79]
  assign _T_60 = $unsigned(vgg_io_dataOut_bits_25); // @[AWSVggWrapper.scala 53:79]
  assign _T_61 = $unsigned(vgg_io_dataOut_bits_26); // @[AWSVggWrapper.scala 53:79]
  assign _T_62 = $unsigned(vgg_io_dataOut_bits_27); // @[AWSVggWrapper.scala 53:79]
  assign _T_63 = $unsigned(vgg_io_dataOut_bits_28); // @[AWSVggWrapper.scala 53:79]
  assign _T_64 = $unsigned(vgg_io_dataOut_bits_29); // @[AWSVggWrapper.scala 53:79]
  assign _T_65 = $unsigned(vgg_io_dataOut_bits_30); // @[AWSVggWrapper.scala 53:79]
  assign _T_66 = $unsigned(vgg_io_dataOut_bits_31); // @[AWSVggWrapper.scala 53:79]
  assign _T_67 = $unsigned(vgg_io_dataOut_bits_32); // @[AWSVggWrapper.scala 53:79]
  assign _T_68 = $unsigned(vgg_io_dataOut_bits_33); // @[AWSVggWrapper.scala 53:79]
  assign _T_69 = $unsigned(vgg_io_dataOut_bits_34); // @[AWSVggWrapper.scala 53:79]
  assign _T_70 = $unsigned(vgg_io_dataOut_bits_35); // @[AWSVggWrapper.scala 53:79]
  assign _T_71 = $unsigned(vgg_io_dataOut_bits_36); // @[AWSVggWrapper.scala 53:79]
  assign _T_72 = $unsigned(vgg_io_dataOut_bits_37); // @[AWSVggWrapper.scala 53:79]
  assign _T_73 = $unsigned(vgg_io_dataOut_bits_38); // @[AWSVggWrapper.scala 53:79]
  assign _T_74 = $unsigned(vgg_io_dataOut_bits_39); // @[AWSVggWrapper.scala 53:79]
  assign _T_75 = $unsigned(vgg_io_dataOut_bits_40); // @[AWSVggWrapper.scala 53:79]
  assign _T_76 = $unsigned(vgg_io_dataOut_bits_41); // @[AWSVggWrapper.scala 53:79]
  assign _T_77 = $unsigned(vgg_io_dataOut_bits_42); // @[AWSVggWrapper.scala 53:79]
  assign _T_78 = $unsigned(vgg_io_dataOut_bits_43); // @[AWSVggWrapper.scala 53:79]
  assign _T_79 = $unsigned(vgg_io_dataOut_bits_44); // @[AWSVggWrapper.scala 53:79]
  assign _T_80 = $unsigned(vgg_io_dataOut_bits_45); // @[AWSVggWrapper.scala 53:79]
  assign _T_81 = $unsigned(vgg_io_dataOut_bits_46); // @[AWSVggWrapper.scala 53:79]
  assign _T_82 = $unsigned(vgg_io_dataOut_bits_47); // @[AWSVggWrapper.scala 53:79]
  assign _T_83 = $unsigned(vgg_io_dataOut_bits_48); // @[AWSVggWrapper.scala 53:79]
  assign _T_84 = $unsigned(vgg_io_dataOut_bits_49); // @[AWSVggWrapper.scala 53:79]
  assign _T_85 = $unsigned(vgg_io_dataOut_bits_50); // @[AWSVggWrapper.scala 53:79]
  assign _T_86 = $unsigned(vgg_io_dataOut_bits_51); // @[AWSVggWrapper.scala 53:79]
  assign _T_87 = $unsigned(vgg_io_dataOut_bits_52); // @[AWSVggWrapper.scala 53:79]
  assign _T_88 = $unsigned(vgg_io_dataOut_bits_53); // @[AWSVggWrapper.scala 53:79]
  assign _T_89 = $unsigned(vgg_io_dataOut_bits_54); // @[AWSVggWrapper.scala 53:79]
  assign _T_90 = $unsigned(vgg_io_dataOut_bits_55); // @[AWSVggWrapper.scala 53:79]
  assign _T_91 = $unsigned(vgg_io_dataOut_bits_56); // @[AWSVggWrapper.scala 53:79]
  assign _T_92 = $unsigned(vgg_io_dataOut_bits_57); // @[AWSVggWrapper.scala 53:79]
  assign _T_93 = $unsigned(vgg_io_dataOut_bits_58); // @[AWSVggWrapper.scala 53:79]
  assign _T_94 = $unsigned(vgg_io_dataOut_bits_59); // @[AWSVggWrapper.scala 53:79]
  assign _T_95 = $unsigned(vgg_io_dataOut_bits_60); // @[AWSVggWrapper.scala 53:79]
  assign _T_96 = $unsigned(vgg_io_dataOut_bits_61); // @[AWSVggWrapper.scala 53:79]
  assign _T_97 = $unsigned(vgg_io_dataOut_bits_62); // @[AWSVggWrapper.scala 53:79]
  assign _T_98 = $unsigned(vgg_io_dataOut_bits_63); // @[AWSVggWrapper.scala 53:79]
  assign _T_99 = $unsigned(vgg_io_dataOut_bits_64); // @[AWSVggWrapper.scala 53:79]
  assign _T_100 = $unsigned(vgg_io_dataOut_bits_65); // @[AWSVggWrapper.scala 53:79]
  assign _T_101 = $unsigned(vgg_io_dataOut_bits_66); // @[AWSVggWrapper.scala 53:79]
  assign _T_102 = $unsigned(vgg_io_dataOut_bits_67); // @[AWSVggWrapper.scala 53:79]
  assign _T_103 = $unsigned(vgg_io_dataOut_bits_68); // @[AWSVggWrapper.scala 53:79]
  assign _T_104 = $unsigned(vgg_io_dataOut_bits_69); // @[AWSVggWrapper.scala 53:79]
  assign _T_105 = $unsigned(vgg_io_dataOut_bits_70); // @[AWSVggWrapper.scala 53:79]
  assign _T_106 = $unsigned(vgg_io_dataOut_bits_71); // @[AWSVggWrapper.scala 53:79]
  assign _T_107 = $unsigned(vgg_io_dataOut_bits_72); // @[AWSVggWrapper.scala 53:79]
  assign _T_108 = $unsigned(vgg_io_dataOut_bits_73); // @[AWSVggWrapper.scala 53:79]
  assign _T_109 = $unsigned(vgg_io_dataOut_bits_74); // @[AWSVggWrapper.scala 53:79]
  assign _T_110 = $unsigned(vgg_io_dataOut_bits_75); // @[AWSVggWrapper.scala 53:79]
  assign _T_111 = $unsigned(vgg_io_dataOut_bits_76); // @[AWSVggWrapper.scala 53:79]
  assign _T_112 = $unsigned(vgg_io_dataOut_bits_77); // @[AWSVggWrapper.scala 53:79]
  assign _T_113 = $unsigned(vgg_io_dataOut_bits_78); // @[AWSVggWrapper.scala 53:79]
  assign _T_114 = $unsigned(vgg_io_dataOut_bits_79); // @[AWSVggWrapper.scala 53:79]
  assign _T_115 = $unsigned(vgg_io_dataOut_bits_80); // @[AWSVggWrapper.scala 53:79]
  assign _T_116 = $unsigned(vgg_io_dataOut_bits_81); // @[AWSVggWrapper.scala 53:79]
  assign _T_117 = $unsigned(vgg_io_dataOut_bits_82); // @[AWSVggWrapper.scala 53:79]
  assign _T_118 = $unsigned(vgg_io_dataOut_bits_83); // @[AWSVggWrapper.scala 53:79]
  assign _T_119 = $unsigned(vgg_io_dataOut_bits_84); // @[AWSVggWrapper.scala 53:79]
  assign _T_120 = $unsigned(vgg_io_dataOut_bits_85); // @[AWSVggWrapper.scala 53:79]
  assign _T_121 = $unsigned(vgg_io_dataOut_bits_86); // @[AWSVggWrapper.scala 53:79]
  assign _T_122 = $unsigned(vgg_io_dataOut_bits_87); // @[AWSVggWrapper.scala 53:79]
  assign _T_123 = $unsigned(vgg_io_dataOut_bits_88); // @[AWSVggWrapper.scala 53:79]
  assign _T_124 = $unsigned(vgg_io_dataOut_bits_89); // @[AWSVggWrapper.scala 53:79]
  assign _T_125 = $unsigned(vgg_io_dataOut_bits_90); // @[AWSVggWrapper.scala 53:79]
  assign _T_126 = $unsigned(vgg_io_dataOut_bits_91); // @[AWSVggWrapper.scala 53:79]
  assign _T_127 = $unsigned(vgg_io_dataOut_bits_92); // @[AWSVggWrapper.scala 53:79]
  assign _T_128 = $unsigned(vgg_io_dataOut_bits_93); // @[AWSVggWrapper.scala 53:79]
  assign _T_129 = $unsigned(vgg_io_dataOut_bits_94); // @[AWSVggWrapper.scala 53:79]
  assign _T_130 = $unsigned(vgg_io_dataOut_bits_95); // @[AWSVggWrapper.scala 53:79]
  assign _T_131 = $unsigned(vgg_io_dataOut_bits_96); // @[AWSVggWrapper.scala 53:79]
  assign _T_132 = $unsigned(vgg_io_dataOut_bits_97); // @[AWSVggWrapper.scala 53:79]
  assign _T_133 = $unsigned(vgg_io_dataOut_bits_98); // @[AWSVggWrapper.scala 53:79]
  assign _T_134 = $unsigned(vgg_io_dataOut_bits_99); // @[AWSVggWrapper.scala 53:79]
  assign _T_135 = $unsigned(vgg_io_dataOut_bits_100); // @[AWSVggWrapper.scala 53:79]
  assign _T_136 = $unsigned(vgg_io_dataOut_bits_101); // @[AWSVggWrapper.scala 53:79]
  assign _T_137 = $unsigned(vgg_io_dataOut_bits_102); // @[AWSVggWrapper.scala 53:79]
  assign _T_138 = $unsigned(vgg_io_dataOut_bits_103); // @[AWSVggWrapper.scala 53:79]
  assign _T_139 = $unsigned(vgg_io_dataOut_bits_104); // @[AWSVggWrapper.scala 53:79]
  assign _T_140 = $unsigned(vgg_io_dataOut_bits_105); // @[AWSVggWrapper.scala 53:79]
  assign _T_141 = $unsigned(vgg_io_dataOut_bits_106); // @[AWSVggWrapper.scala 53:79]
  assign _T_142 = $unsigned(vgg_io_dataOut_bits_107); // @[AWSVggWrapper.scala 53:79]
  assign _T_143 = $unsigned(vgg_io_dataOut_bits_108); // @[AWSVggWrapper.scala 53:79]
  assign _T_144 = $unsigned(vgg_io_dataOut_bits_109); // @[AWSVggWrapper.scala 53:79]
  assign _T_145 = $unsigned(vgg_io_dataOut_bits_110); // @[AWSVggWrapper.scala 53:79]
  assign _T_146 = $unsigned(vgg_io_dataOut_bits_111); // @[AWSVggWrapper.scala 53:79]
  assign _T_147 = $unsigned(vgg_io_dataOut_bits_112); // @[AWSVggWrapper.scala 53:79]
  assign _T_148 = $unsigned(vgg_io_dataOut_bits_113); // @[AWSVggWrapper.scala 53:79]
  assign _T_149 = $unsigned(vgg_io_dataOut_bits_114); // @[AWSVggWrapper.scala 53:79]
  assign _T_150 = $unsigned(vgg_io_dataOut_bits_115); // @[AWSVggWrapper.scala 53:79]
  assign _T_151 = $unsigned(vgg_io_dataOut_bits_116); // @[AWSVggWrapper.scala 53:79]
  assign _T_152 = $unsigned(vgg_io_dataOut_bits_117); // @[AWSVggWrapper.scala 53:79]
  assign _T_153 = $unsigned(vgg_io_dataOut_bits_118); // @[AWSVggWrapper.scala 53:79]
  assign _T_154 = $unsigned(vgg_io_dataOut_bits_119); // @[AWSVggWrapper.scala 53:79]
  assign _T_155 = $unsigned(vgg_io_dataOut_bits_120); // @[AWSVggWrapper.scala 53:79]
  assign _T_156 = $unsigned(vgg_io_dataOut_bits_121); // @[AWSVggWrapper.scala 53:79]
  assign _T_157 = $unsigned(vgg_io_dataOut_bits_122); // @[AWSVggWrapper.scala 53:79]
  assign _T_158 = $unsigned(vgg_io_dataOut_bits_123); // @[AWSVggWrapper.scala 53:79]
  assign _T_159 = $unsigned(vgg_io_dataOut_bits_124); // @[AWSVggWrapper.scala 53:79]
  assign _T_160 = $unsigned(vgg_io_dataOut_bits_125); // @[AWSVggWrapper.scala 53:79]
  assign _T_161 = $unsigned(vgg_io_dataOut_bits_126); // @[AWSVggWrapper.scala 53:79]
  assign _T_162 = $unsigned(vgg_io_dataOut_bits_127); // @[AWSVggWrapper.scala 53:79]
  assign _T_163 = $unsigned(vgg_io_dataOut_bits_128); // @[AWSVggWrapper.scala 53:79]
  assign _T_164 = $unsigned(vgg_io_dataOut_bits_129); // @[AWSVggWrapper.scala 53:79]
  assign _T_165 = $unsigned(vgg_io_dataOut_bits_130); // @[AWSVggWrapper.scala 53:79]
  assign _T_166 = $unsigned(vgg_io_dataOut_bits_131); // @[AWSVggWrapper.scala 53:79]
  assign _T_167 = $unsigned(vgg_io_dataOut_bits_132); // @[AWSVggWrapper.scala 53:79]
  assign _T_168 = $unsigned(vgg_io_dataOut_bits_133); // @[AWSVggWrapper.scala 53:79]
  assign _T_169 = $unsigned(vgg_io_dataOut_bits_134); // @[AWSVggWrapper.scala 53:79]
  assign _T_170 = $unsigned(vgg_io_dataOut_bits_135); // @[AWSVggWrapper.scala 53:79]
  assign _T_171 = $unsigned(vgg_io_dataOut_bits_136); // @[AWSVggWrapper.scala 53:79]
  assign _T_172 = $unsigned(vgg_io_dataOut_bits_137); // @[AWSVggWrapper.scala 53:79]
  assign _T_173 = $unsigned(vgg_io_dataOut_bits_138); // @[AWSVggWrapper.scala 53:79]
  assign _T_174 = $unsigned(vgg_io_dataOut_bits_139); // @[AWSVggWrapper.scala 53:79]
  assign _T_175 = $unsigned(vgg_io_dataOut_bits_140); // @[AWSVggWrapper.scala 53:79]
  assign _T_176 = $unsigned(vgg_io_dataOut_bits_141); // @[AWSVggWrapper.scala 53:79]
  assign _T_177 = $unsigned(vgg_io_dataOut_bits_142); // @[AWSVggWrapper.scala 53:79]
  assign _T_178 = $unsigned(vgg_io_dataOut_bits_143); // @[AWSVggWrapper.scala 53:79]
  assign _T_179 = $unsigned(vgg_io_dataOut_bits_144); // @[AWSVggWrapper.scala 53:79]
  assign _T_180 = $unsigned(vgg_io_dataOut_bits_145); // @[AWSVggWrapper.scala 53:79]
  assign _T_181 = $unsigned(vgg_io_dataOut_bits_146); // @[AWSVggWrapper.scala 53:79]
  assign _T_182 = $unsigned(vgg_io_dataOut_bits_147); // @[AWSVggWrapper.scala 53:79]
  assign _T_183 = $unsigned(vgg_io_dataOut_bits_148); // @[AWSVggWrapper.scala 53:79]
  assign _T_184 = $unsigned(vgg_io_dataOut_bits_149); // @[AWSVggWrapper.scala 53:79]
  assign _T_185 = $unsigned(vgg_io_dataOut_bits_150); // @[AWSVggWrapper.scala 53:79]
  assign _T_186 = $unsigned(vgg_io_dataOut_bits_151); // @[AWSVggWrapper.scala 53:79]
  assign _T_187 = $unsigned(vgg_io_dataOut_bits_152); // @[AWSVggWrapper.scala 53:79]
  assign _T_188 = $unsigned(vgg_io_dataOut_bits_153); // @[AWSVggWrapper.scala 53:79]
  assign _T_189 = $unsigned(vgg_io_dataOut_bits_154); // @[AWSVggWrapper.scala 53:79]
  assign _T_190 = $unsigned(vgg_io_dataOut_bits_155); // @[AWSVggWrapper.scala 53:79]
  assign _T_191 = $unsigned(vgg_io_dataOut_bits_156); // @[AWSVggWrapper.scala 53:79]
  assign _T_192 = $unsigned(vgg_io_dataOut_bits_157); // @[AWSVggWrapper.scala 53:79]
  assign _T_193 = $unsigned(vgg_io_dataOut_bits_158); // @[AWSVggWrapper.scala 53:79]
  assign _T_194 = $unsigned(vgg_io_dataOut_bits_159); // @[AWSVggWrapper.scala 53:79]
  assign _T_195 = $unsigned(vgg_io_dataOut_bits_160); // @[AWSVggWrapper.scala 53:79]
  assign _T_196 = $unsigned(vgg_io_dataOut_bits_161); // @[AWSVggWrapper.scala 53:79]
  assign _T_197 = $unsigned(vgg_io_dataOut_bits_162); // @[AWSVggWrapper.scala 53:79]
  assign _T_198 = $unsigned(vgg_io_dataOut_bits_163); // @[AWSVggWrapper.scala 53:79]
  assign _T_199 = $unsigned(vgg_io_dataOut_bits_164); // @[AWSVggWrapper.scala 53:79]
  assign _T_200 = $unsigned(vgg_io_dataOut_bits_165); // @[AWSVggWrapper.scala 53:79]
  assign _T_201 = $unsigned(vgg_io_dataOut_bits_166); // @[AWSVggWrapper.scala 53:79]
  assign _T_202 = $unsigned(vgg_io_dataOut_bits_167); // @[AWSVggWrapper.scala 53:79]
  assign _T_203 = $unsigned(vgg_io_dataOut_bits_168); // @[AWSVggWrapper.scala 53:79]
  assign _T_204 = $unsigned(vgg_io_dataOut_bits_169); // @[AWSVggWrapper.scala 53:79]
  assign _T_205 = $unsigned(vgg_io_dataOut_bits_170); // @[AWSVggWrapper.scala 53:79]
  assign _T_206 = $unsigned(vgg_io_dataOut_bits_171); // @[AWSVggWrapper.scala 53:79]
  assign _T_207 = $unsigned(vgg_io_dataOut_bits_172); // @[AWSVggWrapper.scala 53:79]
  assign _T_208 = $unsigned(vgg_io_dataOut_bits_173); // @[AWSVggWrapper.scala 53:79]
  assign _T_209 = $unsigned(vgg_io_dataOut_bits_174); // @[AWSVggWrapper.scala 53:79]
  assign _T_210 = $unsigned(vgg_io_dataOut_bits_175); // @[AWSVggWrapper.scala 53:79]
  assign _T_211 = $unsigned(vgg_io_dataOut_bits_176); // @[AWSVggWrapper.scala 53:79]
  assign _T_212 = $unsigned(vgg_io_dataOut_bits_177); // @[AWSVggWrapper.scala 53:79]
  assign _T_213 = $unsigned(vgg_io_dataOut_bits_178); // @[AWSVggWrapper.scala 53:79]
  assign _T_214 = $unsigned(vgg_io_dataOut_bits_179); // @[AWSVggWrapper.scala 53:79]
  assign _T_215 = $unsigned(vgg_io_dataOut_bits_180); // @[AWSVggWrapper.scala 53:79]
  assign _T_216 = $unsigned(vgg_io_dataOut_bits_181); // @[AWSVggWrapper.scala 53:79]
  assign _T_217 = $unsigned(vgg_io_dataOut_bits_182); // @[AWSVggWrapper.scala 53:79]
  assign _T_218 = $unsigned(vgg_io_dataOut_bits_183); // @[AWSVggWrapper.scala 53:79]
  assign _T_219 = $unsigned(vgg_io_dataOut_bits_184); // @[AWSVggWrapper.scala 53:79]
  assign _T_220 = $unsigned(vgg_io_dataOut_bits_185); // @[AWSVggWrapper.scala 53:79]
  assign _T_221 = $unsigned(vgg_io_dataOut_bits_186); // @[AWSVggWrapper.scala 53:79]
  assign _T_222 = $unsigned(vgg_io_dataOut_bits_187); // @[AWSVggWrapper.scala 53:79]
  assign _T_223 = $unsigned(vgg_io_dataOut_bits_188); // @[AWSVggWrapper.scala 53:79]
  assign _T_224 = $unsigned(vgg_io_dataOut_bits_189); // @[AWSVggWrapper.scala 53:79]
  assign _T_225 = $unsigned(vgg_io_dataOut_bits_190); // @[AWSVggWrapper.scala 53:79]
  assign _T_226 = $unsigned(vgg_io_dataOut_bits_191); // @[AWSVggWrapper.scala 53:79]
  assign _T_227 = $unsigned(vgg_io_dataOut_bits_192); // @[AWSVggWrapper.scala 53:79]
  assign _T_228 = $unsigned(vgg_io_dataOut_bits_193); // @[AWSVggWrapper.scala 53:79]
  assign _T_229 = $unsigned(vgg_io_dataOut_bits_194); // @[AWSVggWrapper.scala 53:79]
  assign _T_230 = $unsigned(vgg_io_dataOut_bits_195); // @[AWSVggWrapper.scala 53:79]
  assign _T_231 = $unsigned(vgg_io_dataOut_bits_196); // @[AWSVggWrapper.scala 53:79]
  assign _T_232 = $unsigned(vgg_io_dataOut_bits_197); // @[AWSVggWrapper.scala 53:79]
  assign _T_233 = $unsigned(vgg_io_dataOut_bits_198); // @[AWSVggWrapper.scala 53:79]
  assign _T_234 = $unsigned(vgg_io_dataOut_bits_199); // @[AWSVggWrapper.scala 53:79]
  assign _T_235 = $unsigned(vgg_io_dataOut_bits_200); // @[AWSVggWrapper.scala 53:79]
  assign _T_236 = $unsigned(vgg_io_dataOut_bits_201); // @[AWSVggWrapper.scala 53:79]
  assign _T_237 = $unsigned(vgg_io_dataOut_bits_202); // @[AWSVggWrapper.scala 53:79]
  assign _T_238 = $unsigned(vgg_io_dataOut_bits_203); // @[AWSVggWrapper.scala 53:79]
  assign _T_239 = $unsigned(vgg_io_dataOut_bits_204); // @[AWSVggWrapper.scala 53:79]
  assign _T_240 = $unsigned(vgg_io_dataOut_bits_205); // @[AWSVggWrapper.scala 53:79]
  assign _T_241 = $unsigned(vgg_io_dataOut_bits_206); // @[AWSVggWrapper.scala 53:79]
  assign _T_242 = $unsigned(vgg_io_dataOut_bits_207); // @[AWSVggWrapper.scala 53:79]
  assign _T_243 = $unsigned(vgg_io_dataOut_bits_208); // @[AWSVggWrapper.scala 53:79]
  assign _T_244 = $unsigned(vgg_io_dataOut_bits_209); // @[AWSVggWrapper.scala 53:79]
  assign _T_245 = $unsigned(vgg_io_dataOut_bits_210); // @[AWSVggWrapper.scala 53:79]
  assign _T_246 = $unsigned(vgg_io_dataOut_bits_211); // @[AWSVggWrapper.scala 53:79]
  assign _T_247 = $unsigned(vgg_io_dataOut_bits_212); // @[AWSVggWrapper.scala 53:79]
  assign _T_248 = $unsigned(vgg_io_dataOut_bits_213); // @[AWSVggWrapper.scala 53:79]
  assign _T_249 = $unsigned(vgg_io_dataOut_bits_214); // @[AWSVggWrapper.scala 53:79]
  assign _T_250 = $unsigned(vgg_io_dataOut_bits_215); // @[AWSVggWrapper.scala 53:79]
  assign _T_251 = $unsigned(vgg_io_dataOut_bits_216); // @[AWSVggWrapper.scala 53:79]
  assign _T_252 = $unsigned(vgg_io_dataOut_bits_217); // @[AWSVggWrapper.scala 53:79]
  assign _T_253 = $unsigned(vgg_io_dataOut_bits_218); // @[AWSVggWrapper.scala 53:79]
  assign _T_254 = $unsigned(vgg_io_dataOut_bits_219); // @[AWSVggWrapper.scala 53:79]
  assign _T_255 = $unsigned(vgg_io_dataOut_bits_220); // @[AWSVggWrapper.scala 53:79]
  assign _T_256 = $unsigned(vgg_io_dataOut_bits_221); // @[AWSVggWrapper.scala 53:79]
  assign _T_257 = $unsigned(vgg_io_dataOut_bits_222); // @[AWSVggWrapper.scala 53:79]
  assign _T_258 = $unsigned(vgg_io_dataOut_bits_223); // @[AWSVggWrapper.scala 53:79]
  assign _T_259 = $unsigned(vgg_io_dataOut_bits_224); // @[AWSVggWrapper.scala 53:79]
  assign _T_260 = $unsigned(vgg_io_dataOut_bits_225); // @[AWSVggWrapper.scala 53:79]
  assign _T_261 = $unsigned(vgg_io_dataOut_bits_226); // @[AWSVggWrapper.scala 53:79]
  assign _T_262 = $unsigned(vgg_io_dataOut_bits_227); // @[AWSVggWrapper.scala 53:79]
  assign _T_263 = $unsigned(vgg_io_dataOut_bits_228); // @[AWSVggWrapper.scala 53:79]
  assign _T_264 = $unsigned(vgg_io_dataOut_bits_229); // @[AWSVggWrapper.scala 53:79]
  assign _T_265 = $unsigned(vgg_io_dataOut_bits_230); // @[AWSVggWrapper.scala 53:79]
  assign _T_266 = $unsigned(vgg_io_dataOut_bits_231); // @[AWSVggWrapper.scala 53:79]
  assign _T_267 = $unsigned(vgg_io_dataOut_bits_232); // @[AWSVggWrapper.scala 53:79]
  assign _T_268 = $unsigned(vgg_io_dataOut_bits_233); // @[AWSVggWrapper.scala 53:79]
  assign _T_269 = $unsigned(vgg_io_dataOut_bits_234); // @[AWSVggWrapper.scala 53:79]
  assign _T_270 = $unsigned(vgg_io_dataOut_bits_235); // @[AWSVggWrapper.scala 53:79]
  assign _T_271 = $unsigned(vgg_io_dataOut_bits_236); // @[AWSVggWrapper.scala 53:79]
  assign _T_272 = $unsigned(vgg_io_dataOut_bits_237); // @[AWSVggWrapper.scala 53:79]
  assign _T_273 = $unsigned(vgg_io_dataOut_bits_238); // @[AWSVggWrapper.scala 53:79]
  assign _T_274 = $unsigned(vgg_io_dataOut_bits_239); // @[AWSVggWrapper.scala 53:79]
  assign _T_275 = $unsigned(vgg_io_dataOut_bits_240); // @[AWSVggWrapper.scala 53:79]
  assign _T_276 = $unsigned(vgg_io_dataOut_bits_241); // @[AWSVggWrapper.scala 53:79]
  assign _T_277 = $unsigned(vgg_io_dataOut_bits_242); // @[AWSVggWrapper.scala 53:79]
  assign _T_278 = $unsigned(vgg_io_dataOut_bits_243); // @[AWSVggWrapper.scala 53:79]
  assign _T_279 = $unsigned(vgg_io_dataOut_bits_244); // @[AWSVggWrapper.scala 53:79]
  assign _T_280 = $unsigned(vgg_io_dataOut_bits_245); // @[AWSVggWrapper.scala 53:79]
  assign _T_281 = $unsigned(vgg_io_dataOut_bits_246); // @[AWSVggWrapper.scala 53:79]
  assign _T_282 = $unsigned(vgg_io_dataOut_bits_247); // @[AWSVggWrapper.scala 53:79]
  assign _T_283 = $unsigned(vgg_io_dataOut_bits_248); // @[AWSVggWrapper.scala 53:79]
  assign _T_284 = $unsigned(vgg_io_dataOut_bits_249); // @[AWSVggWrapper.scala 53:79]
  assign _T_285 = $unsigned(vgg_io_dataOut_bits_250); // @[AWSVggWrapper.scala 53:79]
  assign _T_286 = $unsigned(vgg_io_dataOut_bits_251); // @[AWSVggWrapper.scala 53:79]
  assign _T_287 = $unsigned(vgg_io_dataOut_bits_252); // @[AWSVggWrapper.scala 53:79]
  assign _T_288 = $unsigned(vgg_io_dataOut_bits_253); // @[AWSVggWrapper.scala 53:79]
  assign _T_289 = $unsigned(vgg_io_dataOut_bits_254); // @[AWSVggWrapper.scala 53:79]
  assign _T_290 = $unsigned(vgg_io_dataOut_bits_255); // @[AWSVggWrapper.scala 53:79]
  assign _T_291 = {_T_35,_T_36}; // @[AWSVggWrapper.scala 53:94]
  assign _T_292 = {_T_291,_T_37}; // @[AWSVggWrapper.scala 53:94]
  assign _T_293 = {_T_292,_T_38}; // @[AWSVggWrapper.scala 53:94]
  assign _T_294 = {_T_293,_T_39}; // @[AWSVggWrapper.scala 53:94]
  assign _T_295 = {_T_294,_T_40}; // @[AWSVggWrapper.scala 53:94]
  assign _T_296 = {_T_295,_T_41}; // @[AWSVggWrapper.scala 53:94]
  assign _T_297 = {_T_296,_T_42}; // @[AWSVggWrapper.scala 53:94]
  assign _T_298 = {_T_297,_T_43}; // @[AWSVggWrapper.scala 53:94]
  assign _T_299 = {_T_298,_T_44}; // @[AWSVggWrapper.scala 53:94]
  assign _T_300 = {_T_299,_T_45}; // @[AWSVggWrapper.scala 53:94]
  assign _T_301 = {_T_300,_T_46}; // @[AWSVggWrapper.scala 53:94]
  assign _T_302 = {_T_301,_T_47}; // @[AWSVggWrapper.scala 53:94]
  assign _T_303 = {_T_302,_T_48}; // @[AWSVggWrapper.scala 53:94]
  assign _T_304 = {_T_303,_T_49}; // @[AWSVggWrapper.scala 53:94]
  assign _T_305 = {_T_304,_T_50}; // @[AWSVggWrapper.scala 53:94]
  assign _T_306 = {_T_305,_T_51}; // @[AWSVggWrapper.scala 53:94]
  assign _T_307 = {_T_306,_T_52}; // @[AWSVggWrapper.scala 53:94]
  assign _T_308 = {_T_307,_T_53}; // @[AWSVggWrapper.scala 53:94]
  assign _T_309 = {_T_308,_T_54}; // @[AWSVggWrapper.scala 53:94]
  assign _T_310 = {_T_309,_T_55}; // @[AWSVggWrapper.scala 53:94]
  assign _T_311 = {_T_310,_T_56}; // @[AWSVggWrapper.scala 53:94]
  assign _T_312 = {_T_311,_T_57}; // @[AWSVggWrapper.scala 53:94]
  assign _T_313 = {_T_312,_T_58}; // @[AWSVggWrapper.scala 53:94]
  assign _T_314 = {_T_313,_T_59}; // @[AWSVggWrapper.scala 53:94]
  assign _T_315 = {_T_314,_T_60}; // @[AWSVggWrapper.scala 53:94]
  assign _T_316 = {_T_315,_T_61}; // @[AWSVggWrapper.scala 53:94]
  assign _T_317 = {_T_316,_T_62}; // @[AWSVggWrapper.scala 53:94]
  assign _T_318 = {_T_317,_T_63}; // @[AWSVggWrapper.scala 53:94]
  assign _T_319 = {_T_318,_T_64}; // @[AWSVggWrapper.scala 53:94]
  assign _T_320 = {_T_319,_T_65}; // @[AWSVggWrapper.scala 53:94]
  assign _T_321 = {_T_320,_T_66}; // @[AWSVggWrapper.scala 53:94]
  assign _T_322 = {_T_321,_T_67}; // @[AWSVggWrapper.scala 53:94]
  assign _T_323 = {_T_322,_T_68}; // @[AWSVggWrapper.scala 53:94]
  assign _T_324 = {_T_323,_T_69}; // @[AWSVggWrapper.scala 53:94]
  assign _T_325 = {_T_324,_T_70}; // @[AWSVggWrapper.scala 53:94]
  assign _T_326 = {_T_325,_T_71}; // @[AWSVggWrapper.scala 53:94]
  assign _T_327 = {_T_326,_T_72}; // @[AWSVggWrapper.scala 53:94]
  assign _T_328 = {_T_327,_T_73}; // @[AWSVggWrapper.scala 53:94]
  assign _T_329 = {_T_328,_T_74}; // @[AWSVggWrapper.scala 53:94]
  assign _T_330 = {_T_329,_T_75}; // @[AWSVggWrapper.scala 53:94]
  assign _T_331 = {_T_330,_T_76}; // @[AWSVggWrapper.scala 53:94]
  assign _T_332 = {_T_331,_T_77}; // @[AWSVggWrapper.scala 53:94]
  assign _T_333 = {_T_332,_T_78}; // @[AWSVggWrapper.scala 53:94]
  assign _T_334 = {_T_333,_T_79}; // @[AWSVggWrapper.scala 53:94]
  assign _T_335 = {_T_334,_T_80}; // @[AWSVggWrapper.scala 53:94]
  assign _T_336 = {_T_335,_T_81}; // @[AWSVggWrapper.scala 53:94]
  assign _T_337 = {_T_336,_T_82}; // @[AWSVggWrapper.scala 53:94]
  assign _T_338 = {_T_337,_T_83}; // @[AWSVggWrapper.scala 53:94]
  assign _T_339 = {_T_338,_T_84}; // @[AWSVggWrapper.scala 53:94]
  assign _T_340 = {_T_339,_T_85}; // @[AWSVggWrapper.scala 53:94]
  assign _T_341 = {_T_340,_T_86}; // @[AWSVggWrapper.scala 53:94]
  assign _T_342 = {_T_341,_T_87}; // @[AWSVggWrapper.scala 53:94]
  assign _T_343 = {_T_342,_T_88}; // @[AWSVggWrapper.scala 53:94]
  assign _T_344 = {_T_343,_T_89}; // @[AWSVggWrapper.scala 53:94]
  assign _T_345 = {_T_344,_T_90}; // @[AWSVggWrapper.scala 53:94]
  assign _T_346 = {_T_345,_T_91}; // @[AWSVggWrapper.scala 53:94]
  assign _T_347 = {_T_346,_T_92}; // @[AWSVggWrapper.scala 53:94]
  assign _T_348 = {_T_347,_T_93}; // @[AWSVggWrapper.scala 53:94]
  assign _T_349 = {_T_348,_T_94}; // @[AWSVggWrapper.scala 53:94]
  assign _T_350 = {_T_349,_T_95}; // @[AWSVggWrapper.scala 53:94]
  assign _T_351 = {_T_350,_T_96}; // @[AWSVggWrapper.scala 53:94]
  assign _T_352 = {_T_351,_T_97}; // @[AWSVggWrapper.scala 53:94]
  assign _T_353 = {_T_352,_T_98}; // @[AWSVggWrapper.scala 53:94]
  assign _T_354 = {_T_353,_T_99}; // @[AWSVggWrapper.scala 53:94]
  assign _T_355 = {_T_354,_T_100}; // @[AWSVggWrapper.scala 53:94]
  assign _T_356 = {_T_355,_T_101}; // @[AWSVggWrapper.scala 53:94]
  assign _T_357 = {_T_356,_T_102}; // @[AWSVggWrapper.scala 53:94]
  assign _T_358 = {_T_357,_T_103}; // @[AWSVggWrapper.scala 53:94]
  assign _T_359 = {_T_358,_T_104}; // @[AWSVggWrapper.scala 53:94]
  assign _T_360 = {_T_359,_T_105}; // @[AWSVggWrapper.scala 53:94]
  assign _T_361 = {_T_360,_T_106}; // @[AWSVggWrapper.scala 53:94]
  assign _T_362 = {_T_361,_T_107}; // @[AWSVggWrapper.scala 53:94]
  assign _T_363 = {_T_362,_T_108}; // @[AWSVggWrapper.scala 53:94]
  assign _T_364 = {_T_363,_T_109}; // @[AWSVggWrapper.scala 53:94]
  assign _T_365 = {_T_364,_T_110}; // @[AWSVggWrapper.scala 53:94]
  assign _T_366 = {_T_365,_T_111}; // @[AWSVggWrapper.scala 53:94]
  assign _T_367 = {_T_366,_T_112}; // @[AWSVggWrapper.scala 53:94]
  assign _T_368 = {_T_367,_T_113}; // @[AWSVggWrapper.scala 53:94]
  assign _T_369 = {_T_368,_T_114}; // @[AWSVggWrapper.scala 53:94]
  assign _T_370 = {_T_369,_T_115}; // @[AWSVggWrapper.scala 53:94]
  assign _T_371 = {_T_370,_T_116}; // @[AWSVggWrapper.scala 53:94]
  assign _T_372 = {_T_371,_T_117}; // @[AWSVggWrapper.scala 53:94]
  assign _T_373 = {_T_372,_T_118}; // @[AWSVggWrapper.scala 53:94]
  assign _T_374 = {_T_373,_T_119}; // @[AWSVggWrapper.scala 53:94]
  assign _T_375 = {_T_374,_T_120}; // @[AWSVggWrapper.scala 53:94]
  assign _T_376 = {_T_375,_T_121}; // @[AWSVggWrapper.scala 53:94]
  assign _T_377 = {_T_376,_T_122}; // @[AWSVggWrapper.scala 53:94]
  assign _T_378 = {_T_377,_T_123}; // @[AWSVggWrapper.scala 53:94]
  assign _T_379 = {_T_378,_T_124}; // @[AWSVggWrapper.scala 53:94]
  assign _T_380 = {_T_379,_T_125}; // @[AWSVggWrapper.scala 53:94]
  assign _T_381 = {_T_380,_T_126}; // @[AWSVggWrapper.scala 53:94]
  assign _T_382 = {_T_381,_T_127}; // @[AWSVggWrapper.scala 53:94]
  assign _T_383 = {_T_382,_T_128}; // @[AWSVggWrapper.scala 53:94]
  assign _T_384 = {_T_383,_T_129}; // @[AWSVggWrapper.scala 53:94]
  assign _T_385 = {_T_384,_T_130}; // @[AWSVggWrapper.scala 53:94]
  assign _T_386 = {_T_385,_T_131}; // @[AWSVggWrapper.scala 53:94]
  assign _T_387 = {_T_386,_T_132}; // @[AWSVggWrapper.scala 53:94]
  assign _T_388 = {_T_387,_T_133}; // @[AWSVggWrapper.scala 53:94]
  assign _T_389 = {_T_388,_T_134}; // @[AWSVggWrapper.scala 53:94]
  assign _T_390 = {_T_389,_T_135}; // @[AWSVggWrapper.scala 53:94]
  assign _T_391 = {_T_390,_T_136}; // @[AWSVggWrapper.scala 53:94]
  assign _T_392 = {_T_391,_T_137}; // @[AWSVggWrapper.scala 53:94]
  assign _T_393 = {_T_392,_T_138}; // @[AWSVggWrapper.scala 53:94]
  assign _T_394 = {_T_393,_T_139}; // @[AWSVggWrapper.scala 53:94]
  assign _T_395 = {_T_394,_T_140}; // @[AWSVggWrapper.scala 53:94]
  assign _T_396 = {_T_395,_T_141}; // @[AWSVggWrapper.scala 53:94]
  assign _T_397 = {_T_396,_T_142}; // @[AWSVggWrapper.scala 53:94]
  assign _T_398 = {_T_397,_T_143}; // @[AWSVggWrapper.scala 53:94]
  assign _T_399 = {_T_398,_T_144}; // @[AWSVggWrapper.scala 53:94]
  assign _T_400 = {_T_399,_T_145}; // @[AWSVggWrapper.scala 53:94]
  assign _T_401 = {_T_400,_T_146}; // @[AWSVggWrapper.scala 53:94]
  assign _T_402 = {_T_401,_T_147}; // @[AWSVggWrapper.scala 53:94]
  assign _T_403 = {_T_402,_T_148}; // @[AWSVggWrapper.scala 53:94]
  assign _T_404 = {_T_403,_T_149}; // @[AWSVggWrapper.scala 53:94]
  assign _T_405 = {_T_404,_T_150}; // @[AWSVggWrapper.scala 53:94]
  assign _T_406 = {_T_405,_T_151}; // @[AWSVggWrapper.scala 53:94]
  assign _T_407 = {_T_406,_T_152}; // @[AWSVggWrapper.scala 53:94]
  assign _T_408 = {_T_407,_T_153}; // @[AWSVggWrapper.scala 53:94]
  assign _T_409 = {_T_408,_T_154}; // @[AWSVggWrapper.scala 53:94]
  assign _T_410 = {_T_409,_T_155}; // @[AWSVggWrapper.scala 53:94]
  assign _T_411 = {_T_410,_T_156}; // @[AWSVggWrapper.scala 53:94]
  assign _T_412 = {_T_411,_T_157}; // @[AWSVggWrapper.scala 53:94]
  assign _T_413 = {_T_412,_T_158}; // @[AWSVggWrapper.scala 53:94]
  assign _T_414 = {_T_413,_T_159}; // @[AWSVggWrapper.scala 53:94]
  assign _T_415 = {_T_414,_T_160}; // @[AWSVggWrapper.scala 53:94]
  assign _T_416 = {_T_415,_T_161}; // @[AWSVggWrapper.scala 53:94]
  assign _T_417 = {_T_416,_T_162}; // @[AWSVggWrapper.scala 53:94]
  assign _T_418 = {_T_417,_T_163}; // @[AWSVggWrapper.scala 53:94]
  assign _T_419 = {_T_418,_T_164}; // @[AWSVggWrapper.scala 53:94]
  assign _T_420 = {_T_419,_T_165}; // @[AWSVggWrapper.scala 53:94]
  assign _T_421 = {_T_420,_T_166}; // @[AWSVggWrapper.scala 53:94]
  assign _T_422 = {_T_421,_T_167}; // @[AWSVggWrapper.scala 53:94]
  assign _T_423 = {_T_422,_T_168}; // @[AWSVggWrapper.scala 53:94]
  assign _T_424 = {_T_423,_T_169}; // @[AWSVggWrapper.scala 53:94]
  assign _T_425 = {_T_424,_T_170}; // @[AWSVggWrapper.scala 53:94]
  assign _T_426 = {_T_425,_T_171}; // @[AWSVggWrapper.scala 53:94]
  assign _T_427 = {_T_426,_T_172}; // @[AWSVggWrapper.scala 53:94]
  assign _T_428 = {_T_427,_T_173}; // @[AWSVggWrapper.scala 53:94]
  assign _T_429 = {_T_428,_T_174}; // @[AWSVggWrapper.scala 53:94]
  assign _T_430 = {_T_429,_T_175}; // @[AWSVggWrapper.scala 53:94]
  assign _T_431 = {_T_430,_T_176}; // @[AWSVggWrapper.scala 53:94]
  assign _T_432 = {_T_431,_T_177}; // @[AWSVggWrapper.scala 53:94]
  assign _T_433 = {_T_432,_T_178}; // @[AWSVggWrapper.scala 53:94]
  assign _T_434 = {_T_433,_T_179}; // @[AWSVggWrapper.scala 53:94]
  assign _T_435 = {_T_434,_T_180}; // @[AWSVggWrapper.scala 53:94]
  assign _T_436 = {_T_435,_T_181}; // @[AWSVggWrapper.scala 53:94]
  assign _T_437 = {_T_436,_T_182}; // @[AWSVggWrapper.scala 53:94]
  assign _T_438 = {_T_437,_T_183}; // @[AWSVggWrapper.scala 53:94]
  assign _T_439 = {_T_438,_T_184}; // @[AWSVggWrapper.scala 53:94]
  assign _T_440 = {_T_439,_T_185}; // @[AWSVggWrapper.scala 53:94]
  assign _T_441 = {_T_440,_T_186}; // @[AWSVggWrapper.scala 53:94]
  assign _T_442 = {_T_441,_T_187}; // @[AWSVggWrapper.scala 53:94]
  assign _T_443 = {_T_442,_T_188}; // @[AWSVggWrapper.scala 53:94]
  assign _T_444 = {_T_443,_T_189}; // @[AWSVggWrapper.scala 53:94]
  assign _T_445 = {_T_444,_T_190}; // @[AWSVggWrapper.scala 53:94]
  assign _T_446 = {_T_445,_T_191}; // @[AWSVggWrapper.scala 53:94]
  assign _T_447 = {_T_446,_T_192}; // @[AWSVggWrapper.scala 53:94]
  assign _T_448 = {_T_447,_T_193}; // @[AWSVggWrapper.scala 53:94]
  assign _T_449 = {_T_448,_T_194}; // @[AWSVggWrapper.scala 53:94]
  assign _T_450 = {_T_449,_T_195}; // @[AWSVggWrapper.scala 53:94]
  assign _T_451 = {_T_450,_T_196}; // @[AWSVggWrapper.scala 53:94]
  assign _T_452 = {_T_451,_T_197}; // @[AWSVggWrapper.scala 53:94]
  assign _T_453 = {_T_452,_T_198}; // @[AWSVggWrapper.scala 53:94]
  assign _T_454 = {_T_453,_T_199}; // @[AWSVggWrapper.scala 53:94]
  assign _T_455 = {_T_454,_T_200}; // @[AWSVggWrapper.scala 53:94]
  assign _T_456 = {_T_455,_T_201}; // @[AWSVggWrapper.scala 53:94]
  assign _T_457 = {_T_456,_T_202}; // @[AWSVggWrapper.scala 53:94]
  assign _T_458 = {_T_457,_T_203}; // @[AWSVggWrapper.scala 53:94]
  assign _T_459 = {_T_458,_T_204}; // @[AWSVggWrapper.scala 53:94]
  assign _T_460 = {_T_459,_T_205}; // @[AWSVggWrapper.scala 53:94]
  assign _T_461 = {_T_460,_T_206}; // @[AWSVggWrapper.scala 53:94]
  assign _T_462 = {_T_461,_T_207}; // @[AWSVggWrapper.scala 53:94]
  assign _T_463 = {_T_462,_T_208}; // @[AWSVggWrapper.scala 53:94]
  assign _T_464 = {_T_463,_T_209}; // @[AWSVggWrapper.scala 53:94]
  assign _T_465 = {_T_464,_T_210}; // @[AWSVggWrapper.scala 53:94]
  assign _T_466 = {_T_465,_T_211}; // @[AWSVggWrapper.scala 53:94]
  assign _T_467 = {_T_466,_T_212}; // @[AWSVggWrapper.scala 53:94]
  assign _T_468 = {_T_467,_T_213}; // @[AWSVggWrapper.scala 53:94]
  assign _T_469 = {_T_468,_T_214}; // @[AWSVggWrapper.scala 53:94]
  assign _T_470 = {_T_469,_T_215}; // @[AWSVggWrapper.scala 53:94]
  assign _T_471 = {_T_470,_T_216}; // @[AWSVggWrapper.scala 53:94]
  assign _T_472 = {_T_471,_T_217}; // @[AWSVggWrapper.scala 53:94]
  assign _T_473 = {_T_472,_T_218}; // @[AWSVggWrapper.scala 53:94]
  assign _T_474 = {_T_473,_T_219}; // @[AWSVggWrapper.scala 53:94]
  assign _T_475 = {_T_474,_T_220}; // @[AWSVggWrapper.scala 53:94]
  assign _T_476 = {_T_475,_T_221}; // @[AWSVggWrapper.scala 53:94]
  assign _T_477 = {_T_476,_T_222}; // @[AWSVggWrapper.scala 53:94]
  assign _T_478 = {_T_477,_T_223}; // @[AWSVggWrapper.scala 53:94]
  assign _T_479 = {_T_478,_T_224}; // @[AWSVggWrapper.scala 53:94]
  assign _T_480 = {_T_479,_T_225}; // @[AWSVggWrapper.scala 53:94]
  assign _T_481 = {_T_480,_T_226}; // @[AWSVggWrapper.scala 53:94]
  assign _T_482 = {_T_481,_T_227}; // @[AWSVggWrapper.scala 53:94]
  assign _T_483 = {_T_482,_T_228}; // @[AWSVggWrapper.scala 53:94]
  assign _T_484 = {_T_483,_T_229}; // @[AWSVggWrapper.scala 53:94]
  assign _T_485 = {_T_484,_T_230}; // @[AWSVggWrapper.scala 53:94]
  assign _T_486 = {_T_485,_T_231}; // @[AWSVggWrapper.scala 53:94]
  assign _T_487 = {_T_486,_T_232}; // @[AWSVggWrapper.scala 53:94]
  assign _T_488 = {_T_487,_T_233}; // @[AWSVggWrapper.scala 53:94]
  assign _T_489 = {_T_488,_T_234}; // @[AWSVggWrapper.scala 53:94]
  assign _T_490 = {_T_489,_T_235}; // @[AWSVggWrapper.scala 53:94]
  assign _T_491 = {_T_490,_T_236}; // @[AWSVggWrapper.scala 53:94]
  assign _T_492 = {_T_491,_T_237}; // @[AWSVggWrapper.scala 53:94]
  assign _T_493 = {_T_492,_T_238}; // @[AWSVggWrapper.scala 53:94]
  assign _T_494 = {_T_493,_T_239}; // @[AWSVggWrapper.scala 53:94]
  assign _T_495 = {_T_494,_T_240}; // @[AWSVggWrapper.scala 53:94]
  assign _T_496 = {_T_495,_T_241}; // @[AWSVggWrapper.scala 53:94]
  assign _T_497 = {_T_496,_T_242}; // @[AWSVggWrapper.scala 53:94]
  assign _T_498 = {_T_497,_T_243}; // @[AWSVggWrapper.scala 53:94]
  assign _T_499 = {_T_498,_T_244}; // @[AWSVggWrapper.scala 53:94]
  assign _T_500 = {_T_499,_T_245}; // @[AWSVggWrapper.scala 53:94]
  assign _T_501 = {_T_500,_T_246}; // @[AWSVggWrapper.scala 53:94]
  assign _T_502 = {_T_501,_T_247}; // @[AWSVggWrapper.scala 53:94]
  assign _T_503 = {_T_502,_T_248}; // @[AWSVggWrapper.scala 53:94]
  assign _T_504 = {_T_503,_T_249}; // @[AWSVggWrapper.scala 53:94]
  assign _T_505 = {_T_504,_T_250}; // @[AWSVggWrapper.scala 53:94]
  assign _T_506 = {_T_505,_T_251}; // @[AWSVggWrapper.scala 53:94]
  assign _T_507 = {_T_506,_T_252}; // @[AWSVggWrapper.scala 53:94]
  assign _T_508 = {_T_507,_T_253}; // @[AWSVggWrapper.scala 53:94]
  assign _T_509 = {_T_508,_T_254}; // @[AWSVggWrapper.scala 53:94]
  assign _T_510 = {_T_509,_T_255}; // @[AWSVggWrapper.scala 53:94]
  assign _T_511 = {_T_510,_T_256}; // @[AWSVggWrapper.scala 53:94]
  assign _T_512 = {_T_511,_T_257}; // @[AWSVggWrapper.scala 53:94]
  assign _T_513 = {_T_512,_T_258}; // @[AWSVggWrapper.scala 53:94]
  assign _T_514 = {_T_513,_T_259}; // @[AWSVggWrapper.scala 53:94]
  assign _T_515 = {_T_514,_T_260}; // @[AWSVggWrapper.scala 53:94]
  assign _T_516 = {_T_515,_T_261}; // @[AWSVggWrapper.scala 53:94]
  assign _T_517 = {_T_516,_T_262}; // @[AWSVggWrapper.scala 53:94]
  assign _T_518 = {_T_517,_T_263}; // @[AWSVggWrapper.scala 53:94]
  assign _T_519 = {_T_518,_T_264}; // @[AWSVggWrapper.scala 53:94]
  assign _T_520 = {_T_519,_T_265}; // @[AWSVggWrapper.scala 53:94]
  assign _T_521 = {_T_520,_T_266}; // @[AWSVggWrapper.scala 53:94]
  assign _T_522 = {_T_521,_T_267}; // @[AWSVggWrapper.scala 53:94]
  assign _T_523 = {_T_522,_T_268}; // @[AWSVggWrapper.scala 53:94]
  assign _T_524 = {_T_523,_T_269}; // @[AWSVggWrapper.scala 53:94]
  assign _T_525 = {_T_524,_T_270}; // @[AWSVggWrapper.scala 53:94]
  assign _T_526 = {_T_525,_T_271}; // @[AWSVggWrapper.scala 53:94]
  assign _T_527 = {_T_526,_T_272}; // @[AWSVggWrapper.scala 53:94]
  assign _T_528 = {_T_527,_T_273}; // @[AWSVggWrapper.scala 53:94]
  assign _T_529 = {_T_528,_T_274}; // @[AWSVggWrapper.scala 53:94]
  assign _T_530 = {_T_529,_T_275}; // @[AWSVggWrapper.scala 53:94]
  assign _T_531 = {_T_530,_T_276}; // @[AWSVggWrapper.scala 53:94]
  assign _T_532 = {_T_531,_T_277}; // @[AWSVggWrapper.scala 53:94]
  assign _T_533 = {_T_532,_T_278}; // @[AWSVggWrapper.scala 53:94]
  assign _T_534 = {_T_533,_T_279}; // @[AWSVggWrapper.scala 53:94]
  assign _T_535 = {_T_534,_T_280}; // @[AWSVggWrapper.scala 53:94]
  assign _T_536 = {_T_535,_T_281}; // @[AWSVggWrapper.scala 53:94]
  assign _T_537 = {_T_536,_T_282}; // @[AWSVggWrapper.scala 53:94]
  assign _T_538 = {_T_537,_T_283}; // @[AWSVggWrapper.scala 53:94]
  assign _T_539 = {_T_538,_T_284}; // @[AWSVggWrapper.scala 53:94]
  assign _T_540 = {_T_539,_T_285}; // @[AWSVggWrapper.scala 53:94]
  assign _T_541 = {_T_540,_T_286}; // @[AWSVggWrapper.scala 53:94]
  assign _T_542 = {_T_541,_T_287}; // @[AWSVggWrapper.scala 53:94]
  assign _T_543 = {_T_542,_T_288}; // @[AWSVggWrapper.scala 53:94]
  assign _T_544 = {_T_543,_T_289}; // @[AWSVggWrapper.scala 53:94]
  assign dataInAsUInt = {_T_544,_T_290}; // @[AWSVggWrapper.scala 53:94]
  assign _T_1839 = queueIOOut_io_deq_bits[15:0]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_255 = $signed(_T_1839); // @[AWSVggWrapper.scala 64:110]
  assign _T_1841 = queueIOOut_io_deq_bits[31:16]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_254 = $signed(_T_1841); // @[AWSVggWrapper.scala 64:110]
  assign _T_1843 = queueIOOut_io_deq_bits[47:32]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_253 = $signed(_T_1843); // @[AWSVggWrapper.scala 64:110]
  assign _T_1845 = queueIOOut_io_deq_bits[63:48]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_252 = $signed(_T_1845); // @[AWSVggWrapper.scala 64:110]
  assign _T_1847 = queueIOOut_io_deq_bits[79:64]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_251 = $signed(_T_1847); // @[AWSVggWrapper.scala 64:110]
  assign _T_1849 = queueIOOut_io_deq_bits[95:80]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_250 = $signed(_T_1849); // @[AWSVggWrapper.scala 64:110]
  assign _T_1851 = queueIOOut_io_deq_bits[111:96]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_249 = $signed(_T_1851); // @[AWSVggWrapper.scala 64:110]
  assign _T_1853 = queueIOOut_io_deq_bits[127:112]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_248 = $signed(_T_1853); // @[AWSVggWrapper.scala 64:110]
  assign _T_1855 = queueIOOut_io_deq_bits[143:128]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_247 = $signed(_T_1855); // @[AWSVggWrapper.scala 64:110]
  assign _T_1857 = queueIOOut_io_deq_bits[159:144]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_246 = $signed(_T_1857); // @[AWSVggWrapper.scala 64:110]
  assign _T_1859 = queueIOOut_io_deq_bits[175:160]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_245 = $signed(_T_1859); // @[AWSVggWrapper.scala 64:110]
  assign _T_1861 = queueIOOut_io_deq_bits[191:176]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_244 = $signed(_T_1861); // @[AWSVggWrapper.scala 64:110]
  assign _T_1863 = queueIOOut_io_deq_bits[207:192]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_243 = $signed(_T_1863); // @[AWSVggWrapper.scala 64:110]
  assign _T_1865 = queueIOOut_io_deq_bits[223:208]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_242 = $signed(_T_1865); // @[AWSVggWrapper.scala 64:110]
  assign _T_1867 = queueIOOut_io_deq_bits[239:224]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_241 = $signed(_T_1867); // @[AWSVggWrapper.scala 64:110]
  assign _T_1869 = queueIOOut_io_deq_bits[255:240]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_240 = $signed(_T_1869); // @[AWSVggWrapper.scala 64:110]
  assign _T_1871 = queueIOOut_io_deq_bits[271:256]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_239 = $signed(_T_1871); // @[AWSVggWrapper.scala 64:110]
  assign _T_1873 = queueIOOut_io_deq_bits[287:272]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_238 = $signed(_T_1873); // @[AWSVggWrapper.scala 64:110]
  assign _T_1875 = queueIOOut_io_deq_bits[303:288]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_237 = $signed(_T_1875); // @[AWSVggWrapper.scala 64:110]
  assign _T_1877 = queueIOOut_io_deq_bits[319:304]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_236 = $signed(_T_1877); // @[AWSVggWrapper.scala 64:110]
  assign _T_1879 = queueIOOut_io_deq_bits[335:320]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_235 = $signed(_T_1879); // @[AWSVggWrapper.scala 64:110]
  assign _T_1881 = queueIOOut_io_deq_bits[351:336]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_234 = $signed(_T_1881); // @[AWSVggWrapper.scala 64:110]
  assign _T_1883 = queueIOOut_io_deq_bits[367:352]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_233 = $signed(_T_1883); // @[AWSVggWrapper.scala 64:110]
  assign _T_1885 = queueIOOut_io_deq_bits[383:368]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_232 = $signed(_T_1885); // @[AWSVggWrapper.scala 64:110]
  assign _T_1887 = queueIOOut_io_deq_bits[399:384]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_231 = $signed(_T_1887); // @[AWSVggWrapper.scala 64:110]
  assign _T_1889 = queueIOOut_io_deq_bits[415:400]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_230 = $signed(_T_1889); // @[AWSVggWrapper.scala 64:110]
  assign _T_1891 = queueIOOut_io_deq_bits[431:416]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_229 = $signed(_T_1891); // @[AWSVggWrapper.scala 64:110]
  assign _T_1893 = queueIOOut_io_deq_bits[447:432]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_228 = $signed(_T_1893); // @[AWSVggWrapper.scala 64:110]
  assign _T_1895 = queueIOOut_io_deq_bits[463:448]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_227 = $signed(_T_1895); // @[AWSVggWrapper.scala 64:110]
  assign _T_1897 = queueIOOut_io_deq_bits[479:464]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_226 = $signed(_T_1897); // @[AWSVggWrapper.scala 64:110]
  assign _T_1899 = queueIOOut_io_deq_bits[495:480]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_225 = $signed(_T_1899); // @[AWSVggWrapper.scala 64:110]
  assign _T_1901 = queueIOOut_io_deq_bits[511:496]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_224 = $signed(_T_1901); // @[AWSVggWrapper.scala 64:110]
  assign _T_1903 = queueIOOut_io_deq_bits[527:512]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_223 = $signed(_T_1903); // @[AWSVggWrapper.scala 64:110]
  assign _T_1905 = queueIOOut_io_deq_bits[543:528]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_222 = $signed(_T_1905); // @[AWSVggWrapper.scala 64:110]
  assign _T_1907 = queueIOOut_io_deq_bits[559:544]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_221 = $signed(_T_1907); // @[AWSVggWrapper.scala 64:110]
  assign _T_1909 = queueIOOut_io_deq_bits[575:560]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_220 = $signed(_T_1909); // @[AWSVggWrapper.scala 64:110]
  assign _T_1911 = queueIOOut_io_deq_bits[591:576]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_219 = $signed(_T_1911); // @[AWSVggWrapper.scala 64:110]
  assign _T_1913 = queueIOOut_io_deq_bits[607:592]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_218 = $signed(_T_1913); // @[AWSVggWrapper.scala 64:110]
  assign _T_1915 = queueIOOut_io_deq_bits[623:608]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_217 = $signed(_T_1915); // @[AWSVggWrapper.scala 64:110]
  assign _T_1917 = queueIOOut_io_deq_bits[639:624]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_216 = $signed(_T_1917); // @[AWSVggWrapper.scala 64:110]
  assign _T_1919 = queueIOOut_io_deq_bits[655:640]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_215 = $signed(_T_1919); // @[AWSVggWrapper.scala 64:110]
  assign _T_1921 = queueIOOut_io_deq_bits[671:656]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_214 = $signed(_T_1921); // @[AWSVggWrapper.scala 64:110]
  assign _T_1923 = queueIOOut_io_deq_bits[687:672]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_213 = $signed(_T_1923); // @[AWSVggWrapper.scala 64:110]
  assign _T_1925 = queueIOOut_io_deq_bits[703:688]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_212 = $signed(_T_1925); // @[AWSVggWrapper.scala 64:110]
  assign _T_1927 = queueIOOut_io_deq_bits[719:704]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_211 = $signed(_T_1927); // @[AWSVggWrapper.scala 64:110]
  assign _T_1929 = queueIOOut_io_deq_bits[735:720]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_210 = $signed(_T_1929); // @[AWSVggWrapper.scala 64:110]
  assign _T_1931 = queueIOOut_io_deq_bits[751:736]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_209 = $signed(_T_1931); // @[AWSVggWrapper.scala 64:110]
  assign _T_1933 = queueIOOut_io_deq_bits[767:752]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_208 = $signed(_T_1933); // @[AWSVggWrapper.scala 64:110]
  assign _T_1935 = queueIOOut_io_deq_bits[783:768]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_207 = $signed(_T_1935); // @[AWSVggWrapper.scala 64:110]
  assign _T_1937 = queueIOOut_io_deq_bits[799:784]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_206 = $signed(_T_1937); // @[AWSVggWrapper.scala 64:110]
  assign _T_1939 = queueIOOut_io_deq_bits[815:800]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_205 = $signed(_T_1939); // @[AWSVggWrapper.scala 64:110]
  assign _T_1941 = queueIOOut_io_deq_bits[831:816]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_204 = $signed(_T_1941); // @[AWSVggWrapper.scala 64:110]
  assign _T_1943 = queueIOOut_io_deq_bits[847:832]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_203 = $signed(_T_1943); // @[AWSVggWrapper.scala 64:110]
  assign _T_1945 = queueIOOut_io_deq_bits[863:848]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_202 = $signed(_T_1945); // @[AWSVggWrapper.scala 64:110]
  assign _T_1947 = queueIOOut_io_deq_bits[879:864]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_201 = $signed(_T_1947); // @[AWSVggWrapper.scala 64:110]
  assign _T_1949 = queueIOOut_io_deq_bits[895:880]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_200 = $signed(_T_1949); // @[AWSVggWrapper.scala 64:110]
  assign _T_1951 = queueIOOut_io_deq_bits[911:896]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_199 = $signed(_T_1951); // @[AWSVggWrapper.scala 64:110]
  assign _T_1953 = queueIOOut_io_deq_bits[927:912]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_198 = $signed(_T_1953); // @[AWSVggWrapper.scala 64:110]
  assign _T_1955 = queueIOOut_io_deq_bits[943:928]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_197 = $signed(_T_1955); // @[AWSVggWrapper.scala 64:110]
  assign _T_1957 = queueIOOut_io_deq_bits[959:944]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_196 = $signed(_T_1957); // @[AWSVggWrapper.scala 64:110]
  assign _T_1959 = queueIOOut_io_deq_bits[975:960]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_195 = $signed(_T_1959); // @[AWSVggWrapper.scala 64:110]
  assign _T_1961 = queueIOOut_io_deq_bits[991:976]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_194 = $signed(_T_1961); // @[AWSVggWrapper.scala 64:110]
  assign _T_1963 = queueIOOut_io_deq_bits[1007:992]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_193 = $signed(_T_1963); // @[AWSVggWrapper.scala 64:110]
  assign _T_1965 = queueIOOut_io_deq_bits[1023:1008]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_192 = $signed(_T_1965); // @[AWSVggWrapper.scala 64:110]
  assign _T_1967 = queueIOOut_io_deq_bits[1039:1024]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_191 = $signed(_T_1967); // @[AWSVggWrapper.scala 64:110]
  assign _T_1969 = queueIOOut_io_deq_bits[1055:1040]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_190 = $signed(_T_1969); // @[AWSVggWrapper.scala 64:110]
  assign _T_1971 = queueIOOut_io_deq_bits[1071:1056]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_189 = $signed(_T_1971); // @[AWSVggWrapper.scala 64:110]
  assign _T_1973 = queueIOOut_io_deq_bits[1087:1072]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_188 = $signed(_T_1973); // @[AWSVggWrapper.scala 64:110]
  assign _T_1975 = queueIOOut_io_deq_bits[1103:1088]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_187 = $signed(_T_1975); // @[AWSVggWrapper.scala 64:110]
  assign _T_1977 = queueIOOut_io_deq_bits[1119:1104]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_186 = $signed(_T_1977); // @[AWSVggWrapper.scala 64:110]
  assign _T_1979 = queueIOOut_io_deq_bits[1135:1120]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_185 = $signed(_T_1979); // @[AWSVggWrapper.scala 64:110]
  assign _T_1981 = queueIOOut_io_deq_bits[1151:1136]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_184 = $signed(_T_1981); // @[AWSVggWrapper.scala 64:110]
  assign _T_1983 = queueIOOut_io_deq_bits[1167:1152]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_183 = $signed(_T_1983); // @[AWSVggWrapper.scala 64:110]
  assign _T_1985 = queueIOOut_io_deq_bits[1183:1168]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_182 = $signed(_T_1985); // @[AWSVggWrapper.scala 64:110]
  assign _T_1987 = queueIOOut_io_deq_bits[1199:1184]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_181 = $signed(_T_1987); // @[AWSVggWrapper.scala 64:110]
  assign _T_1989 = queueIOOut_io_deq_bits[1215:1200]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_180 = $signed(_T_1989); // @[AWSVggWrapper.scala 64:110]
  assign _T_1991 = queueIOOut_io_deq_bits[1231:1216]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_179 = $signed(_T_1991); // @[AWSVggWrapper.scala 64:110]
  assign _T_1993 = queueIOOut_io_deq_bits[1247:1232]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_178 = $signed(_T_1993); // @[AWSVggWrapper.scala 64:110]
  assign _T_1995 = queueIOOut_io_deq_bits[1263:1248]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_177 = $signed(_T_1995); // @[AWSVggWrapper.scala 64:110]
  assign _T_1997 = queueIOOut_io_deq_bits[1279:1264]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_176 = $signed(_T_1997); // @[AWSVggWrapper.scala 64:110]
  assign _T_1999 = queueIOOut_io_deq_bits[1295:1280]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_175 = $signed(_T_1999); // @[AWSVggWrapper.scala 64:110]
  assign _T_2001 = queueIOOut_io_deq_bits[1311:1296]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_174 = $signed(_T_2001); // @[AWSVggWrapper.scala 64:110]
  assign _T_2003 = queueIOOut_io_deq_bits[1327:1312]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_173 = $signed(_T_2003); // @[AWSVggWrapper.scala 64:110]
  assign _T_2005 = queueIOOut_io_deq_bits[1343:1328]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_172 = $signed(_T_2005); // @[AWSVggWrapper.scala 64:110]
  assign _T_2007 = queueIOOut_io_deq_bits[1359:1344]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_171 = $signed(_T_2007); // @[AWSVggWrapper.scala 64:110]
  assign _T_2009 = queueIOOut_io_deq_bits[1375:1360]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_170 = $signed(_T_2009); // @[AWSVggWrapper.scala 64:110]
  assign _T_2011 = queueIOOut_io_deq_bits[1391:1376]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_169 = $signed(_T_2011); // @[AWSVggWrapper.scala 64:110]
  assign _T_2013 = queueIOOut_io_deq_bits[1407:1392]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_168 = $signed(_T_2013); // @[AWSVggWrapper.scala 64:110]
  assign _T_2015 = queueIOOut_io_deq_bits[1423:1408]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_167 = $signed(_T_2015); // @[AWSVggWrapper.scala 64:110]
  assign _T_2017 = queueIOOut_io_deq_bits[1439:1424]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_166 = $signed(_T_2017); // @[AWSVggWrapper.scala 64:110]
  assign _T_2019 = queueIOOut_io_deq_bits[1455:1440]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_165 = $signed(_T_2019); // @[AWSVggWrapper.scala 64:110]
  assign _T_2021 = queueIOOut_io_deq_bits[1471:1456]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_164 = $signed(_T_2021); // @[AWSVggWrapper.scala 64:110]
  assign _T_2023 = queueIOOut_io_deq_bits[1487:1472]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_163 = $signed(_T_2023); // @[AWSVggWrapper.scala 64:110]
  assign _T_2025 = queueIOOut_io_deq_bits[1503:1488]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_162 = $signed(_T_2025); // @[AWSVggWrapper.scala 64:110]
  assign _T_2027 = queueIOOut_io_deq_bits[1519:1504]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_161 = $signed(_T_2027); // @[AWSVggWrapper.scala 64:110]
  assign _T_2029 = queueIOOut_io_deq_bits[1535:1520]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_160 = $signed(_T_2029); // @[AWSVggWrapper.scala 64:110]
  assign _T_2031 = queueIOOut_io_deq_bits[1551:1536]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_159 = $signed(_T_2031); // @[AWSVggWrapper.scala 64:110]
  assign _T_2033 = queueIOOut_io_deq_bits[1567:1552]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_158 = $signed(_T_2033); // @[AWSVggWrapper.scala 64:110]
  assign _T_2035 = queueIOOut_io_deq_bits[1583:1568]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_157 = $signed(_T_2035); // @[AWSVggWrapper.scala 64:110]
  assign _T_2037 = queueIOOut_io_deq_bits[1599:1584]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_156 = $signed(_T_2037); // @[AWSVggWrapper.scala 64:110]
  assign _T_2039 = queueIOOut_io_deq_bits[1615:1600]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_155 = $signed(_T_2039); // @[AWSVggWrapper.scala 64:110]
  assign _T_2041 = queueIOOut_io_deq_bits[1631:1616]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_154 = $signed(_T_2041); // @[AWSVggWrapper.scala 64:110]
  assign _T_2043 = queueIOOut_io_deq_bits[1647:1632]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_153 = $signed(_T_2043); // @[AWSVggWrapper.scala 64:110]
  assign _T_2045 = queueIOOut_io_deq_bits[1663:1648]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_152 = $signed(_T_2045); // @[AWSVggWrapper.scala 64:110]
  assign _T_2047 = queueIOOut_io_deq_bits[1679:1664]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_151 = $signed(_T_2047); // @[AWSVggWrapper.scala 64:110]
  assign _T_2049 = queueIOOut_io_deq_bits[1695:1680]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_150 = $signed(_T_2049); // @[AWSVggWrapper.scala 64:110]
  assign _T_2051 = queueIOOut_io_deq_bits[1711:1696]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_149 = $signed(_T_2051); // @[AWSVggWrapper.scala 64:110]
  assign _T_2053 = queueIOOut_io_deq_bits[1727:1712]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_148 = $signed(_T_2053); // @[AWSVggWrapper.scala 64:110]
  assign _T_2055 = queueIOOut_io_deq_bits[1743:1728]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_147 = $signed(_T_2055); // @[AWSVggWrapper.scala 64:110]
  assign _T_2057 = queueIOOut_io_deq_bits[1759:1744]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_146 = $signed(_T_2057); // @[AWSVggWrapper.scala 64:110]
  assign _T_2059 = queueIOOut_io_deq_bits[1775:1760]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_145 = $signed(_T_2059); // @[AWSVggWrapper.scala 64:110]
  assign _T_2061 = queueIOOut_io_deq_bits[1791:1776]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_144 = $signed(_T_2061); // @[AWSVggWrapper.scala 64:110]
  assign _T_2063 = queueIOOut_io_deq_bits[1807:1792]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_143 = $signed(_T_2063); // @[AWSVggWrapper.scala 64:110]
  assign _T_2065 = queueIOOut_io_deq_bits[1823:1808]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_142 = $signed(_T_2065); // @[AWSVggWrapper.scala 64:110]
  assign _T_2067 = queueIOOut_io_deq_bits[1839:1824]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_141 = $signed(_T_2067); // @[AWSVggWrapper.scala 64:110]
  assign _T_2069 = queueIOOut_io_deq_bits[1855:1840]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_140 = $signed(_T_2069); // @[AWSVggWrapper.scala 64:110]
  assign _T_2071 = queueIOOut_io_deq_bits[1871:1856]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_139 = $signed(_T_2071); // @[AWSVggWrapper.scala 64:110]
  assign _T_2073 = queueIOOut_io_deq_bits[1887:1872]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_138 = $signed(_T_2073); // @[AWSVggWrapper.scala 64:110]
  assign _T_2075 = queueIOOut_io_deq_bits[1903:1888]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_137 = $signed(_T_2075); // @[AWSVggWrapper.scala 64:110]
  assign _T_2077 = queueIOOut_io_deq_bits[1919:1904]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_136 = $signed(_T_2077); // @[AWSVggWrapper.scala 64:110]
  assign _T_2079 = queueIOOut_io_deq_bits[1935:1920]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_135 = $signed(_T_2079); // @[AWSVggWrapper.scala 64:110]
  assign _T_2081 = queueIOOut_io_deq_bits[1951:1936]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_134 = $signed(_T_2081); // @[AWSVggWrapper.scala 64:110]
  assign _T_2083 = queueIOOut_io_deq_bits[1967:1952]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_133 = $signed(_T_2083); // @[AWSVggWrapper.scala 64:110]
  assign _T_2085 = queueIOOut_io_deq_bits[1983:1968]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_132 = $signed(_T_2085); // @[AWSVggWrapper.scala 64:110]
  assign _T_2087 = queueIOOut_io_deq_bits[1999:1984]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_131 = $signed(_T_2087); // @[AWSVggWrapper.scala 64:110]
  assign _T_2089 = queueIOOut_io_deq_bits[2015:2000]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_130 = $signed(_T_2089); // @[AWSVggWrapper.scala 64:110]
  assign _T_2091 = queueIOOut_io_deq_bits[2031:2016]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_129 = $signed(_T_2091); // @[AWSVggWrapper.scala 64:110]
  assign _T_2093 = queueIOOut_io_deq_bits[2047:2032]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_128 = $signed(_T_2093); // @[AWSVggWrapper.scala 64:110]
  assign _T_2095 = queueIOOut_io_deq_bits[2063:2048]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_127 = $signed(_T_2095); // @[AWSVggWrapper.scala 64:110]
  assign _T_2097 = queueIOOut_io_deq_bits[2079:2064]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_126 = $signed(_T_2097); // @[AWSVggWrapper.scala 64:110]
  assign _T_2099 = queueIOOut_io_deq_bits[2095:2080]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_125 = $signed(_T_2099); // @[AWSVggWrapper.scala 64:110]
  assign _T_2101 = queueIOOut_io_deq_bits[2111:2096]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_124 = $signed(_T_2101); // @[AWSVggWrapper.scala 64:110]
  assign _T_2103 = queueIOOut_io_deq_bits[2127:2112]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_123 = $signed(_T_2103); // @[AWSVggWrapper.scala 64:110]
  assign _T_2105 = queueIOOut_io_deq_bits[2143:2128]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_122 = $signed(_T_2105); // @[AWSVggWrapper.scala 64:110]
  assign _T_2107 = queueIOOut_io_deq_bits[2159:2144]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_121 = $signed(_T_2107); // @[AWSVggWrapper.scala 64:110]
  assign _T_2109 = queueIOOut_io_deq_bits[2175:2160]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_120 = $signed(_T_2109); // @[AWSVggWrapper.scala 64:110]
  assign _T_2111 = queueIOOut_io_deq_bits[2191:2176]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_119 = $signed(_T_2111); // @[AWSVggWrapper.scala 64:110]
  assign _T_2113 = queueIOOut_io_deq_bits[2207:2192]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_118 = $signed(_T_2113); // @[AWSVggWrapper.scala 64:110]
  assign _T_2115 = queueIOOut_io_deq_bits[2223:2208]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_117 = $signed(_T_2115); // @[AWSVggWrapper.scala 64:110]
  assign _T_2117 = queueIOOut_io_deq_bits[2239:2224]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_116 = $signed(_T_2117); // @[AWSVggWrapper.scala 64:110]
  assign _T_2119 = queueIOOut_io_deq_bits[2255:2240]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_115 = $signed(_T_2119); // @[AWSVggWrapper.scala 64:110]
  assign _T_2121 = queueIOOut_io_deq_bits[2271:2256]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_114 = $signed(_T_2121); // @[AWSVggWrapper.scala 64:110]
  assign _T_2123 = queueIOOut_io_deq_bits[2287:2272]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_113 = $signed(_T_2123); // @[AWSVggWrapper.scala 64:110]
  assign _T_2125 = queueIOOut_io_deq_bits[2303:2288]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_112 = $signed(_T_2125); // @[AWSVggWrapper.scala 64:110]
  assign _T_2127 = queueIOOut_io_deq_bits[2319:2304]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_111 = $signed(_T_2127); // @[AWSVggWrapper.scala 64:110]
  assign _T_2129 = queueIOOut_io_deq_bits[2335:2320]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_110 = $signed(_T_2129); // @[AWSVggWrapper.scala 64:110]
  assign _T_2131 = queueIOOut_io_deq_bits[2351:2336]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_109 = $signed(_T_2131); // @[AWSVggWrapper.scala 64:110]
  assign _T_2133 = queueIOOut_io_deq_bits[2367:2352]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_108 = $signed(_T_2133); // @[AWSVggWrapper.scala 64:110]
  assign _T_2135 = queueIOOut_io_deq_bits[2383:2368]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_107 = $signed(_T_2135); // @[AWSVggWrapper.scala 64:110]
  assign _T_2137 = queueIOOut_io_deq_bits[2399:2384]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_106 = $signed(_T_2137); // @[AWSVggWrapper.scala 64:110]
  assign _T_2139 = queueIOOut_io_deq_bits[2415:2400]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_105 = $signed(_T_2139); // @[AWSVggWrapper.scala 64:110]
  assign _T_2141 = queueIOOut_io_deq_bits[2431:2416]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_104 = $signed(_T_2141); // @[AWSVggWrapper.scala 64:110]
  assign _T_2143 = queueIOOut_io_deq_bits[2447:2432]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_103 = $signed(_T_2143); // @[AWSVggWrapper.scala 64:110]
  assign _T_2145 = queueIOOut_io_deq_bits[2463:2448]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_102 = $signed(_T_2145); // @[AWSVggWrapper.scala 64:110]
  assign _T_2147 = queueIOOut_io_deq_bits[2479:2464]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_101 = $signed(_T_2147); // @[AWSVggWrapper.scala 64:110]
  assign _T_2149 = queueIOOut_io_deq_bits[2495:2480]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_100 = $signed(_T_2149); // @[AWSVggWrapper.scala 64:110]
  assign _T_2151 = queueIOOut_io_deq_bits[2511:2496]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_99 = $signed(_T_2151); // @[AWSVggWrapper.scala 64:110]
  assign _T_2153 = queueIOOut_io_deq_bits[2527:2512]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_98 = $signed(_T_2153); // @[AWSVggWrapper.scala 64:110]
  assign _T_2155 = queueIOOut_io_deq_bits[2543:2528]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_97 = $signed(_T_2155); // @[AWSVggWrapper.scala 64:110]
  assign _T_2157 = queueIOOut_io_deq_bits[2559:2544]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_96 = $signed(_T_2157); // @[AWSVggWrapper.scala 64:110]
  assign _T_2159 = queueIOOut_io_deq_bits[2575:2560]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_95 = $signed(_T_2159); // @[AWSVggWrapper.scala 64:110]
  assign _T_2161 = queueIOOut_io_deq_bits[2591:2576]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_94 = $signed(_T_2161); // @[AWSVggWrapper.scala 64:110]
  assign _T_2163 = queueIOOut_io_deq_bits[2607:2592]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_93 = $signed(_T_2163); // @[AWSVggWrapper.scala 64:110]
  assign _T_2165 = queueIOOut_io_deq_bits[2623:2608]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_92 = $signed(_T_2165); // @[AWSVggWrapper.scala 64:110]
  assign _T_2167 = queueIOOut_io_deq_bits[2639:2624]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_91 = $signed(_T_2167); // @[AWSVggWrapper.scala 64:110]
  assign _T_2169 = queueIOOut_io_deq_bits[2655:2640]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_90 = $signed(_T_2169); // @[AWSVggWrapper.scala 64:110]
  assign _T_2171 = queueIOOut_io_deq_bits[2671:2656]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_89 = $signed(_T_2171); // @[AWSVggWrapper.scala 64:110]
  assign _T_2173 = queueIOOut_io_deq_bits[2687:2672]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_88 = $signed(_T_2173); // @[AWSVggWrapper.scala 64:110]
  assign _T_2175 = queueIOOut_io_deq_bits[2703:2688]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_87 = $signed(_T_2175); // @[AWSVggWrapper.scala 64:110]
  assign _T_2177 = queueIOOut_io_deq_bits[2719:2704]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_86 = $signed(_T_2177); // @[AWSVggWrapper.scala 64:110]
  assign _T_2179 = queueIOOut_io_deq_bits[2735:2720]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_85 = $signed(_T_2179); // @[AWSVggWrapper.scala 64:110]
  assign _T_2181 = queueIOOut_io_deq_bits[2751:2736]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_84 = $signed(_T_2181); // @[AWSVggWrapper.scala 64:110]
  assign _T_2183 = queueIOOut_io_deq_bits[2767:2752]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_83 = $signed(_T_2183); // @[AWSVggWrapper.scala 64:110]
  assign _T_2185 = queueIOOut_io_deq_bits[2783:2768]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_82 = $signed(_T_2185); // @[AWSVggWrapper.scala 64:110]
  assign _T_2187 = queueIOOut_io_deq_bits[2799:2784]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_81 = $signed(_T_2187); // @[AWSVggWrapper.scala 64:110]
  assign _T_2189 = queueIOOut_io_deq_bits[2815:2800]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_80 = $signed(_T_2189); // @[AWSVggWrapper.scala 64:110]
  assign _T_2191 = queueIOOut_io_deq_bits[2831:2816]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_79 = $signed(_T_2191); // @[AWSVggWrapper.scala 64:110]
  assign _T_2193 = queueIOOut_io_deq_bits[2847:2832]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_78 = $signed(_T_2193); // @[AWSVggWrapper.scala 64:110]
  assign _T_2195 = queueIOOut_io_deq_bits[2863:2848]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_77 = $signed(_T_2195); // @[AWSVggWrapper.scala 64:110]
  assign _T_2197 = queueIOOut_io_deq_bits[2879:2864]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_76 = $signed(_T_2197); // @[AWSVggWrapper.scala 64:110]
  assign _T_2199 = queueIOOut_io_deq_bits[2895:2880]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_75 = $signed(_T_2199); // @[AWSVggWrapper.scala 64:110]
  assign _T_2201 = queueIOOut_io_deq_bits[2911:2896]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_74 = $signed(_T_2201); // @[AWSVggWrapper.scala 64:110]
  assign _T_2203 = queueIOOut_io_deq_bits[2927:2912]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_73 = $signed(_T_2203); // @[AWSVggWrapper.scala 64:110]
  assign _T_2205 = queueIOOut_io_deq_bits[2943:2928]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_72 = $signed(_T_2205); // @[AWSVggWrapper.scala 64:110]
  assign _T_2207 = queueIOOut_io_deq_bits[2959:2944]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_71 = $signed(_T_2207); // @[AWSVggWrapper.scala 64:110]
  assign _T_2209 = queueIOOut_io_deq_bits[2975:2960]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_70 = $signed(_T_2209); // @[AWSVggWrapper.scala 64:110]
  assign _T_2211 = queueIOOut_io_deq_bits[2991:2976]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_69 = $signed(_T_2211); // @[AWSVggWrapper.scala 64:110]
  assign _T_2213 = queueIOOut_io_deq_bits[3007:2992]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_68 = $signed(_T_2213); // @[AWSVggWrapper.scala 64:110]
  assign _T_2215 = queueIOOut_io_deq_bits[3023:3008]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_67 = $signed(_T_2215); // @[AWSVggWrapper.scala 64:110]
  assign _T_2217 = queueIOOut_io_deq_bits[3039:3024]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_66 = $signed(_T_2217); // @[AWSVggWrapper.scala 64:110]
  assign _T_2219 = queueIOOut_io_deq_bits[3055:3040]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_65 = $signed(_T_2219); // @[AWSVggWrapper.scala 64:110]
  assign _T_2221 = queueIOOut_io_deq_bits[3071:3056]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_64 = $signed(_T_2221); // @[AWSVggWrapper.scala 64:110]
  assign _T_2223 = queueIOOut_io_deq_bits[3087:3072]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_63 = $signed(_T_2223); // @[AWSVggWrapper.scala 64:110]
  assign _T_2225 = queueIOOut_io_deq_bits[3103:3088]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_62 = $signed(_T_2225); // @[AWSVggWrapper.scala 64:110]
  assign _T_2227 = queueIOOut_io_deq_bits[3119:3104]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_61 = $signed(_T_2227); // @[AWSVggWrapper.scala 64:110]
  assign _T_2229 = queueIOOut_io_deq_bits[3135:3120]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_60 = $signed(_T_2229); // @[AWSVggWrapper.scala 64:110]
  assign _T_2231 = queueIOOut_io_deq_bits[3151:3136]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_59 = $signed(_T_2231); // @[AWSVggWrapper.scala 64:110]
  assign _T_2233 = queueIOOut_io_deq_bits[3167:3152]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_58 = $signed(_T_2233); // @[AWSVggWrapper.scala 64:110]
  assign _T_2235 = queueIOOut_io_deq_bits[3183:3168]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_57 = $signed(_T_2235); // @[AWSVggWrapper.scala 64:110]
  assign _T_2237 = queueIOOut_io_deq_bits[3199:3184]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_56 = $signed(_T_2237); // @[AWSVggWrapper.scala 64:110]
  assign _T_2239 = queueIOOut_io_deq_bits[3215:3200]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_55 = $signed(_T_2239); // @[AWSVggWrapper.scala 64:110]
  assign _T_2241 = queueIOOut_io_deq_bits[3231:3216]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_54 = $signed(_T_2241); // @[AWSVggWrapper.scala 64:110]
  assign _T_2243 = queueIOOut_io_deq_bits[3247:3232]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_53 = $signed(_T_2243); // @[AWSVggWrapper.scala 64:110]
  assign _T_2245 = queueIOOut_io_deq_bits[3263:3248]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_52 = $signed(_T_2245); // @[AWSVggWrapper.scala 64:110]
  assign _T_2247 = queueIOOut_io_deq_bits[3279:3264]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_51 = $signed(_T_2247); // @[AWSVggWrapper.scala 64:110]
  assign _T_2249 = queueIOOut_io_deq_bits[3295:3280]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_50 = $signed(_T_2249); // @[AWSVggWrapper.scala 64:110]
  assign _T_2251 = queueIOOut_io_deq_bits[3311:3296]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_49 = $signed(_T_2251); // @[AWSVggWrapper.scala 64:110]
  assign _T_2253 = queueIOOut_io_deq_bits[3327:3312]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_48 = $signed(_T_2253); // @[AWSVggWrapper.scala 64:110]
  assign _T_2255 = queueIOOut_io_deq_bits[3343:3328]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_47 = $signed(_T_2255); // @[AWSVggWrapper.scala 64:110]
  assign _T_2257 = queueIOOut_io_deq_bits[3359:3344]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_46 = $signed(_T_2257); // @[AWSVggWrapper.scala 64:110]
  assign _T_2259 = queueIOOut_io_deq_bits[3375:3360]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_45 = $signed(_T_2259); // @[AWSVggWrapper.scala 64:110]
  assign _T_2261 = queueIOOut_io_deq_bits[3391:3376]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_44 = $signed(_T_2261); // @[AWSVggWrapper.scala 64:110]
  assign _T_2263 = queueIOOut_io_deq_bits[3407:3392]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_43 = $signed(_T_2263); // @[AWSVggWrapper.scala 64:110]
  assign _T_2265 = queueIOOut_io_deq_bits[3423:3408]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_42 = $signed(_T_2265); // @[AWSVggWrapper.scala 64:110]
  assign _T_2267 = queueIOOut_io_deq_bits[3439:3424]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_41 = $signed(_T_2267); // @[AWSVggWrapper.scala 64:110]
  assign _T_2269 = queueIOOut_io_deq_bits[3455:3440]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_40 = $signed(_T_2269); // @[AWSVggWrapper.scala 64:110]
  assign _T_2271 = queueIOOut_io_deq_bits[3471:3456]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_39 = $signed(_T_2271); // @[AWSVggWrapper.scala 64:110]
  assign _T_2273 = queueIOOut_io_deq_bits[3487:3472]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_38 = $signed(_T_2273); // @[AWSVggWrapper.scala 64:110]
  assign _T_2275 = queueIOOut_io_deq_bits[3503:3488]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_37 = $signed(_T_2275); // @[AWSVggWrapper.scala 64:110]
  assign _T_2277 = queueIOOut_io_deq_bits[3519:3504]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_36 = $signed(_T_2277); // @[AWSVggWrapper.scala 64:110]
  assign _T_2279 = queueIOOut_io_deq_bits[3535:3520]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_35 = $signed(_T_2279); // @[AWSVggWrapper.scala 64:110]
  assign _T_2281 = queueIOOut_io_deq_bits[3551:3536]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_34 = $signed(_T_2281); // @[AWSVggWrapper.scala 64:110]
  assign _T_2283 = queueIOOut_io_deq_bits[3567:3552]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_33 = $signed(_T_2283); // @[AWSVggWrapper.scala 64:110]
  assign _T_2285 = queueIOOut_io_deq_bits[3583:3568]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_32 = $signed(_T_2285); // @[AWSVggWrapper.scala 64:110]
  assign _T_2287 = queueIOOut_io_deq_bits[3599:3584]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_31 = $signed(_T_2287); // @[AWSVggWrapper.scala 64:110]
  assign _T_2289 = queueIOOut_io_deq_bits[3615:3600]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_30 = $signed(_T_2289); // @[AWSVggWrapper.scala 64:110]
  assign _T_2291 = queueIOOut_io_deq_bits[3631:3616]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_29 = $signed(_T_2291); // @[AWSVggWrapper.scala 64:110]
  assign _T_2293 = queueIOOut_io_deq_bits[3647:3632]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_28 = $signed(_T_2293); // @[AWSVggWrapper.scala 64:110]
  assign _T_2295 = queueIOOut_io_deq_bits[3663:3648]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_27 = $signed(_T_2295); // @[AWSVggWrapper.scala 64:110]
  assign _T_2297 = queueIOOut_io_deq_bits[3679:3664]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_26 = $signed(_T_2297); // @[AWSVggWrapper.scala 64:110]
  assign _T_2299 = queueIOOut_io_deq_bits[3695:3680]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_25 = $signed(_T_2299); // @[AWSVggWrapper.scala 64:110]
  assign _T_2301 = queueIOOut_io_deq_bits[3711:3696]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_24 = $signed(_T_2301); // @[AWSVggWrapper.scala 64:110]
  assign _T_2303 = queueIOOut_io_deq_bits[3727:3712]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_23 = $signed(_T_2303); // @[AWSVggWrapper.scala 64:110]
  assign _T_2305 = queueIOOut_io_deq_bits[3743:3728]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_22 = $signed(_T_2305); // @[AWSVggWrapper.scala 64:110]
  assign _T_2307 = queueIOOut_io_deq_bits[3759:3744]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_21 = $signed(_T_2307); // @[AWSVggWrapper.scala 64:110]
  assign _T_2309 = queueIOOut_io_deq_bits[3775:3760]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_20 = $signed(_T_2309); // @[AWSVggWrapper.scala 64:110]
  assign _T_2311 = queueIOOut_io_deq_bits[3791:3776]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_19 = $signed(_T_2311); // @[AWSVggWrapper.scala 64:110]
  assign _T_2313 = queueIOOut_io_deq_bits[3807:3792]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_18 = $signed(_T_2313); // @[AWSVggWrapper.scala 64:110]
  assign _T_2315 = queueIOOut_io_deq_bits[3823:3808]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_17 = $signed(_T_2315); // @[AWSVggWrapper.scala 64:110]
  assign _T_2317 = queueIOOut_io_deq_bits[3839:3824]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_16 = $signed(_T_2317); // @[AWSVggWrapper.scala 64:110]
  assign _T_2319 = queueIOOut_io_deq_bits[3855:3840]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_15 = $signed(_T_2319); // @[AWSVggWrapper.scala 64:110]
  assign _T_2321 = queueIOOut_io_deq_bits[3871:3856]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_14 = $signed(_T_2321); // @[AWSVggWrapper.scala 64:110]
  assign _T_2323 = queueIOOut_io_deq_bits[3887:3872]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_13 = $signed(_T_2323); // @[AWSVggWrapper.scala 64:110]
  assign _T_2325 = queueIOOut_io_deq_bits[3903:3888]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_12 = $signed(_T_2325); // @[AWSVggWrapper.scala 64:110]
  assign _T_2327 = queueIOOut_io_deq_bits[3919:3904]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_11 = $signed(_T_2327); // @[AWSVggWrapper.scala 64:110]
  assign _T_2329 = queueIOOut_io_deq_bits[3935:3920]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_10 = $signed(_T_2329); // @[AWSVggWrapper.scala 64:110]
  assign _T_2331 = queueIOOut_io_deq_bits[3951:3936]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_9 = $signed(_T_2331); // @[AWSVggWrapper.scala 64:110]
  assign _T_2333 = queueIOOut_io_deq_bits[3967:3952]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_8 = $signed(_T_2333); // @[AWSVggWrapper.scala 64:110]
  assign _T_2335 = queueIOOut_io_deq_bits[3983:3968]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_7 = $signed(_T_2335); // @[AWSVggWrapper.scala 64:110]
  assign _T_2337 = queueIOOut_io_deq_bits[3999:3984]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_6 = $signed(_T_2337); // @[AWSVggWrapper.scala 64:110]
  assign _T_2339 = queueIOOut_io_deq_bits[4015:4000]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_5 = $signed(_T_2339); // @[AWSVggWrapper.scala 64:110]
  assign _T_2341 = queueIOOut_io_deq_bits[4031:4016]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_4 = $signed(_T_2341); // @[AWSVggWrapper.scala 64:110]
  assign _T_2343 = queueIOOut_io_deq_bits[4047:4032]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_3 = $signed(_T_2343); // @[AWSVggWrapper.scala 64:110]
  assign _T_2345 = queueIOOut_io_deq_bits[4063:4048]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_2 = $signed(_T_2345); // @[AWSVggWrapper.scala 64:110]
  assign _T_2347 = queueIOOut_io_deq_bits[4079:4064]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_1 = $signed(_T_2347); // @[AWSVggWrapper.scala 64:110]
  assign _T_2349 = queueIOOut_io_deq_bits[4095:4080]; // @[AWSVggWrapper.scala 64:67]
  assign sintOut_0 = $signed(_T_2349); // @[AWSVggWrapper.scala 64:110]
  assign _GEN_0 = dense_2_io_dataOut_valid ? $signed(dense_2_io_dataOut_bits_0) : $signed(outputRegs_0); // @[AWSVggWrapper.scala 109:37]
  assign _GEN_1 = dense_2_io_dataOut_valid ? $signed(dense_2_io_dataOut_bits_1) : $signed(outputRegs_1); // @[AWSVggWrapper.scala 109:37]
  assign _GEN_2 = dense_2_io_dataOut_valid ? $signed(dense_2_io_dataOut_bits_2) : $signed(outputRegs_2); // @[AWSVggWrapper.scala 109:37]
  assign _GEN_3 = dense_2_io_dataOut_valid ? $signed(dense_2_io_dataOut_bits_3) : $signed(outputRegs_3); // @[AWSVggWrapper.scala 109:37]
  assign _GEN_4 = dense_2_io_dataOut_valid ? $signed(dense_2_io_dataOut_bits_4) : $signed(outputRegs_4); // @[AWSVggWrapper.scala 109:37]
  assign _GEN_5 = dense_2_io_dataOut_valid ? $signed(dense_2_io_dataOut_bits_5) : $signed(outputRegs_5); // @[AWSVggWrapper.scala 109:37]
  assign _GEN_6 = dense_2_io_dataOut_valid ? $signed(dense_2_io_dataOut_bits_6) : $signed(outputRegs_6); // @[AWSVggWrapper.scala 109:37]
  assign _GEN_7 = dense_2_io_dataOut_valid ? $signed(dense_2_io_dataOut_bits_7) : $signed(outputRegs_7); // @[AWSVggWrapper.scala 109:37]
  assign _GEN_8 = dense_2_io_dataOut_valid ? $signed(dense_2_io_dataOut_bits_8) : $signed(outputRegs_8); // @[AWSVggWrapper.scala 109:37]
  assign _GEN_9 = dense_2_io_dataOut_valid ? $signed(dense_2_io_dataOut_bits_9) : $signed(outputRegs_9); // @[AWSVggWrapper.scala 109:37]
  assign _GEN_10 = dense_2_io_dataOut_valid; // @[AWSVggWrapper.scala 109:37]
  assign queueIOIn_ready = queueIOOut_io_enq_ready; // @[AWSVggWrapper.scala 54:23]
  assign queueIOIn_valid = vgg_io_dataOut_valid; // @[AWSVggWrapper.scala 54:23]
  assign _T_2353_0 = dense_io_dataOut_bits_0; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_1 = dense_io_dataOut_bits_1; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_2 = dense_io_dataOut_bits_2; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_3 = dense_io_dataOut_bits_3; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_4 = dense_io_dataOut_bits_4; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_5 = dense_io_dataOut_bits_5; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_6 = dense_io_dataOut_bits_6; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_7 = dense_io_dataOut_bits_7; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_8 = dense_io_dataOut_bits_8; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_9 = dense_io_dataOut_bits_9; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_10 = dense_io_dataOut_bits_10; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_11 = dense_io_dataOut_bits_11; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_12 = dense_io_dataOut_bits_12; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_13 = dense_io_dataOut_bits_13; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_14 = dense_io_dataOut_bits_14; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_15 = dense_io_dataOut_bits_15; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_16 = dense_io_dataOut_bits_16; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_17 = dense_io_dataOut_bits_17; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_18 = dense_io_dataOut_bits_18; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_19 = dense_io_dataOut_bits_19; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_20 = dense_io_dataOut_bits_20; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_21 = dense_io_dataOut_bits_21; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_22 = dense_io_dataOut_bits_22; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_23 = dense_io_dataOut_bits_23; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_24 = dense_io_dataOut_bits_24; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_25 = dense_io_dataOut_bits_25; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_26 = dense_io_dataOut_bits_26; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_27 = dense_io_dataOut_bits_27; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_28 = dense_io_dataOut_bits_28; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_29 = dense_io_dataOut_bits_29; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_30 = dense_io_dataOut_bits_30; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_31 = dense_io_dataOut_bits_31; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_32 = dense_io_dataOut_bits_32; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_33 = dense_io_dataOut_bits_33; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_34 = dense_io_dataOut_bits_34; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_35 = dense_io_dataOut_bits_35; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_36 = dense_io_dataOut_bits_36; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_37 = dense_io_dataOut_bits_37; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_38 = dense_io_dataOut_bits_38; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_39 = dense_io_dataOut_bits_39; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_40 = dense_io_dataOut_bits_40; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_41 = dense_io_dataOut_bits_41; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_42 = dense_io_dataOut_bits_42; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_43 = dense_io_dataOut_bits_43; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_44 = dense_io_dataOut_bits_44; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_45 = dense_io_dataOut_bits_45; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_46 = dense_io_dataOut_bits_46; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_47 = dense_io_dataOut_bits_47; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_48 = dense_io_dataOut_bits_48; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_49 = dense_io_dataOut_bits_49; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_50 = dense_io_dataOut_bits_50; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_51 = dense_io_dataOut_bits_51; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_52 = dense_io_dataOut_bits_52; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_53 = dense_io_dataOut_bits_53; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_54 = dense_io_dataOut_bits_54; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_55 = dense_io_dataOut_bits_55; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_56 = dense_io_dataOut_bits_56; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_57 = dense_io_dataOut_bits_57; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_58 = dense_io_dataOut_bits_58; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_59 = dense_io_dataOut_bits_59; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_60 = dense_io_dataOut_bits_60; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_61 = dense_io_dataOut_bits_61; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_62 = dense_io_dataOut_bits_62; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_63 = dense_io_dataOut_bits_63; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_64 = dense_io_dataOut_bits_64; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_65 = dense_io_dataOut_bits_65; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_66 = dense_io_dataOut_bits_66; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_67 = dense_io_dataOut_bits_67; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_68 = dense_io_dataOut_bits_68; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_69 = dense_io_dataOut_bits_69; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_70 = dense_io_dataOut_bits_70; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_71 = dense_io_dataOut_bits_71; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_72 = dense_io_dataOut_bits_72; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_73 = dense_io_dataOut_bits_73; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_74 = dense_io_dataOut_bits_74; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_75 = dense_io_dataOut_bits_75; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_76 = dense_io_dataOut_bits_76; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_77 = dense_io_dataOut_bits_77; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_78 = dense_io_dataOut_bits_78; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_79 = dense_io_dataOut_bits_79; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_80 = dense_io_dataOut_bits_80; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_81 = dense_io_dataOut_bits_81; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_82 = dense_io_dataOut_bits_82; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_83 = dense_io_dataOut_bits_83; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_84 = dense_io_dataOut_bits_84; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_85 = dense_io_dataOut_bits_85; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_86 = dense_io_dataOut_bits_86; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_87 = dense_io_dataOut_bits_87; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_88 = dense_io_dataOut_bits_88; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_89 = dense_io_dataOut_bits_89; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_90 = dense_io_dataOut_bits_90; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_91 = dense_io_dataOut_bits_91; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_92 = dense_io_dataOut_bits_92; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_93 = dense_io_dataOut_bits_93; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_94 = dense_io_dataOut_bits_94; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_95 = dense_io_dataOut_bits_95; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_96 = dense_io_dataOut_bits_96; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_97 = dense_io_dataOut_bits_97; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_98 = dense_io_dataOut_bits_98; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_99 = dense_io_dataOut_bits_99; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_100 = dense_io_dataOut_bits_100; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_101 = dense_io_dataOut_bits_101; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_102 = dense_io_dataOut_bits_102; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_103 = dense_io_dataOut_bits_103; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_104 = dense_io_dataOut_bits_104; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_105 = dense_io_dataOut_bits_105; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_106 = dense_io_dataOut_bits_106; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_107 = dense_io_dataOut_bits_107; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_108 = dense_io_dataOut_bits_108; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_109 = dense_io_dataOut_bits_109; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_110 = dense_io_dataOut_bits_110; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_111 = dense_io_dataOut_bits_111; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_112 = dense_io_dataOut_bits_112; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_113 = dense_io_dataOut_bits_113; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_114 = dense_io_dataOut_bits_114; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_115 = dense_io_dataOut_bits_115; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_116 = dense_io_dataOut_bits_116; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_117 = dense_io_dataOut_bits_117; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_118 = dense_io_dataOut_bits_118; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_119 = dense_io_dataOut_bits_119; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_120 = dense_io_dataOut_bits_120; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_121 = dense_io_dataOut_bits_121; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_122 = dense_io_dataOut_bits_122; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_123 = dense_io_dataOut_bits_123; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_124 = dense_io_dataOut_bits_124; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_125 = dense_io_dataOut_bits_125; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_126 = dense_io_dataOut_bits_126; // @[AWSVggWrapper.scala 83:33]
  assign _T_2353_127 = dense_io_dataOut_bits_127; // @[AWSVggWrapper.scala 83:33]
  assign io_dataIn_ready = vgg_io_dataIn_ready;
  assign io_dataOut_valid = vldReg;
  assign io_dataOut_bits_0 = outputRegs_0;
  assign io_dataOut_bits_1 = outputRegs_1;
  assign io_dataOut_bits_2 = outputRegs_2;
  assign io_dataOut_bits_3 = outputRegs_3;
  assign io_dataOut_bits_4 = outputRegs_4;
  assign io_dataOut_bits_5 = outputRegs_5;
  assign io_dataOut_bits_6 = outputRegs_6;
  assign io_dataOut_bits_7 = outputRegs_7;
  assign io_dataOut_bits_8 = outputRegs_8;
  assign io_dataOut_bits_9 = outputRegs_9;
  assign vgg_clock = clock;
  assign vgg_reset = reset;
  assign vgg_io_dataIn_valid = io_dataIn_valid;
  assign vgg_io_dataIn_bits_0 = io_dataIn_bits_0;
  assign vgg_io_dataIn_bits_1 = io_dataIn_bits_1;
  assign vgg_io_dataIn_bits_2 = io_dataIn_bits_2;
  assign vgg_io_dataOut_ready = queueIOIn_ready;
  assign queueIOOut_clock = clock;
  assign queueIOOut_reset = reset;
  assign queueIOOut_io_enq_valid = queueIOIn_valid;
  assign queueIOOut_io_enq_bits = dataInAsUInt;
  assign queueIOOut_io_deq_ready = muxLyr_io_dataIn_ready;
  assign muxLyr_clock = clock;
  assign muxLyr_reset = reset;
  assign muxLyr_io_dataIn_valid = queueIOOut_io_deq_valid;
  assign muxLyr_io_dataIn_bits_0 = sintOut_0;
  assign muxLyr_io_dataIn_bits_1 = sintOut_1;
  assign muxLyr_io_dataIn_bits_2 = sintOut_2;
  assign muxLyr_io_dataIn_bits_3 = sintOut_3;
  assign muxLyr_io_dataIn_bits_4 = sintOut_4;
  assign muxLyr_io_dataIn_bits_5 = sintOut_5;
  assign muxLyr_io_dataIn_bits_6 = sintOut_6;
  assign muxLyr_io_dataIn_bits_7 = sintOut_7;
  assign muxLyr_io_dataIn_bits_8 = sintOut_8;
  assign muxLyr_io_dataIn_bits_9 = sintOut_9;
  assign muxLyr_io_dataIn_bits_10 = sintOut_10;
  assign muxLyr_io_dataIn_bits_11 = sintOut_11;
  assign muxLyr_io_dataIn_bits_12 = sintOut_12;
  assign muxLyr_io_dataIn_bits_13 = sintOut_13;
  assign muxLyr_io_dataIn_bits_14 = sintOut_14;
  assign muxLyr_io_dataIn_bits_15 = sintOut_15;
  assign muxLyr_io_dataIn_bits_16 = sintOut_16;
  assign muxLyr_io_dataIn_bits_17 = sintOut_17;
  assign muxLyr_io_dataIn_bits_18 = sintOut_18;
  assign muxLyr_io_dataIn_bits_19 = sintOut_19;
  assign muxLyr_io_dataIn_bits_20 = sintOut_20;
  assign muxLyr_io_dataIn_bits_21 = sintOut_21;
  assign muxLyr_io_dataIn_bits_22 = sintOut_22;
  assign muxLyr_io_dataIn_bits_23 = sintOut_23;
  assign muxLyr_io_dataIn_bits_24 = sintOut_24;
  assign muxLyr_io_dataIn_bits_25 = sintOut_25;
  assign muxLyr_io_dataIn_bits_26 = sintOut_26;
  assign muxLyr_io_dataIn_bits_27 = sintOut_27;
  assign muxLyr_io_dataIn_bits_28 = sintOut_28;
  assign muxLyr_io_dataIn_bits_29 = sintOut_29;
  assign muxLyr_io_dataIn_bits_30 = sintOut_30;
  assign muxLyr_io_dataIn_bits_31 = sintOut_31;
  assign muxLyr_io_dataIn_bits_32 = sintOut_32;
  assign muxLyr_io_dataIn_bits_33 = sintOut_33;
  assign muxLyr_io_dataIn_bits_34 = sintOut_34;
  assign muxLyr_io_dataIn_bits_35 = sintOut_35;
  assign muxLyr_io_dataIn_bits_36 = sintOut_36;
  assign muxLyr_io_dataIn_bits_37 = sintOut_37;
  assign muxLyr_io_dataIn_bits_38 = sintOut_38;
  assign muxLyr_io_dataIn_bits_39 = sintOut_39;
  assign muxLyr_io_dataIn_bits_40 = sintOut_40;
  assign muxLyr_io_dataIn_bits_41 = sintOut_41;
  assign muxLyr_io_dataIn_bits_42 = sintOut_42;
  assign muxLyr_io_dataIn_bits_43 = sintOut_43;
  assign muxLyr_io_dataIn_bits_44 = sintOut_44;
  assign muxLyr_io_dataIn_bits_45 = sintOut_45;
  assign muxLyr_io_dataIn_bits_46 = sintOut_46;
  assign muxLyr_io_dataIn_bits_47 = sintOut_47;
  assign muxLyr_io_dataIn_bits_48 = sintOut_48;
  assign muxLyr_io_dataIn_bits_49 = sintOut_49;
  assign muxLyr_io_dataIn_bits_50 = sintOut_50;
  assign muxLyr_io_dataIn_bits_51 = sintOut_51;
  assign muxLyr_io_dataIn_bits_52 = sintOut_52;
  assign muxLyr_io_dataIn_bits_53 = sintOut_53;
  assign muxLyr_io_dataIn_bits_54 = sintOut_54;
  assign muxLyr_io_dataIn_bits_55 = sintOut_55;
  assign muxLyr_io_dataIn_bits_56 = sintOut_56;
  assign muxLyr_io_dataIn_bits_57 = sintOut_57;
  assign muxLyr_io_dataIn_bits_58 = sintOut_58;
  assign muxLyr_io_dataIn_bits_59 = sintOut_59;
  assign muxLyr_io_dataIn_bits_60 = sintOut_60;
  assign muxLyr_io_dataIn_bits_61 = sintOut_61;
  assign muxLyr_io_dataIn_bits_62 = sintOut_62;
  assign muxLyr_io_dataIn_bits_63 = sintOut_63;
  assign muxLyr_io_dataIn_bits_64 = sintOut_64;
  assign muxLyr_io_dataIn_bits_65 = sintOut_65;
  assign muxLyr_io_dataIn_bits_66 = sintOut_66;
  assign muxLyr_io_dataIn_bits_67 = sintOut_67;
  assign muxLyr_io_dataIn_bits_68 = sintOut_68;
  assign muxLyr_io_dataIn_bits_69 = sintOut_69;
  assign muxLyr_io_dataIn_bits_70 = sintOut_70;
  assign muxLyr_io_dataIn_bits_71 = sintOut_71;
  assign muxLyr_io_dataIn_bits_72 = sintOut_72;
  assign muxLyr_io_dataIn_bits_73 = sintOut_73;
  assign muxLyr_io_dataIn_bits_74 = sintOut_74;
  assign muxLyr_io_dataIn_bits_75 = sintOut_75;
  assign muxLyr_io_dataIn_bits_76 = sintOut_76;
  assign muxLyr_io_dataIn_bits_77 = sintOut_77;
  assign muxLyr_io_dataIn_bits_78 = sintOut_78;
  assign muxLyr_io_dataIn_bits_79 = sintOut_79;
  assign muxLyr_io_dataIn_bits_80 = sintOut_80;
  assign muxLyr_io_dataIn_bits_81 = sintOut_81;
  assign muxLyr_io_dataIn_bits_82 = sintOut_82;
  assign muxLyr_io_dataIn_bits_83 = sintOut_83;
  assign muxLyr_io_dataIn_bits_84 = sintOut_84;
  assign muxLyr_io_dataIn_bits_85 = sintOut_85;
  assign muxLyr_io_dataIn_bits_86 = sintOut_86;
  assign muxLyr_io_dataIn_bits_87 = sintOut_87;
  assign muxLyr_io_dataIn_bits_88 = sintOut_88;
  assign muxLyr_io_dataIn_bits_89 = sintOut_89;
  assign muxLyr_io_dataIn_bits_90 = sintOut_90;
  assign muxLyr_io_dataIn_bits_91 = sintOut_91;
  assign muxLyr_io_dataIn_bits_92 = sintOut_92;
  assign muxLyr_io_dataIn_bits_93 = sintOut_93;
  assign muxLyr_io_dataIn_bits_94 = sintOut_94;
  assign muxLyr_io_dataIn_bits_95 = sintOut_95;
  assign muxLyr_io_dataIn_bits_96 = sintOut_96;
  assign muxLyr_io_dataIn_bits_97 = sintOut_97;
  assign muxLyr_io_dataIn_bits_98 = sintOut_98;
  assign muxLyr_io_dataIn_bits_99 = sintOut_99;
  assign muxLyr_io_dataIn_bits_100 = sintOut_100;
  assign muxLyr_io_dataIn_bits_101 = sintOut_101;
  assign muxLyr_io_dataIn_bits_102 = sintOut_102;
  assign muxLyr_io_dataIn_bits_103 = sintOut_103;
  assign muxLyr_io_dataIn_bits_104 = sintOut_104;
  assign muxLyr_io_dataIn_bits_105 = sintOut_105;
  assign muxLyr_io_dataIn_bits_106 = sintOut_106;
  assign muxLyr_io_dataIn_bits_107 = sintOut_107;
  assign muxLyr_io_dataIn_bits_108 = sintOut_108;
  assign muxLyr_io_dataIn_bits_109 = sintOut_109;
  assign muxLyr_io_dataIn_bits_110 = sintOut_110;
  assign muxLyr_io_dataIn_bits_111 = sintOut_111;
  assign muxLyr_io_dataIn_bits_112 = sintOut_112;
  assign muxLyr_io_dataIn_bits_113 = sintOut_113;
  assign muxLyr_io_dataIn_bits_114 = sintOut_114;
  assign muxLyr_io_dataIn_bits_115 = sintOut_115;
  assign muxLyr_io_dataIn_bits_116 = sintOut_116;
  assign muxLyr_io_dataIn_bits_117 = sintOut_117;
  assign muxLyr_io_dataIn_bits_118 = sintOut_118;
  assign muxLyr_io_dataIn_bits_119 = sintOut_119;
  assign muxLyr_io_dataIn_bits_120 = sintOut_120;
  assign muxLyr_io_dataIn_bits_121 = sintOut_121;
  assign muxLyr_io_dataIn_bits_122 = sintOut_122;
  assign muxLyr_io_dataIn_bits_123 = sintOut_123;
  assign muxLyr_io_dataIn_bits_124 = sintOut_124;
  assign muxLyr_io_dataIn_bits_125 = sintOut_125;
  assign muxLyr_io_dataIn_bits_126 = sintOut_126;
  assign muxLyr_io_dataIn_bits_127 = sintOut_127;
  assign muxLyr_io_dataIn_bits_128 = sintOut_128;
  assign muxLyr_io_dataIn_bits_129 = sintOut_129;
  assign muxLyr_io_dataIn_bits_130 = sintOut_130;
  assign muxLyr_io_dataIn_bits_131 = sintOut_131;
  assign muxLyr_io_dataIn_bits_132 = sintOut_132;
  assign muxLyr_io_dataIn_bits_133 = sintOut_133;
  assign muxLyr_io_dataIn_bits_134 = sintOut_134;
  assign muxLyr_io_dataIn_bits_135 = sintOut_135;
  assign muxLyr_io_dataIn_bits_136 = sintOut_136;
  assign muxLyr_io_dataIn_bits_137 = sintOut_137;
  assign muxLyr_io_dataIn_bits_138 = sintOut_138;
  assign muxLyr_io_dataIn_bits_139 = sintOut_139;
  assign muxLyr_io_dataIn_bits_140 = sintOut_140;
  assign muxLyr_io_dataIn_bits_141 = sintOut_141;
  assign muxLyr_io_dataIn_bits_142 = sintOut_142;
  assign muxLyr_io_dataIn_bits_143 = sintOut_143;
  assign muxLyr_io_dataIn_bits_144 = sintOut_144;
  assign muxLyr_io_dataIn_bits_145 = sintOut_145;
  assign muxLyr_io_dataIn_bits_146 = sintOut_146;
  assign muxLyr_io_dataIn_bits_147 = sintOut_147;
  assign muxLyr_io_dataIn_bits_148 = sintOut_148;
  assign muxLyr_io_dataIn_bits_149 = sintOut_149;
  assign muxLyr_io_dataIn_bits_150 = sintOut_150;
  assign muxLyr_io_dataIn_bits_151 = sintOut_151;
  assign muxLyr_io_dataIn_bits_152 = sintOut_152;
  assign muxLyr_io_dataIn_bits_153 = sintOut_153;
  assign muxLyr_io_dataIn_bits_154 = sintOut_154;
  assign muxLyr_io_dataIn_bits_155 = sintOut_155;
  assign muxLyr_io_dataIn_bits_156 = sintOut_156;
  assign muxLyr_io_dataIn_bits_157 = sintOut_157;
  assign muxLyr_io_dataIn_bits_158 = sintOut_158;
  assign muxLyr_io_dataIn_bits_159 = sintOut_159;
  assign muxLyr_io_dataIn_bits_160 = sintOut_160;
  assign muxLyr_io_dataIn_bits_161 = sintOut_161;
  assign muxLyr_io_dataIn_bits_162 = sintOut_162;
  assign muxLyr_io_dataIn_bits_163 = sintOut_163;
  assign muxLyr_io_dataIn_bits_164 = sintOut_164;
  assign muxLyr_io_dataIn_bits_165 = sintOut_165;
  assign muxLyr_io_dataIn_bits_166 = sintOut_166;
  assign muxLyr_io_dataIn_bits_167 = sintOut_167;
  assign muxLyr_io_dataIn_bits_168 = sintOut_168;
  assign muxLyr_io_dataIn_bits_169 = sintOut_169;
  assign muxLyr_io_dataIn_bits_170 = sintOut_170;
  assign muxLyr_io_dataIn_bits_171 = sintOut_171;
  assign muxLyr_io_dataIn_bits_172 = sintOut_172;
  assign muxLyr_io_dataIn_bits_173 = sintOut_173;
  assign muxLyr_io_dataIn_bits_174 = sintOut_174;
  assign muxLyr_io_dataIn_bits_175 = sintOut_175;
  assign muxLyr_io_dataIn_bits_176 = sintOut_176;
  assign muxLyr_io_dataIn_bits_177 = sintOut_177;
  assign muxLyr_io_dataIn_bits_178 = sintOut_178;
  assign muxLyr_io_dataIn_bits_179 = sintOut_179;
  assign muxLyr_io_dataIn_bits_180 = sintOut_180;
  assign muxLyr_io_dataIn_bits_181 = sintOut_181;
  assign muxLyr_io_dataIn_bits_182 = sintOut_182;
  assign muxLyr_io_dataIn_bits_183 = sintOut_183;
  assign muxLyr_io_dataIn_bits_184 = sintOut_184;
  assign muxLyr_io_dataIn_bits_185 = sintOut_185;
  assign muxLyr_io_dataIn_bits_186 = sintOut_186;
  assign muxLyr_io_dataIn_bits_187 = sintOut_187;
  assign muxLyr_io_dataIn_bits_188 = sintOut_188;
  assign muxLyr_io_dataIn_bits_189 = sintOut_189;
  assign muxLyr_io_dataIn_bits_190 = sintOut_190;
  assign muxLyr_io_dataIn_bits_191 = sintOut_191;
  assign muxLyr_io_dataIn_bits_192 = sintOut_192;
  assign muxLyr_io_dataIn_bits_193 = sintOut_193;
  assign muxLyr_io_dataIn_bits_194 = sintOut_194;
  assign muxLyr_io_dataIn_bits_195 = sintOut_195;
  assign muxLyr_io_dataIn_bits_196 = sintOut_196;
  assign muxLyr_io_dataIn_bits_197 = sintOut_197;
  assign muxLyr_io_dataIn_bits_198 = sintOut_198;
  assign muxLyr_io_dataIn_bits_199 = sintOut_199;
  assign muxLyr_io_dataIn_bits_200 = sintOut_200;
  assign muxLyr_io_dataIn_bits_201 = sintOut_201;
  assign muxLyr_io_dataIn_bits_202 = sintOut_202;
  assign muxLyr_io_dataIn_bits_203 = sintOut_203;
  assign muxLyr_io_dataIn_bits_204 = sintOut_204;
  assign muxLyr_io_dataIn_bits_205 = sintOut_205;
  assign muxLyr_io_dataIn_bits_206 = sintOut_206;
  assign muxLyr_io_dataIn_bits_207 = sintOut_207;
  assign muxLyr_io_dataIn_bits_208 = sintOut_208;
  assign muxLyr_io_dataIn_bits_209 = sintOut_209;
  assign muxLyr_io_dataIn_bits_210 = sintOut_210;
  assign muxLyr_io_dataIn_bits_211 = sintOut_211;
  assign muxLyr_io_dataIn_bits_212 = sintOut_212;
  assign muxLyr_io_dataIn_bits_213 = sintOut_213;
  assign muxLyr_io_dataIn_bits_214 = sintOut_214;
  assign muxLyr_io_dataIn_bits_215 = sintOut_215;
  assign muxLyr_io_dataIn_bits_216 = sintOut_216;
  assign muxLyr_io_dataIn_bits_217 = sintOut_217;
  assign muxLyr_io_dataIn_bits_218 = sintOut_218;
  assign muxLyr_io_dataIn_bits_219 = sintOut_219;
  assign muxLyr_io_dataIn_bits_220 = sintOut_220;
  assign muxLyr_io_dataIn_bits_221 = sintOut_221;
  assign muxLyr_io_dataIn_bits_222 = sintOut_222;
  assign muxLyr_io_dataIn_bits_223 = sintOut_223;
  assign muxLyr_io_dataIn_bits_224 = sintOut_224;
  assign muxLyr_io_dataIn_bits_225 = sintOut_225;
  assign muxLyr_io_dataIn_bits_226 = sintOut_226;
  assign muxLyr_io_dataIn_bits_227 = sintOut_227;
  assign muxLyr_io_dataIn_bits_228 = sintOut_228;
  assign muxLyr_io_dataIn_bits_229 = sintOut_229;
  assign muxLyr_io_dataIn_bits_230 = sintOut_230;
  assign muxLyr_io_dataIn_bits_231 = sintOut_231;
  assign muxLyr_io_dataIn_bits_232 = sintOut_232;
  assign muxLyr_io_dataIn_bits_233 = sintOut_233;
  assign muxLyr_io_dataIn_bits_234 = sintOut_234;
  assign muxLyr_io_dataIn_bits_235 = sintOut_235;
  assign muxLyr_io_dataIn_bits_236 = sintOut_236;
  assign muxLyr_io_dataIn_bits_237 = sintOut_237;
  assign muxLyr_io_dataIn_bits_238 = sintOut_238;
  assign muxLyr_io_dataIn_bits_239 = sintOut_239;
  assign muxLyr_io_dataIn_bits_240 = sintOut_240;
  assign muxLyr_io_dataIn_bits_241 = sintOut_241;
  assign muxLyr_io_dataIn_bits_242 = sintOut_242;
  assign muxLyr_io_dataIn_bits_243 = sintOut_243;
  assign muxLyr_io_dataIn_bits_244 = sintOut_244;
  assign muxLyr_io_dataIn_bits_245 = sintOut_245;
  assign muxLyr_io_dataIn_bits_246 = sintOut_246;
  assign muxLyr_io_dataIn_bits_247 = sintOut_247;
  assign muxLyr_io_dataIn_bits_248 = sintOut_248;
  assign muxLyr_io_dataIn_bits_249 = sintOut_249;
  assign muxLyr_io_dataIn_bits_250 = sintOut_250;
  assign muxLyr_io_dataIn_bits_251 = sintOut_251;
  assign muxLyr_io_dataIn_bits_252 = sintOut_252;
  assign muxLyr_io_dataIn_bits_253 = sintOut_253;
  assign muxLyr_io_dataIn_bits_254 = sintOut_254;
  assign muxLyr_io_dataIn_bits_255 = sintOut_255;
  assign dense_clock = clock;
  assign dense_reset = reset;
  assign dense_io_dataIn_valid = muxLyr_io_dataOut_valid;
  assign dense_io_dataIn_bits_0 = muxLyr_io_dataOut_bits_0;
  assign dense_io_dataIn_bits_1 = muxLyr_io_dataOut_bits_1;
  assign dense_io_dataIn_bits_2 = muxLyr_io_dataOut_bits_2;
  assign dense_io_dataIn_bits_3 = muxLyr_io_dataOut_bits_3;
  assign muxLyr_2_clock = clock;
  assign muxLyr_2_reset = reset;
  assign muxLyr_2_io_dataIn_valid = dense_io_dataOut_valid;
  assign muxLyr_2_io_dataIn_bits_0 = _T_2353_0;
  assign muxLyr_2_io_dataIn_bits_1 = _T_2353_1;
  assign muxLyr_2_io_dataIn_bits_2 = _T_2353_2;
  assign muxLyr_2_io_dataIn_bits_3 = _T_2353_3;
  assign muxLyr_2_io_dataIn_bits_4 = _T_2353_4;
  assign muxLyr_2_io_dataIn_bits_5 = _T_2353_5;
  assign muxLyr_2_io_dataIn_bits_6 = _T_2353_6;
  assign muxLyr_2_io_dataIn_bits_7 = _T_2353_7;
  assign muxLyr_2_io_dataIn_bits_8 = _T_2353_8;
  assign muxLyr_2_io_dataIn_bits_9 = _T_2353_9;
  assign muxLyr_2_io_dataIn_bits_10 = _T_2353_10;
  assign muxLyr_2_io_dataIn_bits_11 = _T_2353_11;
  assign muxLyr_2_io_dataIn_bits_12 = _T_2353_12;
  assign muxLyr_2_io_dataIn_bits_13 = _T_2353_13;
  assign muxLyr_2_io_dataIn_bits_14 = _T_2353_14;
  assign muxLyr_2_io_dataIn_bits_15 = _T_2353_15;
  assign muxLyr_2_io_dataIn_bits_16 = _T_2353_16;
  assign muxLyr_2_io_dataIn_bits_17 = _T_2353_17;
  assign muxLyr_2_io_dataIn_bits_18 = _T_2353_18;
  assign muxLyr_2_io_dataIn_bits_19 = _T_2353_19;
  assign muxLyr_2_io_dataIn_bits_20 = _T_2353_20;
  assign muxLyr_2_io_dataIn_bits_21 = _T_2353_21;
  assign muxLyr_2_io_dataIn_bits_22 = _T_2353_22;
  assign muxLyr_2_io_dataIn_bits_23 = _T_2353_23;
  assign muxLyr_2_io_dataIn_bits_24 = _T_2353_24;
  assign muxLyr_2_io_dataIn_bits_25 = _T_2353_25;
  assign muxLyr_2_io_dataIn_bits_26 = _T_2353_26;
  assign muxLyr_2_io_dataIn_bits_27 = _T_2353_27;
  assign muxLyr_2_io_dataIn_bits_28 = _T_2353_28;
  assign muxLyr_2_io_dataIn_bits_29 = _T_2353_29;
  assign muxLyr_2_io_dataIn_bits_30 = _T_2353_30;
  assign muxLyr_2_io_dataIn_bits_31 = _T_2353_31;
  assign muxLyr_2_io_dataIn_bits_32 = _T_2353_32;
  assign muxLyr_2_io_dataIn_bits_33 = _T_2353_33;
  assign muxLyr_2_io_dataIn_bits_34 = _T_2353_34;
  assign muxLyr_2_io_dataIn_bits_35 = _T_2353_35;
  assign muxLyr_2_io_dataIn_bits_36 = _T_2353_36;
  assign muxLyr_2_io_dataIn_bits_37 = _T_2353_37;
  assign muxLyr_2_io_dataIn_bits_38 = _T_2353_38;
  assign muxLyr_2_io_dataIn_bits_39 = _T_2353_39;
  assign muxLyr_2_io_dataIn_bits_40 = _T_2353_40;
  assign muxLyr_2_io_dataIn_bits_41 = _T_2353_41;
  assign muxLyr_2_io_dataIn_bits_42 = _T_2353_42;
  assign muxLyr_2_io_dataIn_bits_43 = _T_2353_43;
  assign muxLyr_2_io_dataIn_bits_44 = _T_2353_44;
  assign muxLyr_2_io_dataIn_bits_45 = _T_2353_45;
  assign muxLyr_2_io_dataIn_bits_46 = _T_2353_46;
  assign muxLyr_2_io_dataIn_bits_47 = _T_2353_47;
  assign muxLyr_2_io_dataIn_bits_48 = _T_2353_48;
  assign muxLyr_2_io_dataIn_bits_49 = _T_2353_49;
  assign muxLyr_2_io_dataIn_bits_50 = _T_2353_50;
  assign muxLyr_2_io_dataIn_bits_51 = _T_2353_51;
  assign muxLyr_2_io_dataIn_bits_52 = _T_2353_52;
  assign muxLyr_2_io_dataIn_bits_53 = _T_2353_53;
  assign muxLyr_2_io_dataIn_bits_54 = _T_2353_54;
  assign muxLyr_2_io_dataIn_bits_55 = _T_2353_55;
  assign muxLyr_2_io_dataIn_bits_56 = _T_2353_56;
  assign muxLyr_2_io_dataIn_bits_57 = _T_2353_57;
  assign muxLyr_2_io_dataIn_bits_58 = _T_2353_58;
  assign muxLyr_2_io_dataIn_bits_59 = _T_2353_59;
  assign muxLyr_2_io_dataIn_bits_60 = _T_2353_60;
  assign muxLyr_2_io_dataIn_bits_61 = _T_2353_61;
  assign muxLyr_2_io_dataIn_bits_62 = _T_2353_62;
  assign muxLyr_2_io_dataIn_bits_63 = _T_2353_63;
  assign muxLyr_2_io_dataIn_bits_64 = _T_2353_64;
  assign muxLyr_2_io_dataIn_bits_65 = _T_2353_65;
  assign muxLyr_2_io_dataIn_bits_66 = _T_2353_66;
  assign muxLyr_2_io_dataIn_bits_67 = _T_2353_67;
  assign muxLyr_2_io_dataIn_bits_68 = _T_2353_68;
  assign muxLyr_2_io_dataIn_bits_69 = _T_2353_69;
  assign muxLyr_2_io_dataIn_bits_70 = _T_2353_70;
  assign muxLyr_2_io_dataIn_bits_71 = _T_2353_71;
  assign muxLyr_2_io_dataIn_bits_72 = _T_2353_72;
  assign muxLyr_2_io_dataIn_bits_73 = _T_2353_73;
  assign muxLyr_2_io_dataIn_bits_74 = _T_2353_74;
  assign muxLyr_2_io_dataIn_bits_75 = _T_2353_75;
  assign muxLyr_2_io_dataIn_bits_76 = _T_2353_76;
  assign muxLyr_2_io_dataIn_bits_77 = _T_2353_77;
  assign muxLyr_2_io_dataIn_bits_78 = _T_2353_78;
  assign muxLyr_2_io_dataIn_bits_79 = _T_2353_79;
  assign muxLyr_2_io_dataIn_bits_80 = _T_2353_80;
  assign muxLyr_2_io_dataIn_bits_81 = _T_2353_81;
  assign muxLyr_2_io_dataIn_bits_82 = _T_2353_82;
  assign muxLyr_2_io_dataIn_bits_83 = _T_2353_83;
  assign muxLyr_2_io_dataIn_bits_84 = _T_2353_84;
  assign muxLyr_2_io_dataIn_bits_85 = _T_2353_85;
  assign muxLyr_2_io_dataIn_bits_86 = _T_2353_86;
  assign muxLyr_2_io_dataIn_bits_87 = _T_2353_87;
  assign muxLyr_2_io_dataIn_bits_88 = _T_2353_88;
  assign muxLyr_2_io_dataIn_bits_89 = _T_2353_89;
  assign muxLyr_2_io_dataIn_bits_90 = _T_2353_90;
  assign muxLyr_2_io_dataIn_bits_91 = _T_2353_91;
  assign muxLyr_2_io_dataIn_bits_92 = _T_2353_92;
  assign muxLyr_2_io_dataIn_bits_93 = _T_2353_93;
  assign muxLyr_2_io_dataIn_bits_94 = _T_2353_94;
  assign muxLyr_2_io_dataIn_bits_95 = _T_2353_95;
  assign muxLyr_2_io_dataIn_bits_96 = _T_2353_96;
  assign muxLyr_2_io_dataIn_bits_97 = _T_2353_97;
  assign muxLyr_2_io_dataIn_bits_98 = _T_2353_98;
  assign muxLyr_2_io_dataIn_bits_99 = _T_2353_99;
  assign muxLyr_2_io_dataIn_bits_100 = _T_2353_100;
  assign muxLyr_2_io_dataIn_bits_101 = _T_2353_101;
  assign muxLyr_2_io_dataIn_bits_102 = _T_2353_102;
  assign muxLyr_2_io_dataIn_bits_103 = _T_2353_103;
  assign muxLyr_2_io_dataIn_bits_104 = _T_2353_104;
  assign muxLyr_2_io_dataIn_bits_105 = _T_2353_105;
  assign muxLyr_2_io_dataIn_bits_106 = _T_2353_106;
  assign muxLyr_2_io_dataIn_bits_107 = _T_2353_107;
  assign muxLyr_2_io_dataIn_bits_108 = _T_2353_108;
  assign muxLyr_2_io_dataIn_bits_109 = _T_2353_109;
  assign muxLyr_2_io_dataIn_bits_110 = _T_2353_110;
  assign muxLyr_2_io_dataIn_bits_111 = _T_2353_111;
  assign muxLyr_2_io_dataIn_bits_112 = _T_2353_112;
  assign muxLyr_2_io_dataIn_bits_113 = _T_2353_113;
  assign muxLyr_2_io_dataIn_bits_114 = _T_2353_114;
  assign muxLyr_2_io_dataIn_bits_115 = _T_2353_115;
  assign muxLyr_2_io_dataIn_bits_116 = _T_2353_116;
  assign muxLyr_2_io_dataIn_bits_117 = _T_2353_117;
  assign muxLyr_2_io_dataIn_bits_118 = _T_2353_118;
  assign muxLyr_2_io_dataIn_bits_119 = _T_2353_119;
  assign muxLyr_2_io_dataIn_bits_120 = _T_2353_120;
  assign muxLyr_2_io_dataIn_bits_121 = _T_2353_121;
  assign muxLyr_2_io_dataIn_bits_122 = _T_2353_122;
  assign muxLyr_2_io_dataIn_bits_123 = _T_2353_123;
  assign muxLyr_2_io_dataIn_bits_124 = _T_2353_124;
  assign muxLyr_2_io_dataIn_bits_125 = _T_2353_125;
  assign muxLyr_2_io_dataIn_bits_126 = _T_2353_126;
  assign muxLyr_2_io_dataIn_bits_127 = _T_2353_127;
  assign scale_clock = clock;
  assign scale_reset = reset;
  assign scale_io_dataIn_valid = muxLyr_2_io_dataOut_valid;
  assign scale_io_dataIn_bits_0 = muxLyr_2_io_dataOut_bits_0;
  assign dense_2_clock = clock;
  assign dense_2_reset = reset;
  assign dense_2_io_dataIn_valid = scale_io_dataOut_valid;
  assign dense_2_io_dataIn_bits_0 = scale_io_dataOut_bits_0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  outputRegs_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  outputRegs_1 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  outputRegs_2 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  outputRegs_3 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  outputRegs_4 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  outputRegs_5 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  outputRegs_6 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  outputRegs_7 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  outputRegs_8 = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  outputRegs_9 = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  vldReg = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (dense_2_io_dataOut_valid) begin
      outputRegs_0 <= dense_2_io_dataOut_bits_0;
    end
    if (dense_2_io_dataOut_valid) begin
      outputRegs_1 <= dense_2_io_dataOut_bits_1;
    end
    if (dense_2_io_dataOut_valid) begin
      outputRegs_2 <= dense_2_io_dataOut_bits_2;
    end
    if (dense_2_io_dataOut_valid) begin
      outputRegs_3 <= dense_2_io_dataOut_bits_3;
    end
    if (dense_2_io_dataOut_valid) begin
      outputRegs_4 <= dense_2_io_dataOut_bits_4;
    end
    if (dense_2_io_dataOut_valid) begin
      outputRegs_5 <= dense_2_io_dataOut_bits_5;
    end
    if (dense_2_io_dataOut_valid) begin
      outputRegs_6 <= dense_2_io_dataOut_bits_6;
    end
    if (dense_2_io_dataOut_valid) begin
      outputRegs_7 <= dense_2_io_dataOut_bits_7;
    end
    if (dense_2_io_dataOut_valid) begin
      outputRegs_8 <= dense_2_io_dataOut_bits_8;
    end
    if (dense_2_io_dataOut_valid) begin
      outputRegs_9 <= dense_2_io_dataOut_bits_9;
    end
    if (reset) begin
      vldReg <= 1'h0;
    end else begin
      vldReg <= _GEN_10;
    end
  end
endmodule
