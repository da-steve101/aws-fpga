
module DenseBlackBox0e5d10d8d8(
  input clock,
  input [9:0] readAddr,
  output [19:0] out
);

reg [19:0] rom_uints [1023:0];
initial
begin
rom_uints[0] = 20'h4c;
rom_uints[1] = 20'h3070;
rom_uints[2] = 20'h40303;
rom_uints[3] = 20'hd00cd;
rom_uints[4] = 20'h4ddf5;
rom_uints[5] = 20'h7f10;
rom_uints[6] = 20'h1743f;
rom_uints[7] = 20'hccc5d;
rom_uints[8] = 20'hf7047;
rom_uints[9] = 20'hcdf51;
rom_uints[10] = 20'h1fcc5;
rom_uints[11] = 20'hcf10;
rom_uints[12] = 20'hdd04c;
rom_uints[13] = 20'h30104;
rom_uints[14] = 20'h7000c;
rom_uints[15] = 20'hff531;
rom_uints[16] = 20'hd0c30;
rom_uints[17] = 20'h5fff5;
rom_uints[18] = 20'h57f;
rom_uints[19] = 20'hc01c7;
rom_uints[20] = 20'h3c700;
rom_uints[21] = 20'h15c3;
rom_uints[22] = 20'hd0773;
rom_uints[23] = 20'h70f3;
rom_uints[24] = 20'h5dd3f;
rom_uints[25] = 20'h5f3f4;
rom_uints[26] = 20'hf7131;
rom_uints[27] = 20'h13d70;
rom_uints[28] = 20'h14c0;
rom_uints[29] = 20'h1f40;
rom_uints[30] = 20'h5f734;
rom_uints[31] = 20'h7f01;
rom_uints[32] = 20'h5373;
rom_uints[33] = 20'hc1037;
rom_uints[34] = 20'h14fc3;
rom_uints[35] = 20'hfc0d5;
rom_uints[36] = 20'h4d31;
rom_uints[37] = 20'hc0577;
rom_uints[38] = 20'h131f3;
rom_uints[39] = 20'h4d300;
rom_uints[40] = 20'hcc7d0;
rom_uints[41] = 20'hc300d;
rom_uints[42] = 20'hdf010;
rom_uints[43] = 20'h3c004;
rom_uints[44] = 20'hc340;
rom_uints[45] = 20'h7fc0;
rom_uints[46] = 20'h4f31;
rom_uints[47] = 20'h13c0;
rom_uints[48] = 20'h73034;
rom_uints[49] = 20'h40030;
rom_uints[50] = 20'h7f04d;
rom_uints[51] = 20'h1dc30;
rom_uints[52] = 20'h3713f;
rom_uints[53] = 20'h3f70;
rom_uints[54] = 20'h73007;
rom_uints[55] = 20'h3d040;
rom_uints[56] = 20'h74fcd;
rom_uints[57] = 20'h11df7;
rom_uints[58] = 20'hd7fd0;
rom_uints[59] = 20'h70dc1;
rom_uints[60] = 20'h17ddc;
rom_uints[61] = 20'hf4730;
rom_uints[62] = 20'h3f440;
rom_uints[63] = 20'h130;
rom_uints[64] = 20'h10cf5;
rom_uints[65] = 20'h5ffc5;
rom_uints[66] = 20'h3f141;
rom_uints[67] = 20'h3c50;
rom_uints[68] = 20'h0;
rom_uints[69] = 20'h4f13;
rom_uints[70] = 20'h5f334;
rom_uints[71] = 20'h3c404;
rom_uints[72] = 20'h3c11;
rom_uints[73] = 20'h4fd1;
rom_uints[74] = 20'hc000;
rom_uints[75] = 20'hcc573;
rom_uints[76] = 20'h7c47c;
rom_uints[77] = 20'h7334c;
rom_uints[78] = 20'h7cd5f;
rom_uints[79] = 20'h3000;
rom_uints[80] = 20'h11ff7;
rom_uints[81] = 20'h7704f;
rom_uints[82] = 20'h1f40;
rom_uints[83] = 20'h44733;
rom_uints[84] = 20'hdf15c;
rom_uints[85] = 20'h401f0;
rom_uints[86] = 20'hcf004;
rom_uints[87] = 20'hc43;
rom_uints[88] = 20'h5f3f5;
rom_uints[89] = 20'hf5c1f;
rom_uints[90] = 20'h31331;
rom_uints[91] = 20'h4fd03;
rom_uints[92] = 20'h500cf;
rom_uints[93] = 20'hfc005;
rom_uints[94] = 20'h7f007;
rom_uints[95] = 20'h135df;
rom_uints[96] = 20'h3c70;
rom_uints[97] = 20'hf040;
rom_uints[98] = 20'h5cf71;
rom_uints[99] = 20'hf475f;
rom_uints[100] = 20'hc03d0;
rom_uints[101] = 20'hc371d;
rom_uints[102] = 20'hcc5d0;
rom_uints[103] = 20'hd5cf;
rom_uints[104] = 20'h3c00;
rom_uints[105] = 20'hf4753;
rom_uints[106] = 20'h73c1c;
rom_uints[107] = 20'hc5c34;
rom_uints[108] = 20'hdc335;
rom_uints[109] = 20'h140fc;
rom_uints[110] = 20'hc17f0;
rom_uints[111] = 20'h47f0;
rom_uints[112] = 20'h4df1c;
rom_uints[113] = 20'h531cc;
rom_uints[114] = 20'hc5f0;
rom_uints[115] = 20'h1341f;
rom_uints[116] = 20'h33753;
rom_uints[117] = 20'hd47;
rom_uints[118] = 20'h5f700;
rom_uints[119] = 20'hd701d;
rom_uints[120] = 20'hc0c04;
rom_uints[121] = 20'h7dd03;
rom_uints[122] = 20'h4;
rom_uints[123] = 20'hc133;
rom_uints[124] = 20'hd0c4d;
rom_uints[125] = 20'h35fdd;
rom_uints[126] = 20'h3c1;
rom_uints[127] = 20'hcfd57;
rom_uints[128] = 20'hc00d0;
rom_uints[129] = 20'hd3503;
rom_uints[130] = 20'h117f3;
rom_uints[131] = 20'hc533;
rom_uints[132] = 20'h4c0;
rom_uints[133] = 20'h4000;
rom_uints[134] = 20'hdd71f;
rom_uints[135] = 20'hfcc53;
rom_uints[136] = 20'h7c1d0;
rom_uints[137] = 20'h3fd50;
rom_uints[138] = 20'hf317;
rom_uints[139] = 20'h1d3;
rom_uints[140] = 20'hf7513;
rom_uints[141] = 20'h773cd;
rom_uints[142] = 20'h44c0;
rom_uints[143] = 20'hf71dd;
rom_uints[144] = 20'hc403;
rom_uints[145] = 20'hd710f;
rom_uints[146] = 20'hcc0;
rom_uints[147] = 20'h1777f;
rom_uints[148] = 20'hf3d0;
rom_uints[149] = 20'h43cc5;
rom_uints[150] = 20'h3f443;
rom_uints[151] = 20'h44fc;
rom_uints[152] = 20'h47f4c;
rom_uints[153] = 20'h30;
rom_uints[154] = 20'h714c3;
rom_uints[155] = 20'hfd01d;
rom_uints[156] = 20'h7cf45;
rom_uints[157] = 20'h30f44;
rom_uints[158] = 20'h71f0;
rom_uints[159] = 20'hcc44c;
rom_uints[160] = 20'h7ccc1;
rom_uints[161] = 20'hd1ccd;
rom_uints[162] = 20'hfcd05;
rom_uints[163] = 20'hf51f;
rom_uints[164] = 20'h40c30;
rom_uints[165] = 20'h131f0;
rom_uints[166] = 20'hf4d35;
rom_uints[167] = 20'h1fd7;
rom_uints[168] = 20'h43773;
rom_uints[169] = 20'h4c00f;
rom_uints[170] = 20'hf77f;
rom_uints[171] = 20'hc0335;
rom_uints[172] = 20'h7347c;
rom_uints[173] = 20'h1cc3;
rom_uints[174] = 20'hc1cd3;
rom_uints[175] = 20'hd430;
rom_uints[176] = 20'h3d3;
rom_uints[177] = 20'h45ff7;
rom_uints[178] = 20'h3c711;
rom_uints[179] = 20'h77dfd;
rom_uints[180] = 20'h37073;
rom_uints[181] = 20'hc7df3;
rom_uints[182] = 20'h4cd;
rom_uints[183] = 20'h1cc7c;
rom_uints[184] = 20'h3dc;
rom_uints[185] = 20'h347d0;
rom_uints[186] = 20'h3c153;
rom_uints[187] = 20'h31fd1;
rom_uints[188] = 20'h40df;
rom_uints[189] = 20'h7c1c1;
rom_uints[190] = 20'h4073d;
rom_uints[191] = 20'h1fd41;
rom_uints[192] = 20'h7c301;
rom_uints[193] = 20'h4c4c1;
rom_uints[194] = 20'hf0cd7;
rom_uints[195] = 20'h3cdc;
rom_uints[196] = 20'h3d5dd;
rom_uints[197] = 20'h43f05;
rom_uints[198] = 20'h375fc;
rom_uints[199] = 20'hc7f14;
rom_uints[200] = 20'h11cf1;
rom_uints[201] = 20'h10373;
rom_uints[202] = 20'h15d7f;
rom_uints[203] = 20'h1ccd0;
rom_uints[204] = 20'h3353f;
rom_uints[205] = 20'h37c1;
rom_uints[206] = 20'h77330;
rom_uints[207] = 20'h1f400;
rom_uints[208] = 20'h7340;
rom_uints[209] = 20'h3cc11;
rom_uints[210] = 20'hf7c0;
rom_uints[211] = 20'h300d1;
rom_uints[212] = 20'h370d0;
rom_uints[213] = 20'h10703;
rom_uints[214] = 20'h37573;
rom_uints[215] = 20'h1cc13;
rom_uints[216] = 20'hf7104;
rom_uints[217] = 20'h13413;
rom_uints[218] = 20'h74cd3;
rom_uints[219] = 20'hf747d;
rom_uints[220] = 20'hc0c13;
rom_uints[221] = 20'hc000c;
rom_uints[222] = 20'h4c47f;
rom_uints[223] = 20'h34f70;
rom_uints[224] = 20'hc0f10;
rom_uints[225] = 20'hf710d;
rom_uints[226] = 20'hf50;
rom_uints[227] = 20'h14f3;
rom_uints[228] = 20'hf4107;
rom_uints[229] = 20'hf40;
rom_uints[230] = 20'h31f53;
rom_uints[231] = 20'hc40;
rom_uints[232] = 20'h74c3;
rom_uints[233] = 20'h5ff34;
rom_uints[234] = 20'h40dcd;
rom_uints[235] = 20'h3dc5f;
rom_uints[236] = 20'h4743;
rom_uints[237] = 20'hd7c0c;
rom_uints[238] = 20'h4fc3;
rom_uints[239] = 20'hd7dc;
rom_uints[240] = 20'hf511f;
rom_uints[241] = 20'h40cc7;
rom_uints[242] = 20'h5f33d;
rom_uints[243] = 20'h1300;
rom_uints[244] = 20'h33c43;
rom_uints[245] = 20'h5cfc4;
rom_uints[246] = 20'h4000;
rom_uints[247] = 20'h33770;
rom_uints[248] = 20'h47d3;
rom_uints[249] = 20'hc710d;
rom_uints[250] = 20'h34dd0;
rom_uints[251] = 20'hcddd;
rom_uints[252] = 20'hcc400;
rom_uints[253] = 20'hc4733;
rom_uints[254] = 20'hd403;
rom_uints[255] = 20'hd31fd;
rom_uints[256] = 20'hc003;
rom_uints[257] = 20'hdc073;
rom_uints[258] = 20'h70c4c;
rom_uints[259] = 20'h143df;
rom_uints[260] = 20'h70037;
rom_uints[261] = 20'h313d3;
rom_uints[262] = 20'h77034;
rom_uints[263] = 20'hcd530;
rom_uints[264] = 20'hc3001;
rom_uints[265] = 20'h100cc;
rom_uints[266] = 20'h315cf;
rom_uints[267] = 20'h1d33;
rom_uints[268] = 20'hc17cd;
rom_uints[269] = 20'h7d5df;
rom_uints[270] = 20'hc1307;
rom_uints[271] = 20'h30177;
rom_uints[272] = 20'hc0f50;
rom_uints[273] = 20'hc7014;
rom_uints[274] = 20'hc3f44;
rom_uints[275] = 20'hf130;
rom_uints[276] = 20'hfd44;
rom_uints[277] = 20'h1c43;
rom_uints[278] = 20'h743cd;
rom_uints[279] = 20'hc301;
rom_uints[280] = 20'hd3ddc;
rom_uints[281] = 20'hc0c34;
rom_uints[282] = 20'h33dd0;
rom_uints[283] = 20'hfd57d;
rom_uints[284] = 20'hf010;
rom_uints[285] = 20'hdd7c;
rom_uints[286] = 20'h0;
rom_uints[287] = 20'h570df;
rom_uints[288] = 20'hf70;
rom_uints[289] = 20'hd4073;
rom_uints[290] = 20'hff51d;
rom_uints[291] = 20'hd034c;
rom_uints[292] = 20'h4f70;
rom_uints[293] = 20'h1303d;
rom_uints[294] = 20'hcf015;
rom_uints[295] = 20'hf44f0;
rom_uints[296] = 20'h347d0;
rom_uints[297] = 20'h1ff4d;
rom_uints[298] = 20'hf155f;
rom_uints[299] = 20'h7cf7;
rom_uints[300] = 20'h7335c;
rom_uints[301] = 20'h7dd3;
rom_uints[302] = 20'h5d5f;
rom_uints[303] = 20'h74;
rom_uints[304] = 20'hc40cd;
rom_uints[305] = 20'h5f037;
rom_uints[306] = 20'h4ffd4;
rom_uints[307] = 20'hc0cc4;
rom_uints[308] = 20'h4343c;
rom_uints[309] = 20'h4030;
rom_uints[310] = 20'hf1c07;
rom_uints[311] = 20'hdd4f0;
rom_uints[312] = 20'hd04c0;
rom_uints[313] = 20'hc530;
rom_uints[314] = 20'h0;
rom_uints[315] = 20'h4503;
rom_uints[316] = 20'hf015f;
rom_uints[317] = 20'hc5743;
rom_uints[318] = 20'h1133;
rom_uints[319] = 20'h4f51c;
rom_uints[320] = 20'h14c0;
rom_uints[321] = 20'h173;
rom_uints[322] = 20'h1f0d0;
rom_uints[323] = 20'hd1c07;
rom_uints[324] = 20'h44fc;
rom_uints[325] = 20'hf5d31;
rom_uints[326] = 20'h1d003;
rom_uints[327] = 20'h33c5d;
rom_uints[328] = 20'hf70;
rom_uints[329] = 20'hd1f04;
rom_uints[330] = 20'h3d05d;
rom_uints[331] = 20'h44f04;
rom_uints[332] = 20'hc5cc1;
rom_uints[333] = 20'hc1133;
rom_uints[334] = 20'hc47c4;
rom_uints[335] = 20'h5ff3;
rom_uints[336] = 20'h73c70;
rom_uints[337] = 20'h30dc;
rom_uints[338] = 20'hd4cf3;
rom_uints[339] = 20'hf75dc;
rom_uints[340] = 20'hc7d53;
rom_uints[341] = 20'hf50d3;
rom_uints[342] = 20'hfd1dd;
rom_uints[343] = 20'hc04c4;
rom_uints[344] = 20'hc043d;
rom_uints[345] = 20'h5f3d5;
rom_uints[346] = 20'h4dfd0;
rom_uints[347] = 20'h35dc0;
rom_uints[348] = 20'hccd10;
rom_uints[349] = 20'hf1c04;
rom_uints[350] = 20'h3f53;
rom_uints[351] = 20'hdfd40;
rom_uints[352] = 20'h3f0d1;
rom_uints[353] = 20'h1fd;
rom_uints[354] = 20'hc1d4f;
rom_uints[355] = 20'h75f73;
rom_uints[356] = 20'h1300;
rom_uints[357] = 20'h503f4;
rom_uints[358] = 20'h14cf0;
rom_uints[359] = 20'hc100;
rom_uints[360] = 20'h41f77;
rom_uints[361] = 20'h307f3;
rom_uints[362] = 20'h113cd;
rom_uints[363] = 20'hd40;
rom_uints[364] = 20'h130f1;
rom_uints[365] = 20'h31f1d;
rom_uints[366] = 20'hfd710;
rom_uints[367] = 20'h3d773;
rom_uints[368] = 20'h503d1;
rom_uints[369] = 20'h7057f;
rom_uints[370] = 20'hc1f1;
rom_uints[371] = 20'hf1731;
rom_uints[372] = 20'hcd741;
rom_uints[373] = 20'hd14cf;
rom_uints[374] = 20'h570cf;
rom_uints[375] = 20'h1cc13;
rom_uints[376] = 20'h7d707;
rom_uints[377] = 20'h370;
rom_uints[378] = 20'h1cf4;
rom_uints[379] = 20'hcc70;
rom_uints[380] = 20'hc131;
rom_uints[381] = 20'h43437;
rom_uints[382] = 20'hf754f;
rom_uints[383] = 20'hd3d0;
rom_uints[384] = 20'h1df3;
rom_uints[385] = 20'h15c3f;
rom_uints[386] = 20'h4cdc3;
rom_uints[387] = 20'hd4337;
rom_uints[388] = 20'hc00c1;
rom_uints[389] = 20'h70f1d;
rom_uints[390] = 20'hf1f0;
rom_uints[391] = 20'h33c41;
rom_uints[392] = 20'hfd503;
rom_uints[393] = 20'h7dc;
rom_uints[394] = 20'h3c71;
rom_uints[395] = 20'h1c5c0;
rom_uints[396] = 20'h4335c;
rom_uints[397] = 20'hcfd51;
rom_uints[398] = 20'h573c4;
rom_uints[399] = 20'hd0f4d;
rom_uints[400] = 20'h7d73c;
rom_uints[401] = 20'hcc053;
rom_uints[402] = 20'h73f0;
rom_uints[403] = 20'h5c3d;
rom_uints[404] = 20'hd7f10;
rom_uints[405] = 20'hd13c;
rom_uints[406] = 20'h13d;
rom_uints[407] = 20'hc43d0;
rom_uints[408] = 20'h1c731;
rom_uints[409] = 20'h5fff4;
rom_uints[410] = 20'h4cfdd;
rom_uints[411] = 20'h5ff77;
rom_uints[412] = 20'h70c0c;
rom_uints[413] = 20'h5c0;
rom_uints[414] = 20'h57f1c;
rom_uints[415] = 20'hcd3c5;
rom_uints[416] = 20'hdf1c4;
rom_uints[417] = 20'h377d7;
rom_uints[418] = 20'h341;
rom_uints[419] = 20'h333d4;
rom_uints[420] = 20'hfc5c4;
rom_uints[421] = 20'h301c1;
rom_uints[422] = 20'hcd4c4;
rom_uints[423] = 20'h3f754;
rom_uints[424] = 20'h40c0c;
rom_uints[425] = 20'h7dc1c;
rom_uints[426] = 20'hc4c10;
rom_uints[427] = 20'hfc50c;
rom_uints[428] = 20'h7c00f;
rom_uints[429] = 20'hf0dc;
rom_uints[430] = 20'hc7035;
rom_uints[431] = 20'hd0044;
rom_uints[432] = 20'h140f0;
rom_uints[433] = 20'hc1c;
rom_uints[434] = 20'h3df41;
rom_uints[435] = 20'hc0134;
rom_uints[436] = 20'h11cdf;
rom_uints[437] = 20'hd1c30;
rom_uints[438] = 20'h7754f;
rom_uints[439] = 20'hc40d0;
rom_uints[440] = 20'hc4c4;
rom_uints[441] = 20'h3341;
rom_uints[442] = 20'h11f43;
rom_uints[443] = 20'hfdf1;
rom_uints[444] = 20'h7103c;
rom_uints[445] = 20'h3c13;
rom_uints[446] = 20'hc7743;
rom_uints[447] = 20'hdc017;
rom_uints[448] = 20'hf5330;
rom_uints[449] = 20'h135f0;
rom_uints[450] = 20'h3000;
rom_uints[451] = 20'hf1777;
rom_uints[452] = 20'h3133d;
rom_uints[453] = 20'h4dcc;
rom_uints[454] = 20'hc4df;
rom_uints[455] = 20'hf04d0;
rom_uints[456] = 20'hf513;
rom_uints[457] = 20'h13053;
rom_uints[458] = 20'hf5dd1;
rom_uints[459] = 20'hcc103;
rom_uints[460] = 20'hd0000;
rom_uints[461] = 20'h3c7c1;
rom_uints[462] = 20'h344d3;
rom_uints[463] = 20'hf454f;
rom_uints[464] = 20'h40f70;
rom_uints[465] = 20'hc4c1;
rom_uints[466] = 20'h30700;
rom_uints[467] = 20'hc5f0;
rom_uints[468] = 20'h13370;
rom_uints[469] = 20'h4d770;
rom_uints[470] = 20'h7413;
rom_uints[471] = 20'h30300;
rom_uints[472] = 20'hdd01d;
rom_uints[473] = 20'h5cc;
rom_uints[474] = 20'h4c7d3;
rom_uints[475] = 20'h1cc70;
rom_uints[476] = 20'h3013;
rom_uints[477] = 20'hf7c11;
rom_uints[478] = 20'h34d1;
rom_uints[479] = 20'hf7040;
rom_uints[480] = 20'hc3c13;
rom_uints[481] = 20'h7d0d7;
rom_uints[482] = 20'hc137;
rom_uints[483] = 20'h7c7d7;
rom_uints[484] = 20'h3d13;
rom_uints[485] = 20'h17d4f;
rom_uints[486] = 20'h5ff11;
rom_uints[487] = 20'hd170;
rom_uints[488] = 20'hc1cdc;
rom_uints[489] = 20'h3f407;
rom_uints[490] = 20'hd70;
rom_uints[491] = 20'h5ccf5;
rom_uints[492] = 20'hc341f;
rom_uints[493] = 20'h343d1;
rom_uints[494] = 20'h5ffc;
rom_uints[495] = 20'hc7734;
rom_uints[496] = 20'h7343;
rom_uints[497] = 20'h75c4c;
rom_uints[498] = 20'h447cf;
rom_uints[499] = 20'hf50d7;
rom_uints[500] = 20'h3c40d;
rom_uints[501] = 20'h3cd47;
rom_uints[502] = 20'hd313;
rom_uints[503] = 20'h3d0c;
rom_uints[504] = 20'hf0314;
rom_uints[505] = 20'h40c3;
rom_uints[506] = 20'h40f77;
rom_uints[507] = 20'h443c3;
rom_uints[508] = 20'h577cf;
rom_uints[509] = 20'hd7f1;
rom_uints[510] = 20'h30c10;
rom_uints[511] = 20'hf51fd;
rom_uints[512] = 20'hc15f7;
rom_uints[513] = 20'h3d7;
rom_uints[514] = 20'h34d3;
rom_uints[515] = 20'hd47fd;
rom_uints[516] = 20'h1c7c0;
rom_uints[517] = 20'h131f;
rom_uints[518] = 20'hc7dd;
rom_uints[519] = 20'h7d3f4;
rom_uints[520] = 20'hdd0c;
rom_uints[521] = 20'hd0dd0;
rom_uints[522] = 20'h71f74;
rom_uints[523] = 20'h77c43;
rom_uints[524] = 20'h4cdd3;
rom_uints[525] = 20'h3371;
rom_uints[526] = 20'hc0f40;
rom_uints[527] = 20'h30c53;
rom_uints[528] = 20'h3dc07;
rom_uints[529] = 20'h3043;
rom_uints[530] = 20'h5ff35;
rom_uints[531] = 20'h17f0;
rom_uints[532] = 20'hd1c70;
rom_uints[533] = 20'hf3374;
rom_uints[534] = 20'h3cc71;
rom_uints[535] = 20'h4fc1;
rom_uints[536] = 20'h7f47;
rom_uints[537] = 20'h33701;
rom_uints[538] = 20'hf7c0;
rom_uints[539] = 20'h7d0;
rom_uints[540] = 20'h4fd7d;
rom_uints[541] = 20'hf04c1;
rom_uints[542] = 20'h4530;
rom_uints[543] = 20'h470d3;
rom_uints[544] = 20'h7d7c;
rom_uints[545] = 20'h407d3;
rom_uints[546] = 20'h437c;
rom_uints[547] = 20'h740f7;
rom_uints[548] = 20'hc1c0;
rom_uints[549] = 20'h303c1;
rom_uints[550] = 20'h34f71;
rom_uints[551] = 20'h100c0;
rom_uints[552] = 20'hcdddd;
rom_uints[553] = 20'hcd77;
rom_uints[554] = 20'h4f7c0;
rom_uints[555] = 20'h14c13;
rom_uints[556] = 20'hd3f01;
rom_uints[557] = 20'h30c01;
rom_uints[558] = 20'h17c3;
rom_uints[559] = 20'hdc5c3;
rom_uints[560] = 20'hf740d;
rom_uints[561] = 20'h4cc07;
rom_uints[562] = 20'h30004;
rom_uints[563] = 20'hfdc15;
rom_uints[564] = 20'hc40;
rom_uints[565] = 20'h70dc4;
rom_uints[566] = 20'h3d4f3;
rom_uints[567] = 20'h7007c;
rom_uints[568] = 20'hd0c44;
rom_uints[569] = 20'h4c00c;
rom_uints[570] = 20'hd0df1;
rom_uints[571] = 20'h3f73;
rom_uints[572] = 20'hf41;
rom_uints[573] = 20'h1c073;
rom_uints[574] = 20'hf170;
rom_uints[575] = 20'h7ccc5;
rom_uints[576] = 20'h7f537;
rom_uints[577] = 20'hd4f73;
rom_uints[578] = 20'h43730;
rom_uints[579] = 20'hd340;
rom_uints[580] = 20'h37070;
rom_uints[581] = 20'hddf1c;
rom_uints[582] = 20'hf433;
rom_uints[583] = 20'hc71dc;
rom_uints[584] = 20'hd043f;
rom_uints[585] = 20'hcd0d3;
rom_uints[586] = 20'hdc707;
rom_uints[587] = 20'h77cf5;
rom_uints[588] = 20'hf7750;
rom_uints[589] = 20'h330d0;
rom_uints[590] = 20'h313;
rom_uints[591] = 20'hf4434;
rom_uints[592] = 20'hf307d;
rom_uints[593] = 20'hf4743;
rom_uints[594] = 20'h774fd;
rom_uints[595] = 20'h4733;
rom_uints[596] = 20'hf00d1;
rom_uints[597] = 20'hc4d30;
rom_uints[598] = 20'h1cddc;
rom_uints[599] = 20'h1c130;
rom_uints[600] = 20'h7dfc;
rom_uints[601] = 20'hfc010;
rom_uints[602] = 20'hc11f1;
rom_uints[603] = 20'h71fc4;
rom_uints[604] = 20'h350c3;
rom_uints[605] = 20'h33fd1;
rom_uints[606] = 20'hfd1dd;
rom_uints[607] = 20'h7f74c;
rom_uints[608] = 20'h17003;
rom_uints[609] = 20'h54fcd;
rom_uints[610] = 20'hcd0d0;
rom_uints[611] = 20'h335c0;
rom_uints[612] = 20'h1d343;
rom_uints[613] = 20'hc70;
rom_uints[614] = 20'h5cf0;
rom_uints[615] = 20'h774d0;
rom_uints[616] = 20'h13c0;
rom_uints[617] = 20'h1c4c3;
rom_uints[618] = 20'h300;
rom_uints[619] = 20'hd310;
rom_uints[620] = 20'hc71;
rom_uints[621] = 20'hd17c3;
rom_uints[622] = 20'hc0000;
rom_uints[623] = 20'h54f7d;
rom_uints[624] = 20'h477d3;
rom_uints[625] = 20'hc1f47;
rom_uints[626] = 20'h44c0;
rom_uints[627] = 20'h3d71f;
rom_uints[628] = 20'h30430;
rom_uints[629] = 20'h10c30;
rom_uints[630] = 20'hf0434;
rom_uints[631] = 20'hcd177;
rom_uints[632] = 20'hcc0d0;
rom_uints[633] = 20'hfc10;
rom_uints[634] = 20'h730d3;
rom_uints[635] = 20'hd53dc;
rom_uints[636] = 20'h5fdc1;
rom_uints[637] = 20'hfdd05;
rom_uints[638] = 20'h33c75;
rom_uints[639] = 20'h3f11d;
rom_uints[640] = 20'h5033;
rom_uints[641] = 20'hf74d1;
rom_uints[642] = 20'hd0f00;
rom_uints[643] = 20'hd0c44;
rom_uints[644] = 20'hf40f4;
rom_uints[645] = 20'h4d3f7;
rom_uints[646] = 20'h375f3;
rom_uints[647] = 20'hf0d0;
rom_uints[648] = 20'hf4c;
rom_uints[649] = 20'hc44f7;
rom_uints[650] = 20'hdf050;
rom_uints[651] = 20'h11333;
rom_uints[652] = 20'h74fc;
rom_uints[653] = 20'h3c53;
rom_uints[654] = 20'h3340;
rom_uints[655] = 20'h7300;
rom_uints[656] = 20'h3fc14;
rom_uints[657] = 20'hc7d0;
rom_uints[658] = 20'h1730;
rom_uints[659] = 20'h4df0;
rom_uints[660] = 20'h3d5d3;
rom_uints[661] = 20'h47dcc;
rom_uints[662] = 20'hf5fc4;
rom_uints[663] = 20'h30353;
rom_uints[664] = 20'hdc343;
rom_uints[665] = 20'hfcc45;
rom_uints[666] = 20'h51d3f;
rom_uints[667] = 20'h4c7dc;
rom_uints[668] = 20'hc4df5;
rom_uints[669] = 20'hd05c0;
rom_uints[670] = 20'hc5030;
rom_uints[671] = 20'h1c003;
rom_uints[672] = 20'h77c1f;
rom_uints[673] = 20'h33d04;
rom_uints[674] = 20'h3fd11;
rom_uints[675] = 20'h3cd3;
rom_uints[676] = 20'h5d7f7;
rom_uints[677] = 20'h457fc;
rom_uints[678] = 20'hf7531;
rom_uints[679] = 20'hccf15;
rom_uints[680] = 20'hc7cd7;
rom_uints[681] = 20'h53f3;
rom_uints[682] = 20'h45f13;
rom_uints[683] = 20'hf3dd5;
rom_uints[684] = 20'h3c13;
rom_uints[685] = 20'h1c70;
rom_uints[686] = 20'hcdd31;
rom_uints[687] = 20'h3c44;
rom_uints[688] = 20'h1ff41;
rom_uints[689] = 20'hd1f;
rom_uints[690] = 20'hdc430;
rom_uints[691] = 20'hf573;
rom_uints[692] = 20'h14f43;
rom_uints[693] = 20'h3c1f1;
rom_uints[694] = 20'h4330;
rom_uints[695] = 20'hccc53;
rom_uints[696] = 20'hcc110;
rom_uints[697] = 20'h4f4fc;
rom_uints[698] = 20'hc7573;
rom_uints[699] = 20'hc341;
rom_uints[700] = 20'h71f7;
rom_uints[701] = 20'h34c0;
rom_uints[702] = 20'hfc470;
rom_uints[703] = 20'h353d3;
rom_uints[704] = 20'h4071c;
rom_uints[705] = 20'h3d13;
rom_uints[706] = 20'h17c3;
rom_uints[707] = 20'hc1d3;
rom_uints[708] = 20'h4ff4;
rom_uints[709] = 20'hff411;
rom_uints[710] = 20'h73;
rom_uints[711] = 20'h70340;
rom_uints[712] = 20'hc000;
rom_uints[713] = 20'hc40;
rom_uints[714] = 20'h3c4d;
rom_uints[715] = 20'h3c51f;
rom_uints[716] = 20'hc5f34;
rom_uints[717] = 20'h45f3;
rom_uints[718] = 20'hc0cd1;
rom_uints[719] = 20'hdc1d0;
rom_uints[720] = 20'hfd710;
rom_uints[721] = 20'hfdd03;
rom_uints[722] = 20'hc1;
rom_uints[723] = 20'hc04f1;
rom_uints[724] = 20'hf01c7;
rom_uints[725] = 20'h71f40;
rom_uints[726] = 20'hc7d0;
rom_uints[727] = 20'h30d3;
rom_uints[728] = 20'h33471;
rom_uints[729] = 20'hc04c0;
rom_uints[730] = 20'hdd1f1;
rom_uints[731] = 20'hd7cd1;
rom_uints[732] = 20'h0;
rom_uints[733] = 20'h47d31;
rom_uints[734] = 20'hc3753;
rom_uints[735] = 20'h130f;
rom_uints[736] = 20'hc3c71;
rom_uints[737] = 20'h33d40;
rom_uints[738] = 20'hc47f7;
rom_uints[739] = 20'hcf470;
rom_uints[740] = 20'hdfd01;
rom_uints[741] = 20'h403;
rom_uints[742] = 20'h10c5f;
rom_uints[743] = 20'h744f1;
rom_uints[744] = 20'h504f0;
rom_uints[745] = 20'hc5c7;
rom_uints[746] = 20'hcf3d4;
rom_uints[747] = 20'h13f10;
rom_uints[748] = 20'hcd77;
rom_uints[749] = 20'h3f51;
rom_uints[750] = 20'hffc45;
rom_uints[751] = 20'hc4f40;
rom_uints[752] = 20'h31d3;
rom_uints[753] = 20'hc3c0d;
rom_uints[754] = 20'hfd70;
rom_uints[755] = 20'h3745f;
rom_uints[756] = 20'h40cd7;
rom_uints[757] = 20'hf7703;
rom_uints[758] = 20'hf440;
rom_uints[759] = 20'h4f53;
rom_uints[760] = 20'hf1375;
rom_uints[761] = 20'h3ddc;
rom_uints[762] = 20'h5c34c;
rom_uints[763] = 20'hd703;
rom_uints[764] = 20'h400fd;
rom_uints[765] = 20'hf1430;
rom_uints[766] = 20'h707c0;
rom_uints[767] = 20'hcd530;
rom_uints[768] = 20'h71c0f;
rom_uints[769] = 20'h0;
rom_uints[770] = 20'h430;
rom_uints[771] = 20'hd0c31;
rom_uints[772] = 20'hccd;
rom_uints[773] = 20'h1f100;
rom_uints[774] = 20'hd70;
rom_uints[775] = 20'h1300c;
rom_uints[776] = 20'h1c40;
rom_uints[777] = 20'h3;
rom_uints[778] = 20'hf4717;
rom_uints[779] = 20'h13fd;
rom_uints[780] = 20'hcd55f;
rom_uints[781] = 20'hd3d1d;
rom_uints[782] = 20'h104f0;
rom_uints[783] = 20'hd0730;
rom_uints[784] = 20'h5317c;
rom_uints[785] = 20'h13f44;
rom_uints[786] = 20'h3c5d3;
rom_uints[787] = 20'h30345;
rom_uints[788] = 20'hfd77d;
rom_uints[789] = 20'h40;
rom_uints[790] = 20'hcf114;
rom_uints[791] = 20'h130;
rom_uints[792] = 20'h1c00;
rom_uints[793] = 20'h74f00;
rom_uints[794] = 20'h10f5f;
rom_uints[795] = 20'h7007f;
rom_uints[796] = 20'h1371;
rom_uints[797] = 20'h30003;
rom_uints[798] = 20'h771cf;
rom_uints[799] = 20'h407f4;
rom_uints[800] = 20'h7cd0c;
rom_uints[801] = 20'hcd000;
rom_uints[802] = 20'h3f771;
rom_uints[803] = 20'hc7537;
rom_uints[804] = 20'hcc7c4;
rom_uints[805] = 20'h73403;
rom_uints[806] = 20'hc37d1;
rom_uints[807] = 20'hd04c0;
rom_uints[808] = 20'hcd3d0;
rom_uints[809] = 20'hd077;
rom_uints[810] = 20'hf57cc;
rom_uints[811] = 20'hc10f0;
rom_uints[812] = 20'h4f1fc;
rom_uints[813] = 20'h53cf;
rom_uints[814] = 20'h74c7;
rom_uints[815] = 20'h3c1cd;
rom_uints[816] = 20'hfd45f;
rom_uints[817] = 20'hf1d50;
rom_uints[818] = 20'hf7c0;
rom_uints[819] = 20'h1c3c5;
rom_uints[820] = 20'hcc1f4;
rom_uints[821] = 20'h10c30;
rom_uints[822] = 20'hcd17;
rom_uints[823] = 20'h3df0;
rom_uints[824] = 20'h4f433;
rom_uints[825] = 20'h74df3;
rom_uints[826] = 20'h31;
rom_uints[827] = 20'h34103;
rom_uints[828] = 20'hf5d03;
rom_uints[829] = 20'h310c0;
rom_uints[830] = 20'hf71c4;
rom_uints[831] = 20'hcf4c4;
rom_uints[832] = 20'h1130;
rom_uints[833] = 20'hc4c40;
rom_uints[834] = 20'hdd003;
rom_uints[835] = 20'hdf7dd;
rom_uints[836] = 20'h3f75c;
rom_uints[837] = 20'h300c4;
rom_uints[838] = 20'h10f0;
rom_uints[839] = 20'h53fc5;
rom_uints[840] = 20'h3f744;
rom_uints[841] = 20'h1735c;
rom_uints[842] = 20'h53c34;
rom_uints[843] = 20'h0;
rom_uints[844] = 20'h334c0;
rom_uints[845] = 20'hf1fd4;
rom_uints[846] = 20'hc7f5;
rom_uints[847] = 20'hc43;
rom_uints[848] = 20'h3c5f3;
rom_uints[849] = 20'h4c30;
rom_uints[850] = 20'h4073d;
rom_uints[851] = 20'h7c730;
rom_uints[852] = 20'hc1331;
rom_uints[853] = 20'hf7100;
rom_uints[854] = 20'hfc53;
rom_uints[855] = 20'hd1f;
rom_uints[856] = 20'h74dfd;
rom_uints[857] = 20'hc3f57;
rom_uints[858] = 20'h43f5c;
rom_uints[859] = 20'h4330;
rom_uints[860] = 20'h3131;
rom_uints[861] = 20'h3c4c;
rom_uints[862] = 20'hf3715;
rom_uints[863] = 20'h31cd3;
rom_uints[864] = 20'h43d3;
rom_uints[865] = 20'h74f30;
rom_uints[866] = 20'hff54;
rom_uints[867] = 20'hdd703;
rom_uints[868] = 20'h1c03c;
rom_uints[869] = 20'h403d;
rom_uints[870] = 20'hd737;
rom_uints[871] = 20'hcf431;
rom_uints[872] = 20'h35033;
rom_uints[873] = 20'hf3301;
rom_uints[874] = 20'hdd00c;
rom_uints[875] = 20'h0;
rom_uints[876] = 20'h40c0c;
rom_uints[877] = 20'h4c0;
rom_uints[878] = 20'hf5dc;
rom_uints[879] = 20'hd03c0;
rom_uints[880] = 20'h1747f;
rom_uints[881] = 20'h30d44;
rom_uints[882] = 20'h400c0;
rom_uints[883] = 20'hc4434;
rom_uints[884] = 20'hc03d0;
rom_uints[885] = 20'hc00;
rom_uints[886] = 20'h3d14d;
rom_uints[887] = 20'h1000c;
rom_uints[888] = 20'h331d3;
rom_uints[889] = 20'hd000c;
rom_uints[890] = 20'h1f7c1;
rom_uints[891] = 20'h300cd;
rom_uints[892] = 20'h474c;
rom_uints[893] = 20'h377c7;
rom_uints[894] = 20'h753dc;
rom_uints[895] = 20'h5df77;
rom_uints[896] = 20'hc0134;
rom_uints[897] = 20'h3370;
rom_uints[898] = 20'h7343f;
rom_uints[899] = 20'h4f43;
rom_uints[900] = 20'h7c7c0;
rom_uints[901] = 20'h44fd;
rom_uints[902] = 20'h5c07f;
rom_uints[903] = 20'hc0404;
rom_uints[904] = 20'h1f703;
rom_uints[905] = 20'h1dc70;
rom_uints[906] = 20'hd30d7;
rom_uints[907] = 20'hfcd0;
rom_uints[908] = 20'h4c5f7;
rom_uints[909] = 20'h1ccdc;
rom_uints[910] = 20'hf0315;
rom_uints[911] = 20'hcf10;
rom_uints[912] = 20'hff440;
rom_uints[913] = 20'h4d7f7;
rom_uints[914] = 20'hf370;
rom_uints[915] = 20'hd10d7;
rom_uints[916] = 20'hf0103;
rom_uints[917] = 20'h40fd7;
rom_uints[918] = 20'h11ff4;
rom_uints[919] = 20'h317c0;
rom_uints[920] = 20'hcdc1c;
rom_uints[921] = 20'h57330;
rom_uints[922] = 20'h1c0;
rom_uints[923] = 20'hd1cf0;
rom_uints[924] = 20'h300f5;
rom_uints[925] = 20'h371f7;
rom_uints[926] = 20'h7d77;
rom_uints[927] = 20'hc350;
rom_uints[928] = 20'h44f0;
rom_uints[929] = 20'hc1cd7;
rom_uints[930] = 20'h735f0;
rom_uints[931] = 20'h4700;
rom_uints[932] = 20'hcd743;
rom_uints[933] = 20'h7f513;
rom_uints[934] = 20'h5f43;
rom_uints[935] = 20'hd17c3;
rom_uints[936] = 20'hdc31c;
rom_uints[937] = 20'hcd71d;
rom_uints[938] = 20'h10c73;
rom_uints[939] = 20'hcdd71;
rom_uints[940] = 20'hf431;
rom_uints[941] = 20'h3c4d3;
rom_uints[942] = 20'hc0777;
rom_uints[943] = 20'h31f31;
rom_uints[944] = 20'hcd310;
rom_uints[945] = 20'h33c43;
rom_uints[946] = 20'hc0;
rom_uints[947] = 20'hd174f;
rom_uints[948] = 20'h7cdf5;
rom_uints[949] = 20'h407dc;
rom_uints[950] = 20'h0;
rom_uints[951] = 20'h3101;
rom_uints[952] = 20'h4fc;
rom_uints[953] = 20'h41330;
rom_uints[954] = 20'h1cc;
rom_uints[955] = 20'h13c3;
rom_uints[956] = 20'h3dd1f;
rom_uints[957] = 20'h70f13;
rom_uints[958] = 20'hf0713;
rom_uints[959] = 20'hcd147;
rom_uints[960] = 20'h10f0;
rom_uints[961] = 20'hc1743;
rom_uints[962] = 20'h1fc1;
rom_uints[963] = 20'h5f773;
rom_uints[964] = 20'hc44;
rom_uints[965] = 20'hcc1;
rom_uints[966] = 20'hd3403;
rom_uints[967] = 20'hcdf;
rom_uints[968] = 20'hf1f51;
rom_uints[969] = 20'h4c33;
rom_uints[970] = 20'h3dd7;
rom_uints[971] = 20'hf1331;
rom_uints[972] = 20'h445fc;
rom_uints[973] = 20'hc4c3;
rom_uints[974] = 20'h14fcd;
rom_uints[975] = 20'hd71c7;
rom_uints[976] = 20'hcc34d;
rom_uints[977] = 20'h3c71c;
rom_uints[978] = 20'h403c;
rom_uints[979] = 20'h40c4c;
rom_uints[980] = 20'h431cc;
rom_uints[981] = 20'h7c300;
rom_uints[982] = 20'hf71;
rom_uints[983] = 20'h3c310;
rom_uints[984] = 20'h1f10;
rom_uints[985] = 20'h43;
rom_uints[986] = 20'h37dd0;
rom_uints[987] = 20'h3ddd1;
rom_uints[988] = 20'h4f1ff;
rom_uints[989] = 20'h114fc;
rom_uints[990] = 20'hf1dd0;
rom_uints[991] = 20'hf0;
rom_uints[992] = 20'h31331;
rom_uints[993] = 20'h1f343;
rom_uints[994] = 20'hc7731;
rom_uints[995] = 20'hcc74;
rom_uints[996] = 20'h433;
rom_uints[997] = 20'h14ccf;
rom_uints[998] = 20'hd4d33;
rom_uints[999] = 20'h30;
rom_uints[1000] = 20'h41ff0;
rom_uints[1001] = 20'hcd7f1;
rom_uints[1002] = 20'hc0417;
rom_uints[1003] = 20'h3f051;
rom_uints[1004] = 20'hf71;
rom_uints[1005] = 20'h4c0;
rom_uints[1006] = 20'h34cc1;
rom_uints[1007] = 20'h5fd07;
rom_uints[1008] = 20'hcdd;
rom_uints[1009] = 20'h73dc4;
rom_uints[1010] = 20'h3100;
rom_uints[1011] = 20'hf5d4f;
rom_uints[1012] = 20'h71033;
rom_uints[1013] = 20'h7530;
rom_uints[1014] = 20'h1c3;
rom_uints[1015] = 20'h43f74;
rom_uints[1016] = 20'hf131;
rom_uints[1017] = 20'hf01c1;
rom_uints[1018] = 20'h375f3;
rom_uints[1019] = 20'h344f0;
rom_uints[1020] = 20'h13;
rom_uints[1021] = 20'h1c07;
rom_uints[1022] = 20'hcc1c4;
rom_uints[1023] = 20'hc043c;
end

reg [19:0] outputReg;
assign out = outputReg;
always @(posedge clock)
begin
  outputReg <= rom_uints[readAddr];
end
endmodule
